��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��^A�-�;]Q�S/�pK�:�b����ԏ�1����N9�w�#l�w�Q�@D���G��4;�`/��C���Լ?B�ś3��
YR*/�Kfi���=��Սl���� �diA<ꞝ��d�g�ܲ��I�7!���U����߅����E��_5 ���dդ�\�a�������q=��"�q�8QON��Pҿ����)��g��f����.��"����j��aS
԰�e@� �am��M���=q~t��;���s�۩��1�G�<Q����=�t!Pd���!XI�����>� �|e[��O��0�=�t$�ڄu�W�����v@�`�G��^S��ڶ�$t�!��~K�X	
�S��o��`�[�c���8n	�)��֣&UŰAH��O��NH�[=:X�0,壆7�i1��9c8��MC)�7F0u�:}��HXcD�j�$t+
�-��l��h�?V���O5 �V���"���������kϸ��H#,�&���V�~��`��tr ��g:5�kLdkή95�@e�0/[ S�����}�N���i�n��3:3��~[v�T�s��j��V��H-Sb@�Y]@�)��GX�]���y�UaZ�r����q��y���;q����
B4UѰo����T4q�G�/}ۑ4d2�#��B���W�h#[ɪ��ߩB��u<����z�t����K���l<��a]�^:�=t�s��;[}?a�J����^�y? >�N:��,�3���;~%.�^{N�l��&�n����u_�5��z�pu�����;�k����;l��Z�]Xo�z�;ɬ����ٶ-|?sѢ㉫� [h� �uA�\�Aہ�;R�[#��]
����	�O�/|�uoi�����o���X�>��Џ��,ݫ2�q+�7�qS"��N�_	?�βy@���\C�?0�1��˦�5� ��2Mh�W���P!��M��?z���s�ɳx�����K�⮆?1���wn�X�Y���Li8q(}�$g0���ϫ�>�LX���a~��Sba��6��No��Q�]�T'3���n�����[n|$1ƙ|س�#�#�����Q�-i�U����9�96֌I
�U��.�KJ����)����L�������w.����	�����RA�6ٌ4=AŠ(s�.�7=Ȓt���N�H|詮ػ���_��8�F���V1����DS9����*b ��3͚���%�����l��/��:��L�Õ9�*���M��Q�����ۜE�F�"vM����lKCYa_�CuWܧJ�Q	�@D�=j"Y0<�(�h!���v�.z��D_T��t��kcz�5Z79ϙ?�|��$�z1evu98<�tw"��� đ����'��,ZY��QK \�Х�@*�fg���M�H��W���� bcx�f���V'����$�]�6�� �i�`�Ɇ��K[���Z�������o�y���3ڶ�a?�]�k%t�4ua��{	|ӯ�C�Hu3ql��?�>����A�@�'�t��5�|���D���26N��Q����{P&���:���(�}qzg���-��y��t�hK�;�7���g�C[xamu?`:�� �QP��Ӎ�B� $�k��3�f�����0�<(L�p"G���nax��r�))R&���d��Ǣ�X�ț��������±d���XZ�b2a�"�%�,��h�T�ӈ�{m�=4N�� t^���49���.ǅ\8���#��#�U���G4��T��u�IN|�!���vC�;v�~�	FMD�~WC���/г!r,U���)�i�)�]��$��a�}w_�jYÞ��r�!h�޷Nl���3�>�%V�;�'!W7>f��4VD����٫���b��Ap{��b$����#[�>��Sn�l�6�4CD�Tc^m�Q��?oA�	%z��3ˠoݎ*�:���%W2Ș�S)8$/�YM��,j���w��i�h�(�5�:��?V��@����a�N�_3�A����.$��y�KD�ӕ��дW+/���Vz]l�RmlL¯ţ��G���V��T�8k�9��W��il�ْ�=�&{b�oI�.5[�-\6�����x* x8�������B�6�d�y#��C�s]�8�����n~.Ֆ8�/_�L�����c�k������P/�|0u1������CB�Ϯ:nAҩS�2�M���� �ݭyns�rr�T ɽ���ɥ�ܓ��^�b���Q	�����M����f��'��_�����:��O?��_�����>�n�S�	��bV�f�
�\M���E�2����c�t�.{�M���e䏞�yEM�a_�R�K�b4M"Ί�7�n}�a�[v�gP�q�%Bw(6�j�����ÒG���NM����,j�A��wM(�Ǭ�q�\뫉_@XR�ll)��x�,O<��z��P|����r&/��b=��Uc+m)��c�����g��\ی'H��0+��-��x.!ΛG,�1ƩB�E�{�ˇ���g^��A����L��Sw�(*R �#��1�����h\���E|X�'�A2��U��d0���_V��G���>������ wb�{Ͳ��%���}Ŕ��`e���.)�),K5��_���uyS�<2I�RNKƦ��=L���X�L��mm4
�p�3=�d
���&����I*3��j
ZX/t��B�s���^o�&|�R����)Jr>� ��ܶ�y
�o�A'Ol�����F���E�C1��}��a��Ţ��%0�=s�C�1j=K����3��(˗��nW'A��e�/��'�:g������im�-���R�Ñ��8��\�]<�x��]�Q{�&�����&�Vs����3�\�&���|���w��`��DӘ�ƺ;Ox���MT��a���{6�W���pnw��n^��+^���T^?={O�
`4Ȁ5����-z�[&�w�=�O�%Iw�"�g�� /��O�Δqo�lG��qfL�վC�%֗�	�� l`t�L1(wq�o. �ʸ�|A�*dor�fm�|��V����m��҈/P�?��\��&�����6j�+��ڳ�y�BP��u�x
��#�e�J��Qr92�y�r��Ɔ�S�2OI$�?[V���_h�����N{k	�<~��i�u����N�-*��;^%\�Vwq��Ȕ�5\� x���q�V�Zy�T��Bf
�`x��_=�D�������e���̰�ss�f��U�I�^*h��:쭝_�t���ym|�p�6��z�)OB�!YN���0�u6��f9�k��Г��k��OB7}�^�g���ϝ��Ж�ߖ
Q_zd�a�n�9��@'�q��[�`+s�|��o.;�`)8��t��~��	��,�ՙN	�S'�#�5�sR��W��:���7�g���v����q�A�-�n9�n��?|;�{��H]�����6��-��謕�7�֒N�
�.s�n��S_/��H��ϭ�X�?,�vaf
a3%�Jt
���I�����a pY���P�
�d]NM��1d !�a=�'��)��n�"~�O��*��Yg1�*�ֵ�����4�{�aA�y9��٢C�A��\��I��'�b��;�^������::���L��[,���p��#/E�7���7"�0��i-`Ы}�b�͢�^�p��3�d�F�%#Ǯ�T��
�D�!ד����՝��fO��|���0(
x�/&G���-nv]�A��~_TO��+�������A/�:v�t�d�X��H���v������Q�Zm�vt�*7�&e���P�,�|<�j&�ut�R��g@&��xiN��i�EnV����EMG�r�/@_{]�{�8w�mn��`x�5>>Rzk�%�
N���\��S~
H��̘.Bkϻ�'�|t���YQ]~W���dsn�s���B*�M�y��ӿ},�'&�#���QX�Lt�e� ��V���p/> !���<�	oS'+��%*b��]8�jNL�Q|��(?�w�}u,V�A��0�2��`3��˃!��R�m:����X�D�⌒ q�z"3*��N ����D�v�f�G�?|��y1���MA[,%�<$��#�Ț��8�(f�p�n�n�B��`3W���ңm����8��!0k�-'�W�7\r�nf(�[�b�%�tg���I�Y��bo�v��1�\2#L��X��\�=�{M�R�Ō�m>�L>h�7�Jl���]��XlǱp��y]7�nܑM��K�椾[x�*�yN�����5�^ '�l�W�G!���N�b|�6�r��<�#1��gA� �K�?8��62��\=�����v�zX�g�:�d0�F"��	��gO���N���H�EMY�T�.���w�&��e@
��D ���l/�꣭ m�_w/M���H�[z�+��5p9�`9?�6��lA.��8i�k��ܘ�����8�N��ꢀv�}|]��o�Y���#@b��Z��sJ#�!?S�~�DD:���[����a�o
.yz��3c�$Wq������K	�Bf$��>Ko�D�d��@���$��EPl�o#c���q���v��kB�^o�"9[P18��� �A��,ogވ��z������!J��x���-Y�u�����V��mf�bྑ����e0h� ���p,vZNm�K-�j�O@�n�%���Ĝ*���tZ�0`�͵W�C��Tc�xW�%��l�aT�C^���CŚ����s�c�~<3�	���H���hp��jZO�hA��a��� I���.�ԭ���Ԡ\�zʼ|c��d5ے���l�����}�&��K���*
�J� ���[�מ4:���2$�3�CU�\��[[���R�e#�k1-�՚r�=�����ϴ͹���7'�����)�s�::g�wr��Y�xz!��Rbf�'��@�'��<�n鵭>];�i_�`�+g-�Rk����-Lm���6�P�S���m^�e�Vb�I�l���� �M�.4ܞ5��&[&l�wm��n|�+�����We��W	�ǵ�8��S82��<rK��.?LSa�qI�9�.�mR=�!S��/�3����X,�=� � r4��Y�8�Rh2g0_��S:oL��&�M9O��zk��X,gC3IN�c�����F�W�m�n'� Q7�Z�?p��}���)|��d�H|[+	��iB/�ϊ�������h08w��ݞ��!i{³��k�(c��������ص�b*�r��3"y�
W�m���a.��Ug�Q��럐~�P����)lI2��lA��§ U�s�~��������}��V���<�^�䭬��/����)Q�W����ڃi�0�<�r��h��H>-��{0'���QZ�g�C�oA�;�6PbU ;j�ױt}��/rl���;�1�-c_T��[4Vk��;jmJ�R%m�9Q����F�g2G(x��N�CU�%Z�vR�q����+�'$#���P�#�u�_�_�r�7|#�\�Snx5��Ц�{R
�N9�e��1�*�V��]�)v�����:�<�H�⟜��Mw�Q�%A]�&�Iu���i��4�G=~J��z?,���^ל%���%�b�У"9*,�K�6e+�E�#�9H�2���d�����ΰ`'���j0�ͦFޒ��Q���ŭZ���:��W�4�E�*]}�>��$9��
�_�)��/!>�u��a���mK��MG!*8`� sq��Z�$�{�	�Z�BY��v�Ye||Y�\F��Ǌ��6��P���T-�ağ�N�"Ż��F��Iufd��j��23z�.¶kA��ǝ���xn���<o������)e'�Dln�#�$���&�����k��n���#\py������z�������cW�6]� ;讶�G���㒫)���2'@���k%�EAP��O�R|�S<v�>EPQF�tg��k��Va�@��rԢ[$�`�\���h
E��c��X�7�rq���@��?�5?e_ck�4����׉}\�
Hy�D�z��E���c�;;K�����=��pĜ��F������O��d�a�4aLɎb� ��D���G��D���,?Xق#	
����j�I}̏�7��%%ſ����n��(C8�,[��Cנ��1_N �b�V�}�ql�}ޫ� ��~.��Rj���;QTYbw��kn����Zf�M��0JU@�P�D�,�y3o���y�9#,
S08����Ŷ���Y�w/��(��f.Evv�7��g�OA-�C�.�:�@�Xg�]��t���l��`��ʿD��;'������U@4֒E��t��O��sRuZ�y�a�M���=*�_��--мÏ1�%�)�L3�c�0�M�G��-7/n����dV���tx�稚^z��c�����e4R5�'A��@���`+k~΂�eJQ
z��Lpj�D�UGLF�N�A�jAq52]�;�]k�P���x�2���R?�N��AHZu�Ĥox ��nҀ���E`��tNQ#J[@[���D^�C$S�ܒ�H��2CG]�vҐ��^P"�%:[f�:N��[�x�?W�\T'q��@H�������=���
BJ�3�3��>n��֗{��r;�5�i.l_I�aX�(���u`aƂ�˥��QBm��?ur�b߼5��*D�j7B)�@�y��:8����_�哣%�̼��BMH�~��ۈ���&���V�>4��6v�lef����G��p/
�3�}��?њgZ:�WB!��Q����BI�!�������:x�����_s3��0�B��}��+�� n �<�=�S��y��(.a��4��I�,ƣ@�#;����}�i�����\�^Ս��D�v}o(|�3�w`<���,}�5T�3����ѝi�= ���yf*8:	е'.*�_u�~ׇ��#mF?EZe�q��k@)#�Bg�pG{!{�C4��C�~,�����@��v��NrOؕ .ގ�b<���Mq���x����Є����AWAw�:�`wFY�C*d'㴩���f<ã=S�dߏ�7����C�9E�K�ܸ���dY� �y�*u
^-��y�:�u_]K�j9���M2�-S�];�K�������xJj�R`a��7R{�� ����htq[�"�	��l�D�L���?%��pG$!�?D�u�����>���7NU!=M�i%���v�����T`6iAFi�BC^�b{��6���g�]�� fa;|XG乧�Y���j#�oB��-��;#�{�<��ŋ��D�n���!��NeX�c$�g���Z�y�D{ή;�M�[Թ�8A�>�?��$D�?�5:(v����&�uG�<�8.M�xV��&�u�R5���;�&�e��ؿ?+O-z_+�:��NE�}�u�n�$�=B��\�\	I��#�E���sD�E��\�;��{F+�~��֐D�
>P���u�_2p��؋&��C���I(��S���,)�鏝YzA+�͜�}Q	������:d��eA�h�3�!O�f�A�JbL�6H�ܚ:�xGێ��O�<-f.����B�!<ݐU�S��P��'�]h��t�˴1S��4a�L�*��h0U7��q#��	�)���\����>S�-(y�S�-b!��3m� Ј���4�J$��4=���.s`"�m��K���ƣ
��e�1�-:�k���A���8��u���9V�����-�'�>� Y���H��n�L������5�o�-�e}�,��>-��bG��Ɠ1�|B�9��,/R�h���q<p�sC^�=��S�*�:���s���&�9��Lv��j@rR4Ben�ͷ�d^cP� ��7w,�&�w��3��� H���8���c���@�n��e��a��ǹ>茧��ߪ˟���哤(�m��=��%�d���?�T�,4�rW�Q�9w�qN
O��6)2GZ/�z2"L!*V8}\a�|fV2�w����D�q��8��nͽi��Hx~$�	-Erz�&0? 	|���D��!��>4P���K��$3I���+,�^�y��	�Q��z`;tLo�G����� ��k*�E\��@�v��q5���!��.�hR��L�˟�_�����84T.����)}�m)�N�4Ԋ��>sԫ3y�j�U��Y�ȓ��B�r��;Xa:��J�֗f�:�[�|��}98e�(���b]�>�S�|��e�Ŋȗ
���n�|�X���$�������B��N$eq_�L�(Hv�rf�4w���q��rB_�1�hW�������P@�k�4��?;}�M<y�^�.n�h'������HM���}z3�a�5VL�`q�jl�٭�����_+�N����Sf���j,J������}B^�vy�#��Pqbpp[s�#�t���!�bA ��k�0 'v�?��=*M��q'h.Go����Jg� �!No8yh��TaS��!r�9!�Ѹp$c`g���J�Y]�<
Z!�@�/,�U�O��yd�^��8��S��g�y�T�Q�j.6���y��m�d;XI������1�~͐��c��It-Ѝ$`�W6s���.3>9�%f��A"]eE{��[IG���.Tn�{�wi�<v<�)�VTM���ܶi
��f'C�<�}Ϫg��u���U��ҫP�_�{�b[�E���%b���N�؅D�[����,�|,�M��r���p�L�������S#�p�(�����KP��I�e.�k#bG��d(F[�<�љ���&Uʔ�!������y�l������AlQC��*;�]�6�p���������iq^��c�

M�	�P, ��M[y���*�M?���@�����~y˙0�B{"y߀2Y���PO�E8�4$
ƬL����kb^����~�8�)��.+�N�`�Dx�^���䥁k��&��
\�S��}+i�Յ��<k�ltM�0քR��H�l�f��?�kGx�t����M���} ��8��'�	F��
�tC|����1se�ձ��4�>ϋ��V3�;���!��W.��ɥQ<��)�t�m!F�}I��S�[Y'$B;�|���N7�y�;h�9�I��ai�
���5�}�OS7��KasRn����?zA:��R�bkk45�֨7Rn��,�6zN�������V�;���]B�缩m���j[��8�LC,t�:WT+���9�5z��A�cZPYXG=�}�h���r��LmF\�@y\�<�┆L	�Pv�0�1}�?dc՛��|����v� x
]����&p�jE�T�щ���v�@���#l�����>�����T�G#7��c��z��<�n�mܕ�ީq�qA<ڃ�u���ʻ�����B���2�W&���sG����e��M�7�VV�w�Nyz�I�����j���ssx�/�����,��.z�T]Y��Z�ڔ��/�;*s-�N��{Z���De����5��8��;3�ã!�(&�4�yi�7M�b�����1GuXVn-����g�� �CT����3]��Q8�4RJJ*����B��m�b���(�Q�=.\�Ef���5�Bl���diW.<-S����r��C�%f i�w ��j�3��W:�b�׺�ԇO�	�h^"6��Y���aO~Q1�%˼\�D+�����-f�V��S�d��8�dYp$Yϻ�l��g;�\�������.�
e��0al����׈�K`�C�\ĄrÕ>�CȤ��B�), �9�7�.G�����q��5yD������֞m�ए�¡��L���/�3F)he�N��	9��ܠ?`�9>���g�\�����E�ZҕZ8�j@((���&����e��MO/��s �j�H����0�ON	{�v��y]����D���n���^C�X�\=ۭ�2�c\���-�G��S���0Ǿ��{��>�ی���YPh�2P��V�K?;eWfF�v�w)�/�B�i�j�߫9@����*'Mv��HQ�Q�P�;��jy�jjC��r���8Y���䊳ͩ�wXw`� V�?1����4��b[��t�j��@�eC01�6M�]���{R05�1�o��h�^��_��1�H���(Տ(�^�x,��
���B<��9ܤB�߾l��u�F��M�f�5"�	����P+D;L�Ĳ�Z�(�e���;�8�� �_d}���F�m�-Q{�FW�Ȓo�ܰ��6��g�& �.e\&�+;4t�d[�`<&0B�RY˨ �;L���������E�����V�)e�&0��o�Y-�]�]�FZ��M_`��N�f��q5&r��d��y��GM�ҘI��:q֑��K�Q����34j���Bx�)����d�Sk�C 7��4�PD�r��*��a˩�@��{��q�D�қ�5"�S\O�!/,2k@Q��ٻ����|]0t��(�2� �����0�7I�$U�h�GKz,����1�pM"�f���Z�~t8�@r�y.�xp]�^��$;0����&('�[�.@���K�=7�U�a1}L8���6�"���\��?R�H��pDi�8�& ���$����F�������kmf�*G�=�H��lP�%��qvѮ_&Νɐ�z��G-���d$LZ������B?�v�<��Ǯ�q�BN�xn�PW, ;.�.OgySHV�Z"t�����fd\���k�GӘj����Z���L Th�䯎]��钟%����'Ag		�(:�.����/5Quh9��T�d�(�I���ՓR2�LE�����@���N ;[�-�g��9��|�n��l%��N�SO�1|�CZ����[���Bܫ�'�'�?MR�&��{+�l���A0��
�:T���,�� >���c���=�tX�"�܌�&
*�{�؃K��B���:Al����W�%�d���$��,���0��͛΁�5��0g[xz�(�����[��oV�t+
ц���ɳ�W�&�7(wJO��ov�>e�L��q2��Jgx.{��v�JՎ�-���'֞�D>�s�f� �S��Z�PS}ո�`�R�ӵ<$6y�	_[�PIIb2�B�\�yS��!VmY����X�'*�s)�2,��F	 �;�`��4��T
'3���V�[
'�N�[|t���������^��Xc�����~N�A���ԕë��G��ߤ��*b�#���$���SOz�R��0����!*���l5��.O�4R?a&P �һ����`�ݸt6����qk�	L-�J|��%���ʮ� R,a�ꊨ����h񾜘0���c�t@��2�ubo�ߔ�&����U�B���:���{�� ��HD8�t䄣)���K�w�.`��$��pM�h\��\!�J�1Զ&���)���as��X�D�RYJ������`�rYL�@M�q�Lrޢ�nZ7_�y�\���9�������s���cz��5Ҥ�히�cpđ�Y�7�6C\���m�����"?���Q/[��_\��O#Tܿ���Q1�L��I��Y��DE��=���s��Н ��[x���f-}[9G*��:��'�����2�Q����|�p����, -�w�a��2t�)Y�o�9���Y�ˇ��b��٧�d7����q�k6�}ٺ�� P��X��ڋ�zm�1���^AlHcT��e�j'�_�#-BE{�4?Zp4	��͂-4��z�me#�j�ȹ�����A�̈ém_pBy�	�}Ζ�$(n�|\�;�,�e��n�K ƓO�?����*��^�R�l�F`�0tP��B���oEf���6��L�����Ǿ���"W�f�2֤Z�FYiO;��a�ꑵS�D��(>6A��|gg�YA8�ĉ���l2���Er��4�^���d�H��y����Zr��h�˫���(?�<x�7�C(��r��h	��:-��Y��=�ѕ1�0g��� ��=���M�z��Qޅ�*�]�5!���t��䷅���'�S���a��f�LAo%���lޛx��;I��]�
6 C,;gIñ�����e'��y����B/Zp-��t�f�G���#Y`�z[�����}�K���哂�U�Lu��"?V6�����d-t� ���f�{� u��oS ��4K���R@�m�{�?���Q�PwY *wd�s�%�"�8��A4B
y)/�R��!��Çg�_�:e10 �Q�8:�H��Z�o�2#�
TyB ��sZq��="���֤��V��45��6�wOS�@)4�Ky$�3�ت8������t_����	r'����03�Z�ݞ#�6�.mmG:�V,hf�P8�ΏG�cP�kVCn<O���e#��R�c�T;�􆻫��@���-I�ܗaP ��kޙՃ�r�a�I��$�M��N�Z�FjIWEFܴb��\���&���_$�.�@�OAviB�d�s�)�zxV^�`֥�{C��|�x�N�e�@b7��.�D[��nh��Pn�/qw��+*_�kʨj
5>����nZs�룈yMxD����2�+�zY^�lgsr[ZNC������wj���ǿRq��ҟ�+!Yc�\J�����
\����`H���ЙA]3+Q�i��i�s[	�yF����E�ҰR�S Zf�3W�N���'CF�˘F�l�L�g�!rd���������FNsy/�oP���;"��V��(ܰ�
V�^Ý�*qkU��c�>�^��2���^AKa.���Z=�=|כ�!�n�$9���k^߶�y�੉w0h�|�o����q�8�s9Yj7���c�Y�R.�d޼�W��y�;sĠKyz�)���p|�JI���@)���c]}�	U��Ϡw$po�;$�8��=D�腚Բ�R�a��U�r�Ț[��m+:��&���Uݞ!nL��ش��c�sqZ�pDlm��`ݨϿ�"Οɻ����=�r�%KG;�"k��s�p�Ez�n�wYW��31uY�qV��}���"�We\|Xq��U�#�Z�U|�O��kƾ[ �,L�D�gK+Pܓ����j�ه={��%��M*���
�ꄖ^�>C_��P`]�����֑�Lh��zl���V
�w�?��.�7�ɜH
`Y�F&�Iz�X
d"9���g������;�7���9�����WL�z/'c�J~>�?;n4��g�~h�#��3o��ͥ�x��8Y[@sS�]�����%�V:%^�B����uDOH��4C��|1Y�|�Q�.�U��J�"V|w�n��a���g�CCz��h�Ѹ+T�]{a�Mn��jyW'�?��9'l�At�CY9˫k��U�M�r�'���
���f������� K<w��=�eiQ���g�X�s����;5���~:��'c$��,��n����Pq�$�@���'��Upx
��Y�L�喝��Rf�Ы��(�9ݣ2�|�[�QTo�=-����͡4���=v��0~/c@�ͶEow����R���V���C? �w�B(`+���\ѱ�e�jL�ʁR.ݚ�g�D[�.0�|�h�k���'�ZȐţW���0J"GϩQ�M|yد�L(]�6��@�P�_�b\�,��^Xl���#L)�����gD�X�����Y ������������O����;��M?6�����G�X@��I�p9�����t4 ��3�JCGԞ]�P1�umq�E�C���Sw�q#�;��1��V�0d ��[��+��0XD&�@�r���؏��<�	.�����a#�+�=�W�5B�bz�[%	�(��*�)�x4�b>���Wc�r�T>��]+���x1m�m��̕f2���m�DXh��������i���b����YT�^����/D��d�
���3�6�+��z��G�h:�5F	j*������Ӧ�0j�v��a��9��,O�.�YL�����<�ͽ%܇������(��g�G��]�{�lI�}����p�dn(����N�y
�����5^x�!_aQo�Rk�H��T�X������L�r3L͖��*T��ϨTu���%n�X��+���nkb���]*~p�[� �K��@#�KeQ�7�p)}j��EZ]ܼ���I#�Х�k��
HHk}y�a�҈�K?���>|os�ڦ�R��M�@��b���fW���6&���]��h垀`��d��Y���f���ε�lUoo8%����#��q�(��n�4շR&I�ȧu0������Y�T��ו�����I��6����}l%螪���I�*m	�UgeKQ�q��m���_��8!�^;�?f� 7���M�5��� �u���W���&;��Sx ��Z�h՘�]�@�����t~�TW}I��\8�ֺ�Ώ��T�eR�m��vh�+�T�j�Z洢���vJ�VA����\��$���P����瞲�z�������c&2'�yG�9��3����k�ȶ6li����a9��l��%��Q��+xhb�n	��?1�JMl[���Ol�O)�4=���s�g.�ܺ ok۟x�$��qtq�-�^)�n�}�mH�U�ܐ �!�:�C�	�h��n\�@_Kw���-�><m��}�n��Ee�9�R�C��;��6�{%�	�e�<#��|�k)�N����8��QݖT�3mi�B�5Q�(��U�X1����ֈ�X$����u�~p�.�"�L�)o'�edUAť�W�N�r�.a����6��i��\N�\sQ�����얬�?c�<�;�~���r��UO�J��b�h�{r����<ݟf�����7Ѝ����EC�Vd���"a-.�o~b�F����)�	��l:�h�.�kS���4@�@u���1�������]�+�#a�K�>$b� �K���R��$�Ih�%��#���g�X?�]��m쒷�ȣ5��EC��(��qR�� ʈ
�-#}�D1t��6J�E4��u�?����z��\�z����p���4���<:����]Шwa��|�}��ʱՊ����'�Ӊ����~H`�|���F�߹�G6 v�A�k��z-��Ń�6w��D*�v��N��aA��d;e�d)����[B�nB�ȫH���xXq~r��γ�9�⤖;4m>2��LD������ގ��Jczy�<2�}p���t�vC��Re�e�5����&Uh�l��>Kw8~!st���Wa��8�霾1P ���Z>|CM-!�b��@>q��~jM�L)��k��U�=�Y�I.J��M�����7����h?H`"h�SjI�:�4(/*Nq_�+S�ĊcY����ߒ>���V�E�=R��"�g��DB����ZR��t,��֔����Dq8�Qp�p�5�c���Gn���L�$���m������O69ӟLl6'������,��C�B+}bZ�F�}���F��� �~X�b)�-��߲�D�XJR�J�f^�3�<���dv�4C!	��H>2�ࡎ�h��aĥiܛ�W�Y�����nf�gg��2ψmp����K�T6��F�y@6?W�<�P�!��
(f�{8�+l�탁-q� s@͈h��(ԾŶ�Qٗd����x��2�f
sf�����ѡ`iP�&B���|�D{sF��j�=��G�{��8��i��lm)*�=W��1S���[b�u�["���Q�B:����v��}�r���VZ\Bm?�Wgo��ަ5t�1�lP���3�P��/Y�0���ᦀ����ʥЇ&�ʛb �&�R��<J14-��TCp��b?��S���Ti��Q�TbMKA��U"�!��ްZ�n��ͥR����:�D-�k�N�#г��Uf�V�dY�ZDb�>�hv�{��������L���\M8^MTcE4 )���;A�ks�6�͋���ga������\m�7��d�oC��t�:m^A��ɲ���L$i���/�l�0�$w��rm��6VaMU�)�����!|˸������^ҹ�
ѕj��x1_����w�3F�v���p�=.= �B��g\S��St:5�e�wCA���C'$����o9�hhn��IX?��g��ؔ���M�j|ղP ���z��������5�G&dMgg�#Ĵ�8�E�#�1���H��h�v�C���nO^�"��j���ށ�(KԿ�^<�g*�@2��;ʸ���Sq�>����=���$RWP*&�0����M�7u��Yɴ�3��kxe5�GQ-h^'�
����b��dl%b܌�u'�]��}�)O �"�9ႆs��į�+�t��y癌_L�R���X'��#�d��^	���!�QVV��k���	����Y��Y�k�T�H=�����6�ʋ9��pM��d�c�~�ۿ]Ub�0q�/�i� �E!�Rb��>�[�">"疁�Қ�����:b��Gez1~�H�����F�[D]�R�c�P�GPmVV������	2z�>�Y�i[y�7R�`ևi�X����r��)�Q�XO�%JQw5F�qbU�B�+���G��P�
xX�H�pÅ8d������x /�H)_-��,�(��'�f��c^��N�`�K�	o�_��^�O��^|�y�ŨK���C�n���N&&t�G��oK�ӎ�Ų� ;��
��d��d�Jxj/�/w~. ��K��F>b?�!�����c�w.v$�v�B�oMx���}�j�br&�[?��/=T�o�g���w$:������&��~�;^�t{�m�k�9�O�h����fgw���r�R}0qx0����X�b�ξ�Aa$��OG�<y�:]��_FiT&u�"�=�Ǵ��%PJ�p����~z򸆋���������p���8��f����ݤbgR���F�0���箦�횝����/cϵ��'
$�%��"�t��Q�cN� &?du��%�'�;�JQ�
�Ow��d�Ĵn*�m�=�*E�a�P��8�+y��¤��4�h��J�[/�/��8�x��c�V˫�Z>���D�Dس���<��ae*jR��@���e:��`6N��v�c#(��3c�N�WIw�t�ơ|#u4p.��U����у)V4
�J¦����|G�:�7��1�;$��D0�	}��x�U1�>�C0|V�X�gZ'zf�XGi�`qc��L��L�/�,�:U�'����@:�s߲�K�f�<X
pZ��7�P����z��s��K�E��O��fB��&��\6��(���&H��Eg��	B���`�;�y�h2p�ZJ����U��v�U$�g2�Oy�ad��Λ�=T���"R��>���@ s�角G�q�����v�m6dp�#�O_CU%v�%_����ǝ�l�V0�D�S��=fPb�R0�W":�e �_~���B3�Np%zsL���� QUE�z���=V�6��Cѓ#��4����<�1���D�N�{�h��J��y�@�f*[�8�s�l�Y֟�25z+����u�o:I�_2U���4�aHF$�y�Z�����Ԕ5u-s
Àީ���B��oT�Uƶ�q�ȩ�s �S02��i�k5N�:��Ws7�g#�x�&
b�o��� dD��=}* �m�U�+����>�Կ�5;x��,4����"�7�����/^BVg[qMc����͂���%S�._?��Ș��ra����I[�"6h��}�����{+DZ���̯���ȍ�b�~4��kn��)R޸��4b�!I��4�t���]���] �v�O����7�(�TĎ�1~\F��~���.���w��8��Xy:��Y3���_x�4�٫�J�a�H5PO-qψ����SJ�"}~���C���6��>�J6�v[�������(���\iR(�V
n.S��b����p�tbL/��?�>}�
�����v����ޑW6�^ꭄ��ѺT��AI����a/�Ճ�yM�P�Y�+�֒���#����K'h���q]jW�8��2Aw�Tr�!��?1d�p�����Z�W��j8�����y��y����e��J�r�gzPF.F׎��{9V��O��{�J&�b�A�ӝ]n�(թ�#���:Y��u' w�ǂZ/�-12�t����ݺ�Zc�>�r����܌d�N��Miѻ�:V�˸Q)��TQG�����`����m���p��i��~?�wnR"���OSա��5xu��g��
R����hLz<hW�'D�H�|O�7���x��{Q����rV�f��!k "#�z�I�z�Z	�W,�%ޮ���:����E���/��kw���T9+�$ V����q�F-v��=�b��4�q��H���lt~���ێZ�[h������kܵ�����%��(���'6��#/��w�zK���5���#�&ă��v�~̮U��!���T0\�+����ס�Q��Jo3����՜F�b`��erˆ��<����>�\Ǉ�X����vC-ܣ{����H��v꾍
xT�ݷ�6����m-@��w�lfǫ�ל���UcU��;�ȇ|�K����qv).��Gg�i�_��Ee��������^r2ջW.�?飽�b�	y���j:��"͘�F3dx|���,΢��%�y
��z�&p[x���fx"@�����F�3%�ƌ�T���Y]�3As�X�s�2e��oN?*��d}�GV����㶍$�)3Zp�BV�v;���k����<r��lڧ����2�<%�1 *�Ge�ǖb �+]�c��L�"��7����j�%�l�k���m�'�Մ=���V�5$����(y6yM�Lt���(��W�V���,e�[;�:ʏ�Ƅ ��Q�|K���$ٖ��v
,��ń�B<��~#����S��G-���\�?M�4�ǘ!(��$����գk;�}h��L��M����ղQ0�x��r�8�1k��¤P}:���3�/!�����J������x�S�n>f)�=�O�X�a~j+@�	��]O[G>���TdK[�;�(�a2+'n��dtXd8n�������|�%�Ә�F#�0*��՜RwS�_U�kwߜ��Q�N��J\ⰳ�{�nQ�S��ͩ{+P@�YbQ~˨��]�{�Q�f�t>�kx��r '�@M�e]H2.,�&ɺ?\��)�
D�E$��U!U���6y�C߬�=.)�^|vm�`����^�/1Vp�y;k�2_{,uo�=�}�$!FS��hϷ����J^&��b������X�$	yxJ�!��U������M3�N:��o��9����>��{l�Dx�a�>�������j���&�����k���7�>_���7v�3[��q�4f6vjeM��&�#���@̵:�/����&��:0 �����.#�;[����*�Y�MR���ZĪ��@���'rO�Q�rC�C���h�ّ #�w��4t��#��������Be>�����I�sb�\*��BLDs�ba�g����9֩�� (���~�߾En�|v;���|��q�����ۘ����	y���0�4fO��ڰ�K[5��'ѺY4:Ⓢ�~�N^���^��UG��� Q5k���d�*Z�=��_66aJ��w=��^f=�v#�Y>����Phu�(ς=�xՖ�s𹂱=�Q���T�i�&��ٍ�X��
�[fv����ey�S�+o�y��i?xL����;wl;���-{zp
ӹ� �̪a�/*�{,bo�A��f�ͧ����L(���Yy���IRn�|zZW��̂<.jR^�9�8���/��9��J�E�"=ԞX���g�4��O��	�Cr��t�=M�*K�\�I�6/�����r�Yc�B�)0]��e��M�	�p�7Y�eA
˕7�%�Ud9@��鋒No+/E�����_�$*�Z@~��e��h˿7L0M�@*�HO�u��7w^�5ض���&�A<i����I��7�{����:�(�&��ﶫ�#v����P���)%�.ѩ%P~m~�\�~���ha<qԅ�~�٩��c��C����~��ɜ��������G��!2�X�u�@AX}�xf��m?�[��(X�,J=x�+��o��%u��}��	D-�3,C|�*}`�?�(P���l6[&cm����G��@=G��	�cR��� ��fpd��T�	��j��%� a�UI�$�s�^�ħ�^Q����L)� T���c��:rGC�ʞNޞ�z6�N��T#����8�u _�T��n�f4_\a���-�ۜT>����=R9� ��v�;t��/�{O1���rI�yBK��Za�JQMK���5�����Vʨ���Z3ƈG��͑�����.�ɹ�V��DT���l���d�m��^��1��:ϑ4�Ȯ��|ރ��u��t����x�W}F���/[��2s���K�s��&���DQ,$:�q�Q��XӴ�H=��b��1g%�&���y��t:d.�g.>��&����(�yr��02��DOm����?�#�P������M��D��IL�@Y����q�0���۾�d]8e.cC��Msc4�T�L��o-g��b��yɕL�k9�2
�+����g���Ֆ^�A"��	<A���2�:S�wk��~���#�0D�%V����6);����!q�3�@A"~c�l�$�z��B��T���e��Mm�"�l����0�9�FU�Qj� �0]�IdOE2򍏝���(���x_�a�txn�����,�5�\G��T�35��qH��AJ#��'�UZC�2d_r�{f��o7�_�਻p�8��1W�����֤T\�j��Y��\.X�R�e�a	Ⱥ��kR��;#�H<��*�Y"{M-7��m˷���p#�K|p�}0�i���L�W���Y�M��'|i���/0�[E�!���=N��C#{�����z�.��D���xy��7^�q���ۥ�_+)|�몉�k�?�.�&���_�o���ӔC�K:]RT7�1���@�	�F��ႆ�r^7$'e����O��j&�
L���#�xv�I��"���1�Mn6�ʸ�?{Vs��aM�i���ǪV����e�����+�PRƥ�P�d�O��+ 7��󜞺RM�'ꬭ�Ҟ�C����
ꋎeA��1��{�[}`'�ŠuNdN�h�\��Q�~�I���Vuͣ���ҕ�g�j<�XN��]�����|�t�!8߁X�:Q�1���f�g��_lc���c�J�AE�>l�"���'��M� _�6�J֘�RoC`���l���8r% W�1��-B>1��k�ᘠA-,��܁�k<2vUR#?�a+�����U�/]�?�@�]H6^�U�1Ew�G�0�Lj��TVX�eE���$����h��(&���crn7���N̓�����Zپ���~H3�hb^���ٻ�-����i �S����9W_�N�����lS�^�<�z�{V��
�`b�6+.����]�A	ᓶ�>���r�S�7�ήc���� �'��n پ�Δ��Pf�*Cuǣ�1ਿ3�y�/�ż��5�z�+X�G����p5f��Ύ���������q�<���&���V����R}�� �����;����q���*���k��I���ϣ9�9	r�@#�z�+3^쟀��چ�����'�O:į��A�L�~gyN�#|�b����%y8�?a��������O�xu�,
E�/�#Kڳ2����0P��n|rR�{����*�KX?��^h��)��#@;k:m�fL�d���ĩ��=_��d��g�V�(�T`Ϥ'q����42��g�cw�rbGv�\:g��@�'f�Zz��
�Am��	����T���E�(x)y�߼�+��#��!/(�ft�>������D���c�Q���X��)m�`��RJ�ʬD�9";�? ��Z/\g�BOr��`�wH�X	�@��Om�\����Ƥ�N���\&��aa�K��=��А�9���Oּ^��L<VOW����rj)�R�@�3T��nih�����,�f������,��ƃ�#�(�g7~��&'����+�^>E�C�?��y�#l.���k����:�Es&ZF �<���r���驛^�^���� ��k��w�Q{䥈*2����W)78����`2̇�o���[�^w�E��pƙ�5�(�M7"<h�lnr�ߢ�%���;��J�4yǈ�ѳQ<:p<�z6�ÊVa��-�^^�6vQ��7[Z�k��d�!>5��-C�b6/&p��S�Fٜ?����h��Ib4�;a:l��L�.�Zl4����G��nxI��P�4��d��ʛO�i������.�&xF��)���a�����i���`�0���_51G���sG�%�vn(���2��w�	i:[�C�ۢ��f�g��S0[4b������^�0�a�B\)�w�����H>UN��R��)�68���槈��Ʒ���r`�l ���:���u ��OT�O�}~=8���T�n��O�b��Ҋє���Ѿ��, �	aV/�	�)k)�]̥$�H��5i�Ȑ�4˸~�W��%E���0��17�0��Ϊ��Є P�3H��z�d����]��sp��>���E���SC�~�O����9�ڜ���L9����� &��t}���d�PP��h�\�A�_/>]�|p�*MA �.�[΢�h���#������^'����;Q�RGy�_MZ'�/�/8�\��&���Na"&19�!9�>��r�VMܟ�+�!Oo�":�t3��~�E�6�hZ���#���,��;� j��`%9Sy�����[� T��g�� 3Y���/�L�,��_��sD(sC�_�43%��J�aK6�uUd+�	u���}���o�-�:�Q�X��B�q,�K�xO�*�:\6��8y�Ǧhr���c%�cQ�5�kɤ�b��'��X���2���7���c�����f�L
�^�&�>��S��c���&�*��'<�UH!��S�MJ=(��:��,c�yHj�F;� /�fs��)&䬟��}�N--o��xr��h�J�f�z�9kt3�.j�l{O�n���H����Guk+��3ȇ�uý ���2���YK_���eN��������V��N�2Z��T]ͻR�ơEٮ*�'�t�r�bH�G}�ꤓ�5	�[!�z��m}|O6m��g���T#�&xs���01��.��i�2�ľ���h���a��������&_� s�.����K��>�~"N`g�@0�=Q3��{ d���.T7����DQ�׼�bp-C�a�ڽ@h������\��ò��3��G��Q�h�l����Z�3������F(/f��M$�k�,�Qȗ�a�Y�W⫰K��q@�NƏ�
(}g6��[䗩����|�CAvӗ �cdo�H(lO�-LK�JԠ�-�geԗ5�����c ��t����c���em����z���oԝ�k�9�����e	�����^������(��PUV���=u�2�I$�ɷE깿�[�Q�C�&
&K�9[&&/7;ǫ�/�v����]�p' &� &�{����F�:�E��'��+�t�Ό�;̣����-�|��/�xIſ��@'딶U�)���$��<^���Ϊ���VC!|�SYR3��*�ȹprK�J�!^��-��C�w�8r�|����ϟ�܊�����Px��$���ǜ���|�O��s�$��S���W*����V#���-X��3nc�b4�m�m�}Y���ι_����b�>�o^%���� a˿菛"8����u��ᗿs�[م�����	���94��A`񟺁�WMx�/B=Uz}M��)�&�����Fi[�*x�������N��#x��:�g���:�@{����!��2*#�:�SC�A�	�!�sVXc�&jj���_z0_�Tщ�4�>��$��Kف�b��5K��,�X,�6y�0xc�Bbz\$�H�Y;�d��İ�tcLy!W����hP����֏k��0͋D��H��_(��
���@(��Xg4;�.癓F�6�of�=��1���N���6�®�r]8m��p��BwhD��k�\?]����(tL ���݄2��Ҽ�;"��4-7�834OjY�{ͲI��؇�Z��L����۲_�fX���ɮr>�B�'�~N�8ѻ���=�3��i:N�F$�H���rKpe$���yx&Ԃ�~ ;_�Zw�D;pIU`�8=s����ڈ��_)%:�ΰ�b�mi��Q��l*��\K���h*�]�nJ�H/tjx�YEƀ���s��JpI�1�Hͦ!���Z��X7e֯Uj���X�;�58�-]�ѐ3I�a
OL��=�#�Kv\R�:(ڲ���?���B�����S�"?�мӈ�wN΄���c��f��mCZ~�Voc~|�FMh��Ķ�>��0F ��&i��R_�#��p�-���U������M�[�V�^\�nX6�}<#�2(�2�^�l�ޑ��h�P>��
��hL��	krUP���)�?��g�Ӝ�b�Zc�%14��}$�U�3K��uB��
����S��� ���&Rq�C�$�G�U�1��RpEZ�>&۾����'���=W88I�+	��=�5�h( N���"h�T��<+/^����b��q�7���$&A1����_�E+�S Po,~.	��_1�i4k�a�lV����T�ކ��M�{^.31	�������(�F�߀N�ԧ���
�Z@-�/����>�D�g�z0Z���>��|��̴�H'S'�c�a�8o��u(��/�eX|�7xy�c���N�1IZ�@oe:�m�_&���D3͜���hC�H��|���{:�?�MzaV�Ci��7~𳝢IZ�d�{;?�2
���w��5��A**ةN�FT�f_W��t�����ӊ[�o��ߴ�LMen �4�ۆ3�E�7A��p2\�(���^(0kv�G"��HߖݽfK�4�V~\.CϱE���'�ҧf�|"z46$ܺ����_Y�v�3����
��P�a1����6���I\c-����y��R���w7��do��E�01���ǣ�1�#[A�VO&���R�|������"�jO�CM�*��W�[h�4b�nZmP��(�=���X���N���]_���x<�i.J��U��
�bNS��m�@�C�1@MB�c�C��mg�D:[P��5P��`�ƭ��8O�j0�;�[��<(;v�Ә��.��� ~�٧	��f�nM�UG��������`��&0h������:6�V��R[�1��[�*��첨�N,�����Ƒݫ^��3��#�l=�w�%ũ�������kwR�_�E%0O�A������OR�d��;�z^vj]wy�P�x�T�US��d�FPlI�ǔ�E�s������@ %ʹ!Z���l{�e��7/~�ѭ�(7��6.Ez�j��Q���#	�p�K�ߓ0hb&Q�d�_������7%�*%�sȔ�r���.d���@�L�䜰�"(�A����<��$�v6�^�[L�v:���譼�/Y��aGc��`zH%���'g*3�����ƥ6��W�]�5�^��kj[x軜砫�˾��#��-�U�������~/�}ݫ�h2�X���Ѱ +���i�� �6Ni�caָ�Su����6���x�y�o�B�"���j�q�T�/�q�E�o��1�I>�v!�����^�F}/>����'?u+�X�X�sW���;��0��׭��yi&T�D�Ѹ���Jv 9<�܆��z�P�n���ߍ��J� uG��}[(��h�E@��ӥ�l��f�2�xс.Ӊ�t���Ò(*!9߉E���ie�B�y!��*����^u�����`���l�S�3r��8���xf�c+,�����av���j*�}��3}�r��Gc�����i�%�*���[c�s=�
�*�u�=�����X��T��͋��̞ǃv����>M8S�Rי���Z�ΘЀ7�.[tq���ҧ|a0��,ܑ�[��D�K�E�KxC�Unxf<�Ս��LA���5��<�6?��{$;S��o�q"�*�^��P��5�ݑn�@�g�lm{D�d�
�:R˅�V>�����ȏ�ݶ+ 6`�(.}>�+�_[�Ř�֛p���� g�͸<��K��t����8�~�T2AAU2LWJ�;�=��cg
D��b&`^*�WH�Xm:��Ag��ڡeZ��D��u�fr��.����7[!@L�M����m�H�{���S��6g��a�b�>#xTb�\b��!{���(�J{��(�ܝ�c%W�ǡ)%��B}w������� ��@��'˯�l���P��T�˱6���6�
̓��A�Q�5�,+��b�"TL{�m�1�)�jQ��v%��O�K��]8��?�?�� ��A�-;SC7�M��mXW|�·4�;������@@�qҾ\"J�3F�8�Kڗ{̔02��$:�<�ͅb%����ޫ�8l+�u)8,	ĲY�pm�A(�F���Mߗ嫚*Ա�����q�[P���C���(��[�ve�
��z�}x��}�[�`�'=��0ooge���=��:��_���}߄WP�u��(ތXJ*@�Uo��o�p %��;��|v�?A�jtPн��������o��� ��G�G={�uM�ҌI\{�ښ	�r�bJ1xgՅz? �Q��hO�@ ܞC���qϬ�_V�m���1�K�k$&���\�4�
H@@�����X�T���)�56����+�e��s��L����#��"Ӥ+���sv� ��`#�?Qh9�I�j��T�~�J�@&��x�6������A�uL��N&��%8��q&��:���~ۄY��q�N@2��v�7vf�Z���j ��ś����=�	YQ�M�J��݊a>E=Ѝ�p�?<��,|�kvs+{��@[�D6Ψ"���:�'AG
',Z�m���&ZT���*��}�-����<�x��-*�VƵ��}�_(KCZ�N}���&�Ri��B��m����/Sׇ
��'!���}�6�^9H�qw�	Gh�9c��Y�sd���N�d��b	�@f��x|t�@ڸ*�
i��%��;nN�k���B9��A��C7�t��c�v&�����v��MC�R�nធ��Ci_5W�JF���0��=�+a�AZ��H-�*
W��H��1���3�@.�:tn�V*>'? |b���hx|3kmٺu'�0��M4)�8cU��X�^\I;ݷŒ�p��ahV0�ug�t˦<v&B��^���(������r=��N�(x�\�4:x�C\2&���o�KO
ux��[����a��O-߲{��l�]�?�"s�3e�Ca�D\�cJaaS{mB3����MFƗ+;�M�
�E�0���,�A�D� \S�9���Ϋ�9�]�� �\�ز5_{����X�Hy���{Дhi1���\�p�?}�_ZD���t��"k=�$:��i�v:�OX�Y��>٠����)�g?�QoV��; V����^X�eԈ�V[#���/�PC�4}t���8�6���\\R\��_+g���tC�o}L�wU�w���LS"�P)�c�X�
��Z�f��V� n���:Ix��Oͬ��e���H�#U�_XO����߿��o�g�Sڿc�?x��N���Ć}�\�c��$5���^yMj��M!��a�YO�THa�1V�ͱ�Q��!�&�&�����[:���i� n����h�V���\!)Kb�k8J����޷`�tdH�Y<��m�Ő�.��&e��!��h���Kt	o-��~�f��}�	s�}�lEL �d�Y��@��ؽ/���E�����卦��3�%�h�!�ى�Ğ���o��m�K�w�Uns�QI�����.ic����"w\���d�l"���In?"Q���F˖|�P&�D
��D�	�Oe���;���j����;��EkL���I�n���`��V x7�8^T�z59�bmxf�ofVQ	�E�(̎}����u"�x�?�7q���Lz^1��g�Ɏҏ��TCQ�D׸�W��$�Z~�Q���z�b�_j�b0�0��z�r�����E��|5�i�����nm*�{(!��	�.�������Llo3�wx,�3��!-9������W;F���8W�.롩Þ����2ﻣ9��c	2��Q@��n-�W�0m��-��%�.Jt#S�z��p���	�i3�Ҳ�8���X7�g>�%�K���A�u2H� �t��wY��Gۘ�_X��������¸���\u�tFÚ9�-[��_VW~=�fN��`�K�T�n#�J�w��_vl��c0���|�Q���};>�V�*���'���MWL�?����yg鐠�dd�@�G�*���ԋ�E��բQk����>y���Ha��r��o|�M�@�Yb�l�O*��P@�㡶�<��V��\w�N�`��c/�1�Q��@��6��aUcxx��6#Wי����m�~��\҇^#��M������_'e��Yo��\�aN�1���vd����G=���(�����MX��i�'d��^%�_w\����:�īD��pq ϕ��Jv/��	lW99w�u���hv�6�;$7�D��ud_��)L
��~:��+W绋�:��Ѝ~�]����HNdJOK��Z��.X�}���A�z8us�u_�o:`�͞��5���\�t��Y�֘���<�����`&6��b2�y��@��" � % ߂l��`4��3�T�Ř(Q:��1nS>�(��/�@&��b*���M+? R�:��f�����e�]?����_�46�5�╙�Kz�6����Xk�AC�B�$b�x�z� A��R�C��j��_�>�-��Jэ����0�����c�(�	 z�&p�n�i�ҽ��I���Q~c�����|���J=<�-"���N3%CWIP�Qz�,h4n�>���,�������Z⼻�U��Zl���"�ܑ����j���wz�0/�϶|3�p���=9A��,!��B�C�9�Eꪀ(�����>�fl�^��N�3!S���M��)H�[���V�S:�����Z��H����")��^��`,/"�@��l�;����Ľ�/��G1U�;uH�����z|�0��kэ���>~����@�~���gQ��bl�0[��_7�������*(;;N���c�rw��ޚ3$�r�^�C��AK���n���S��uD� &�郣,�`��u8��^&��dڻQVѓHMhz�A��&_ZB"�}�kI�k����_�V���I!j���ϟً���3r;Nqg{��6꺭�,��>vupOU�r��sW��#��c��S�ho��9�
I��Hy�܄��6��t`{��OTC�X�Q��0�Py[è7C�����~���N*��X������MӼ-��6c�5g!wKC6s�T�X袒t���Xn�;�~��6��y��J���.��VY�ܰ�ݶN���u 1���Gb�72`�<KC�� �u�Ch��T�{F�H�+�2��U�~ւ����T4@B��g��B�I����1`�Z�X.���ш�;����^p>����"���A��0����U�x1j�Z�3�$I3*/FF�Ьp�D_�j̠7�ڧht�U�t�~�iE�d�xW������:TŸ��ዲ}��1�v����u��|yÆ����c���Mx��#���a�y:���&����K/�@��� &Ov#"oK*�J��-��c[e� ߎC� ����Rχ�`*�i�L?Kv������Э����){��d��:T���f��;������i����$6j�����{��=Ka���l����a�;��w~�,��U��(������R6�]���x�}�S��Q��D[W�J��;�X
+�z�Pӣ�~�[2._���ǖ]� S\_�ț�V�U>E»�=D;��1��F@e�h2���囟���9@m�T��q�[�h�x� �\�f�c!�O��3�r���Hi_2��q(��_��֫��"rH�޳���I�A�W��m6�|��#���t.�5��"�8���!)�ý�̞�,���D���{s��WU����wS<ܶ���Ob4_ r�``�����):���O^�ޡ����l��9�T[�klr�Љ,o�P��qra��Nb�v�t�����Ɨ�������n�!� �΁�'Krc�(A��z�Y�g���:f�/U�8��[�6۲-�QN���si��
|j��i%�kS�֌�x��%H�i��s~�E�:
<��c�jBr�[|�U~���0W�܏^���Yg��U��Q}e�3.�wzd �$���������A~��Bd�,F|1��=Ĺ�>��X���3�l�Kx�����n'�b�ǿ(�hU���ؕ�̑� �O�i���=����PGP�P���ق������;���0������_7 9GMyP����e��~�t�]|G$^����&d��S�h
�JN0AQ����9���fh��>f�[mm���pw2�9��4���4#;�l��6іj�.v'Ԍ�����O�&�Z���H��~����q-�jw�{�A4ɂG0�K���$�؂{Bj�Tv��]�w�?"�����cI?�=bۗAJPao6Ƴ-8����A�,�6A�)_���
��/�f�l�V�.�fy��]5&!���_A�y�^kŠ~J	�,O>J8�(d=ħ���j��5�f�.AbSr�,��l���O6���e�\��~)��T-�f'O�s��@i��x�[)7��S�p�R:q�_{��0ʔ�~�$_<+_�7�h�Yt�����Ǟ�|�?Wp�������[�U6����=ֹ�\-������=��O�S��a�b���k��`KY׼<���!�=d� IUy/��Fh[�j��X�E�C�o�Y0_�R������
�J�3F��?N�
AM��-���#��(�7f���t�N:-ʯƃ
J���~��O�Α@�EX�~�3@Њg�[�����|�_���Y�3tN@��M��9�_�r��p�`�ZTm�mT�^�5�B��!$���Ѿ/��iG�C���S:�������^���N$�~��z�u��˝��)�`��{��=���D�5�B��-[J����i�g�BS������U�~��6
Ի��6�*O��`��I�M�A�X!��Em��KD}W�V^�lΕ��gb����}�p�R�<b�f���=W�7���?�K��� T:
	�c�u8{��.iB��#m/�\����J|�Q��!r^�](H�(r��8J!�'�suӺ���ex��i���s�Z��$�y��z�h����'^)��@³�Z��J��2��	|�����l�o��@>x�veJ�#1�ֆ�v��X�j��e.�`�K6��n[���P�:����?��#�3��+�[n��>��߱0yL
��@� F ��>�"E��k8+Ӻ_ӬGr��4�{'U�i�v�eKD�՛�Q�kId�ٺ�0�I�=o�l�Z��=��I>��XuiY�"*`f�6s%��'�{G��ANO�"p���b��mZ�[�����x;�(w*�!l׻�<���ҁWP߶�Z��a�Z����]��s+�2��e�f�ܮ�l#xt�yرÁ/+Ӂj0しμMD�o�\,����Ʀ/# 5�����4@�x��M��t6�����gG���o8��+�<2��~KY ����.
���}��,G�e��x�v��16M��fO�#��"���~B&��9���Ȉ�G|����@;
�!�~��?g]���:�ѿ1�u���7"��ɅM��*F������p¡�(A���e�[+z�<b�|��1a*˛&��M��l�裕����^<�rHt­���hZ�쨒��t�̪ZDϣ3C���*|s�+`��+-���O���ڛ�mQ��V{ 9Z��˘�(Rr����9aP�eaqZ�eL�����/�B D���F���B�%�Ң/k#��
�N��Gb��ƽs��(-�it�;C>��>�v�_���#J��$e��u��l�	��Tʶ��`��d��?��l�<���d�OV,B��f+�uz8��c,�ynՌ��/�A���h��9��^�'��(��|��rhX�:� �O�{���1���L�)�ă���FnX���6a��M"|،��:�'S;�BOG�(���K"���I��6`��eo�Vm�jܥ��
9N�1Mg���k9��j��'��	�gkV���9a�N7bZSf�d����2���J�#�d���v���� �[��~����Q����0`����:
�����BJHg�t���-.�_.���
|�֬`O�����"r��������@�D�7���Y�[|�7}NE����Q��l����k��^'����*a���y^�._�BU<*��Ո��#�;}*��qq�����ma�'�]���0��߈_��|�.zgj�Fh�P�s,�����t\�@F�RB��"�cq?Y�L���*�eRG��=��[:��M$�[��>������3����� K�y���$��eǾ۠kTg2��R��>� $fS%u�VL}-;e��b��{��
�	�&��Xx�s�K6�K�M=z� �ZN�ȭQ��o3��1��z���q���xoj�r'n P��uJ*l�v�.���	�&��2V��F�����k�G���9N���d)���ȃ���V�c�$�o���!'>��!�K�YJJa]�qoEE\N?Xh�Br�Ch�7��F�#�a�{%f��sW�\�}	&�Ǻ�ix��P���� K��t����zWsA{I kq��t�Z\>a0U�+:u�g�X�w�O�5C�w�ڭ�N !=��/j ���̕��8������s���ro�vs��Hď^/�k� y�|B�v>w�֮x����k���sHr�+Nt]�B1;�[�F��D�5� ��w�.<5�;Ȁ^�O�Z_!�=�%��w�d%�E���o������W��e"Uw@^�1�PN��`wZg�S2�2`�/�nx=���b�n�X�k��r��b��_�I$Fw�[�q��O��f*�G�]�r��2ȷs�l�-��FM�Џ��� Y�-C��g�B�����$D�R��KIE���=�g}�
@= i�Zn��Q-5�+���2&��/��e����,=i�QMY뙻����<����Ȱ�<�����:�͵!���%��2^��ۛН?�.��_Lc�rK؆�;��i��������[�~^�|IY���k�x��Jh�gЮ���b�(,L�S,�U�.����Q�6�k�p=�:e�d	hPK��F!�_	 �E�3j�?N�}q�j0v�Fp��K�r!1vl+�D�IV�R���i��P�P,ݧ�u�Hѵ�W�n�eŌ���]ɽ�5��ÛC+��ǝ�1|���FEݳ����b�.h�C��P!Y߮���u�5��x�-�+���m��(��{BS�dʢI��j؃�(�iN��v\8nB9�I8n�NvN:��]�AH~ڸI�L�!W�Q�B�c&[���'HPJhm���N�*�vF\�9�����m�t�E'�Q-�c��sW'�QSɱ7&m�{ʟ͇�:u�&Fg��r{��Ao�ވ���پ�11t�lc�2�רiK��ݲL/��P��$4,�^�5h1l� ��T��C{�_��-��_g&��=|\I��=f�E��O��Z�j^LпJ��_@ � *r�N(o�rk-�+��2��o5p*#��Ǘ��^�[�F�#�:aD�2�X|�b@�5�#J��?"� ��$��w�/��� �4X���
���<湏�j���;My���ؖ�- �x����G�͘b\?|f�e	KMd�$���F[��'�G����'.��@�+aQ�!�8���h-��jǯ�j�P�����A��y���[a��Iٔ��S��$j�L\7K6C�0u+}k�����*q�$ָ�b�Y�����/��ߛy�Ջ�HU���|m*o$�\�QkJ\j����I^)�ʄ]��X⏏�n�`v�m<�ʨ��~������<[�[ƓX������T�|�(�H�}��w�wk�M+u��IQ�Ys��X���"�wC���@�&��#�_�K	���s 8ŏ�;��Y��X�v"c�����:�o4-4�6���5�����LtS����x���<C�w6�8,	�Y�\V���P�Y�'��V��*{��R(�v�i����3T��X�*��>p��b%M��bǺ�l�g���ӭBЧ��K�y,'Q7��xX=�*�ϕbL'@��/(�i-e����<uޢ��z����ƴ;�n�4�M�U�~5P
"G@3����l�@�o���Uu���Hk��$Ґ�◨�~��(�U��a���j�G��j�u�R	�E<���_��P;�ҡT��dAWB�R�~�GJ���sy����hI�l�+Y��@r���oD��X��+�@R�o��K5��]^B�|���8��$�W��W�;��~~�����C�nx���㴀I<G��ꄰ�ޢ:\��'^�� ���h�N��(	Bf�A��q"S�j3!p�$J�cW$��;w�*��Z|�s4��2��쑹��snR|QG�MG��0�}���+� �00/X�=coB�@�A�Q�Lr��+����0-�Fj�>�����A��ˌF
�v%���A����:��!��z���RX�ST��Y���S* ����Cn!ThQV��Ģ��$�8��.�LI䊀�r��,yD~��HQ�~�v���!X�m龜��'�r�N���B����,Wa������4b��&}d�8 16�&#g~ڧr+���ݔz���h�.�yiЈ�?D�hQ�����>�e��c�|H����c�8>��O��|���B�(�b��`#Ō"d�X��r� l��8�́��������Y�?1.1];����q�j��~Ĝ/v�!5����Y�o)�>��z^�/9�K�X��pWE���7%�b���[��XqK���7�pĖc�"'�I��D���OA�Z���u��qI����l��
�fEѴ��%)�K����|v�m�Nɠ�w��-�֊ ϩ��7��U�ѿg�[q(܈nhk�%�%��d�ϴm[��1̩��=�Þ-/��v;1ZK{8��y;Wؔ���a�m4��!�ıY�x�|������Kh��\Ӓ�m��� NL�ק�˛� ���s2�E)�������q���MKO�<�]�|�w�?5�m��Dt�vi؈��"ex����aLrY���஄���>�'�K7����r|@��D9;�u��	���z��:�؃U�]An�,�j��<�n,S8�H�s��gX��X	|� ��Մ�t���5\j��i�н�?�\���l7[�,�MЉ����ի�R��7Me�qrD��AoD,"<8�+s8#3ɚ_^X�x�]��pЃC_ԥ����?QP:�)�$y�M*�܏TpIǩ�(*7u2���.yQF�ܫ�r�J�-36�5�k���R՞�����1Pq;+/�#D���K�ߐ�6dD��Z��{\��/��#���\M��1���{>�"Q�Ȟ[���]�&��ԋQ��rћ�h�J�b���Q6�9a��AE��������z��h6���T���%"��j\T8n�"!8ŪD̛A�ٌݴ,>�Ĝ`e/�ӻ��|I:�	hG�;�U�΀8��<؜M���}fj�D$��^T�$���I�E�;s[GT�ݘ����j�Qv�qYe�,ڳ��x0�*ק���MS�w�����I��N]�Z�@h���|��!���~��Z���nC;'�oD��%�/[���}CkZ:,�d�
ȉ���O��H��Un�B�J"��(SP�hj��$oc���*v[@t��[&��.����=8�WY�	�,�|��:�"35YGY��N�b�֕q���J�p�j�C��,�!�<����ԥ7ަ�U�8�r��ʨ�.���#��������h���eL��U>���b	ﰁ]B>��#�������f�����6���Y�ܲwk�oP�(��cZiB��,us�I��������%5���-��#hB}޸���
��Pw��EN-�w�N�g��{p��d7L���TgmPM�Y�K�L���OS�'��k�� ݟe��׽~�� ��Jq�r!�3U�W$��[b�j�����{!�@>P�Q�7�vw�+�n#~��n(�RA���߆D9Ƣ�iv0��	�syp��=B!��0���� [!���PW���,bQ�>�f6K;��q�5O�?V+�ZϪ^��b*��,�[֞���s��U�ic���k�,�"`:>?�lȢ��K���_��j�X2P����XЩ��Wda��g�a��[Ç�jJS(�5���[�O��_r��|�:����UN��#9�&H��߅�Z/�r��	��P]>�>�J�؅�²�/�)_Ju�M8�^%���G><���]��W�Y+�VC������SgX���ϼ3m�:I@���6��Nm>�
_r:���lj,�W�/�Fy�β.VO�>\�V�3�|gD&K���$�q���u"ԅ�%q@�馃մ8P��/�E�׷�SG����\W�K���C��Yg��ZdA��M.g+O0� �G�<<"H����?���N��rs����\���Nd�X�J=l3�W��GG?�n��/�O\��/8�_����.ggvߛc�4�4u,��
�W=��iRdT��K ���,���e��rv�R�{جK�h$����˳�����+��c�?aDUa�'�9~�e<Ӱ��4	���˸ 9����MYΒ����eji܅D��y��8���x&��v޲�����P�[��^�NH�I�(��)��->n�7��xg��ߍ i��	
+�2��T���e���$v�+a�[��_ʞ0���_8����K)��~hoVF�+9����ո�w����j���%�v��߀���tci�'�q>cյ��H��3�[��=�Z�觞C����#͸�*~�����<��SKܸ�V�P��^J	� ]������=��
���6a��nz6��ȆS������,�>���i���_�	Ml���A��qAr<4����F�vH�I��x����G���<��BЊc�Q��{.T����hcH��8�s�!�,��a���7��|���=�0BR{V�^�cxԠۍ�hFyK�P}�s'3��hZq�L	Om� ��:�dV�?{���.���?Z�]�l���V/�9�KZd�s�L�\˔��sY�Y��y-�X9#���_s}H5-���L=�@M{~�hz�j��"�ţ���9t��+_{��Q�
xa�����h�3�����E#���U'����4�+E��ڢzk�����^��.73^�pY�u`YA��!�se�<�^IA.8�a�~������=�ۀ�����dR�<��P,7���O�D��H5��\��s����R���w��yp�h��� )7)R���o%��d��n���ToO"��-ضZ���E�m�5��#V���X
E���d��k��#5����[#�7���a2���=X��#x���MҜ�O�$�\e���+Y�m�U<��º�����������m�B���3tkY������k���y��-�߉~��"�Dvh�bi�4/�l䔧�Sh<�����ְ��Ps�h�3��D�>�w�_2����K��2��]�-ǵL��BZ�����=��z�&�����?�X_g�Y�7��Y����8
�H"ݖ�1^��v�F���hw���6j�r֚�x��-f�S��K�/r��F���*�%"���<@$�UG�.�q�F�R�O��<���t��7(�iZ��%��PQ� a� c��Iv$J��
Fx`zD9��m�'Ԑ��+�i����=W1W���jGw�����`����5��#	Dc ���I�����V��֟�t����y�TF:1��X���A=��=lA��'���M��N����1�I����t6�=��\@�өQ*R0����Y��Y��8�4�:Z~*�tLJf���� �f�w�p�Eɺ_�j ���@OJ��ݍt�׋z��.h��r~.��~yEy���b��ڌD��?�X̡^Z��f^��9v��9���r�3����k�Y���:_�m��CT2cr�GeHτ>���Hq0�̳�|^Q�Y�u��/�$V##��̡���U�*F���Z�a]�6ԼF+^�Ѱo�:���K�42��/M벅$BKVF򛄿����?U�u��aՁ���Zu;JBt�#�5�Dj׀)�\O��^�iJfD�bn��T0��^�SǗo�^/i'���GG��r��sȲ��I>ŀ|�'ˈ�{+'K�	r��C���Z-ĹEE&|��"��%[w�Yh쳀�®96�4���yH�3���� ��2uPՃ��4E���^P���� �p���^h������P:$>p�bXƿr�L{�Q��I�)G���vL���9�Bz{��%������DH��k�!Z^�oV�ue�[0��AJ}5��p�ܾ�LpH��?b�5c[7u;�_�FI�q�_��u���4�P~ ��t/�4K|��٘����ٙ%ZfO��&yJ�w�Tb��l&;�1�ͅ�ߘ!%^0	«G�¶�j����mɇ�Ԇ!�6�����?�Ĥ��I%W+�ධ��,\9ۿ��6OND��gؒX{��s)M��}ބ]�}3���`�]�S�i��3b���,�
\!?�5���/�pF�캒�/����S7f�d��_�pe ���X$nV"mN��thc0t,,n�����4���i��<����˖�%��zV����b�:�A��GQeQx�lf�{.~��`��@k d��R�פOqDO�`Z �'��_��т����g���^XN_h�i���h1�؍h(>NZ?��2A��=�V�<������#B��myw7�u�j+�49p���̐Ë�L�Ԙ�fV�w�_ ����1#K�)����*�_6�l�r��`߱�*�9����5M�p�J���8+(��j�M����L�
{ k��W�z�_yVq����o�}�Oi����O�q�XR[^{�x��x���y��Hǵ���.�S��$��zK΃�bo{z
�YI����H���hgb�U,�>�p~�M~�Kt9�60l�r��
�ez/�ɮ� D�.w���v������8�Ƣx� z?�� �K��pn�k{�Ցʵ��I���_;�\!F��Ef�{06\nh�X��.�eaǉ5��&R{���l(:��c�Zy(�;����J���tshc�`�Ik����۪tv�Xr�f(4S��Q,�h�9z�i�J��g�'�W�uqS5���� (��o_�aK��L%�Z&!��mѧ4`����<K�0j���#������CԤծ��s�����e'8�*�f���}V����8���JA_o^l�:-��ቧ;����-�ޏa���I��)