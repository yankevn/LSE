��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~ށ;�|
�����6,�pk�N���WIVq�湭z��O&��4� T�:J�V��t�~9u�{4�`4�]j�CO�c���5?;DX��1�����r��如ػIEI9���̾x�_]<�d�����;f�G�W}��� \s"�Y���
~vE�\t��ұ�r���ȗ%N(�
�(8�,�IJ:�1��L�I�#�!��i�l��@��T���XQ��F�}"^yug=V8�����a4w��]���܂z3��ϩ�ub�c�F�p�`���'��@.<Bo1�$��+"�E�q����snec�e��y�����|�!t�i�}xp0�.T���z.M�i�&LL ���#����b����V������<�|v�����p�\M�ʎ<�ѻ�3b��+��1�wM�['.��&]�ǋ4��-��>�	�4)���~�z
�;;� �a��e�[P�d�"ߜ����Hb��B��'��Î�`h��E�S80P�;%x�K��ŗK�m.*���g�Ak3�A$pe�<M�!9�S��͆�.N��G��������\��9}-�e�ywf	h/ڴ`(8�Mc��R�o��?���?7'�35�'TH�!$��z�}?~y�;�|)�"@f�֥T�}}nCǄ&]�	��B�c�ӵ�5ȐyNh~�XdT��{��#hī�ӊ�����"I�b������@�a��6������U���tYfQ[�T6���K���A�ٷٽ,�^.%ja��`�1:ۖԀJ.'.v�k_6�@���$��T��ߎHFC�(3�o��gD�z9�c3��q��!��63f:7��#��f��Xj�6��d�L�FPϜ�w���w�D�r�erP.fAt����n�'B��:�>F���+�����ݼ�� ¹�M1 W�>tcT]*k\9��2$���o��V<l�?��#����1��#zhd.+8��W�5c�j�Cl�>>�x3f�����t�����3vH;x����zׯ�6n�D�A�vJP���λԠ�0�����c�HC�Cb�Ao�]|����Զwk��Hk�m��_�A�ܪr�{�>iJ�+�H�YW�?N�X�싩��?�y^� #�������|q���YnnQ� �Ʊ��"�@�Y?f��.����u�����������(��؛MVzkW�\�c㗽}sC�~�}3��1�[J�� &=ˋ5b���a���D~Pfײ��V�М����.;vު�C.U:����;��H��ե����Z���{=-V�����[��Ն�P�s(�Ȥ$l�k�L��ޥ�I��h��s��#�!8:.�6~�Ѯi���[\�-�o������ 	U�J���*�����&Y
�c\��P�3�B��נ������0��'n�囫�=�.v2Z����fgԲ��/�/���������Z43i�xH�{��T�A�5'�P��Y5܁ �R��ב�VR�2�\���#CqM�r1�׆2��8�W�,!�����	�R�In`h�^ �S	�kdrYbc�5�ٟ�G�Ā �(�4�:������o�H��/�bϻ��K�qb7���S�Z��8봐����T�x��:>�##Q���e"Wo�vJpĮ� ��7fũ�Xs�P�9Y��V<���JZ4���ր7�}�#xu[c�s�RP@ۉ���}|;���.�����e#uo5~��v���8AǗW}�[_*��&b��O��+Q.#@�!*�4m"nʑ�gO�蝅��v\J�����
 ��>4�6��Y�5�Ἱ��z�)>c�q���,�/�AJ=<��U�h��X&����/-�R')�ٞ5����V��u
�Đ����M�`c�S$rj�b�1��Q��i�ޔm��6&�#��?�#��&�A�iڅ�4�R�A�׳��Ւ��3j�[�[����N���Лz?������T�a�	Ӓ��g� ܒ#q��e���G_�{�@&Ü��I}�H@��X,�!��O�M�i6U(��L��g�q萬"��J��+1�$Ue\���am8�#n6Խ`�*�����L�r-��`�dY@�x� ����Mj��6[3Uap4܍��n�;����LȊ=<�U0��%ߗK 8��V���R=��+د����K!v۽Ơ'���`�I�%��[:������5���?���������|:�hWf�3��D��I�*��Y��������4)C^�e�pb���4F���a�1��bq�𴇑>����g�����4dH=��+�q[��-рdķ;%�p�0�dG2c�s�����qW��@�����$BP��w��ן:^r�%V_�a�-�E$����Y����;����)�:t.N�I�aF��W4��eXO�<�R��Ͳ�\5P�r@��?#��M����B��Q� 8\��]�E��mܺ�a�{����3��l��c��M�|���/�ׅ�Q؟<c���[�q�3���
��LY��ZFtA��+��
�|D�0�Z×w/g���Fk-\�{�[L�0~��҈t�G2.�e�Y��ـ@c�)"|V
+�u��e����f��� '��R����YQ�܆�f5��[�Ƥi�eY>�~t?��_l�̜̒v�̩��O�g3�����4�J�"��Ϡ������0˫r�� �Y@�fP�W����� �	�;c�p��ɜ_��94�C�P�Ti���/�a/��;fRy�ܼ<DiB�[���գ$��i��h}S(�UQ/s�_�}�S��h��"�h��<ϼ �� �H�J,f�;�ԷQS\��(�f�$>�3��������+�f=4��"�a��0
�vH���>��DY�)q�T�3_���Ʃ� 1[;T��A36��\��)fgY�C��
DR����eA��G��߄���m�H[��T_��O�&y�-�R�iILv������oޖ5�e~A�o���@f�0�\T�߯e���Ɋ�P5�ٿ��I�ý���8�^��)��k�f-o]F=Bg�9]bO��8�ZF���#p��t��r�}~%��K9_K�SD�QML���U��ɭۥM������H���AK[w���������O7�� �Z���'k�~Z�pj�Z0�o9L��$�l�Ζ@YaB����>t�"�^� �Crh��g^EX��99|���?��G�4 ���\ ��"v���sa��CS<m�>��/�i��CR	5�{p����W0P�v��+Q���D)AI3�+�]��:�̾}�@K�v��W�I�o[>���'��jQ��;���&�˔���N�`�Z?������dl�[�x*�2�5toӂ�=�(l K=�G��zsl���P�������َ� f�4�,eW��~����������k�D���Tw�zH��.64���{eV�c�{Tm4As
�;Is�au�<�+���J�ҙ�i�W��ӊ��gdһX�^�Pe�3�3�vtҼ��d��2S+a�e]���?b���)� QF,�U?{W�$R�Ȕ5|
���7�+��c�_i�\�ek�d��僕���M��I��BїE&ϒ,ъ~o���P�%q�͸fH�[xI<j�*�L�
���`�Rs�d胳�H�/DO�ț�$�� �Ÿ�7���|d�E�m��~Ԣ��;�?hE/�VA�%�E�=l�4���;��K*���1D5��Bв[�\W"�=���4Ml�LuE�`]v�(wJ��X�¢F	���4�
�e|�['A�%��<#Y�zG���� 29�}�dmNqnC��} [d�S_a�Z�
��s5���R׻POZ}��j�ץ�hl;=�$"C��~�|�Gj�Ð���Ku�ðm��CCa����ш�d��u^Dq��{7��|�#�ݼ	E�/Tt�*��iO��^#sB~��笃"t��a��i��'Q~�p^�+p��V��e�tV�k������/%o��<����z	 �:�ȑ��T��v
'�.h�IJ� 32	�C�C��l���-��i|kg�����<T�S��'l" �*��gs;�7i
��D��NIkRv�X�jž�6S�H?TOTG�{s|9ǜ��0%�\�]�L �N��}�=9,�$>���?���Q�@�f�R�c�06�+�E�~�]���o}��>�Au��{U�����n�;8a��ȥ�̛�/+��8\�.�>s������ٟ�}�
+�����tc=��)f��:��-c9�[z����:�!XAS��_%ü�03h`p�3�K�䶶�����	wяy��FR{��\M��e$��/# 
�� �@��Nd�"�H��_?
�F�D�D�-��N_�B�j1_,	ؓ����݋a�}\tA��g3��Έ=�Wor��'�3��@E/E�l��_������O�-��������	�ĺ���YKy<�2�~�������)�A:��� v^�`��V�=s��R�	L\���֑;.?GUB���iP�~����]���B$L�������]%kh�C��[��\�@]��x$�ߝ�r�t�3�i�2GY��P��y�	+�x��Q�?M!h�� :��p-���H��A���E�P��
ENIy��QSr�p��OgԞ��*oBh��$��@1� �Xubª��򽙎Q	<(&F�G���Ock�S^U�*Ĕ�<��8\�����&���LI�3)��sG��"/�z@2A��[<�ە��+�U	��'�x+�\���W��(��	�w2%���C�m�N��ށ�*���ow+���>c��e(��#w_2���Mn!���9���ξ�>s�����JoG����6��f�@[(�Ke5M�]����YHc1G���@�P�x�z8��g�+TzK�4��H[�7����aQ���n��C�1��{Q����+@�Jpd��;3h�ġ��K�o��87��&D�k��$�ː�u��Ȧqh���h���|�xo~�6�31��-�uW�*F�mI%�I���yH����=�[�n���X��8���bɧ�H���ު0D�xC�"�7�x���L	�9U��c���Oe][.��*��?�(���6E������6S��.F��+�FP�rZs�[�=�Ev����+�qR��x����#�x�v��n#�:���N���}�K-����m&�p�u���j�IK |��<Z��ު�3m�rdlh,V�x��@�-����oכvw�6��?Qa�Y(Y�?c���3���Z���<�����S�;!���TW]�'1��hoS3�m�7�3���Td��6�o���嗩��WM�%�v F�m��Sƀ'����]�2�OL֦���gB|kq�9ɓU���(�)u��G=��ow��wP�?�"!��,�f[����ṡ:��y�l�/Kx5*��s�߮�������� �ldn ��>J;~���j-�>+�b$ʹj�S��T�A;ޕJs�F\f��{~؆�J�~�.X;,ܥho��7��v?(�8T�޶c7���=��eS������ U�����0�V(�A�"|J�u!�w5�<��Q~�V�
y��]��qjߨ>s��{Hn��ߐ x�+
d�^=�*�׏�u��x�oa���j�U��_�$�v�¢��b��%t�F���v2�I���*��AC�%%�޳�����`�]�"緒j8��yJ��쨯}��?�z�`�$���76G�P�8I�u�����˸��ags�Tg�?X	?pO�5T����*�K���Sh? �gl��9v-#?���+�b��,��qVG.�q+��6,�mi�v�@�1Bl�99y�7S�c�X䪭xB6�T�N0v����y��c78U�qnZL�q�:E(�2GSb�]�siU�X�,)�Ur� wʍ
+���Z-�Ƃ�8�*i�a+M�� ��I��9w�AS4���tڕE��;���#�>�[+�����Y=N%�;gƿy|��zP��EM6����C�R��^O4C[_��%�N�W�����lu��X��z��>��0���O�])�PE�%_�W=i��(y�4��x������QC�r)`�G���?��ɸw�6T�����|t@�[2^�RFJK:���'K�4e��/L�PAT���`�?y0����d�A�=6xa��h�^��g`*�2�}Z��e7�-��9Z��R�B:��4�,nE���π��>�#��Kx����¶��gYwu~=�g�z�քS`ٗ�E�;ܟ1(<u��cx�.��v�2�f)�+y�"�����ek�hTQ��f@���{`�d��Y�Ο<�MZj��������ժv�ƫ�_���
P}в�{�1Y�y��%�K2
h�0�=[-7>e<�~�ND�[���'��Q�1Y�O�ꗕ��9g���_�5'��~��BkE�Ag#���S.{�8�$ϧ��t -���8�%]\�v=^j�;�f��!P��Z5N.tޕ���WO�oI8�m�J���ȳ���^~UF��qr`"U\뮄}�l�\��2�L���/)Ͼ���\���ɩ�TD���Z L%�v6���C�U��xl�5�1�``�R*����TVŚ�8�#���o����3sB�sБu�)�H!��<*�j�����G�&D6�'�FG�h�����u�q�����z�Q>_��A�k��,Y����>��Y���y�o{1W��خ`�钃l�pbB�9�oz��2�K��s 9��\Ny姘�M�@� �Fą��rZ}WL���g% �?�8_m���{&��k���m�l�{��v��N�Z/fd�$�~ON	�1��!. ��C7���9�W�FZ��hq�X���B���e�I V�QZCB��V��Z�����ҺP��N��Lf�n��ͫ�eP��T���|���KM�����7��J著�A��r�\�$��[i��� � �
�8�ه�(x�/!���Y���,�k$��&�h���s��X%\̩��.y�<��t�Ffq�tu<	��7!�8$�-[z����Н=)<hB��Vw#�Id��nL&w�p���2�E��
�#�=�ta�^[�!d ���D貴
zQv�])c�;�.djc�y��'�����Y��A���ۡ�X��ʬ;>{����M��Hc�j�a
�����~��??��}��ˇ������e~$�]�Ef9�����^��U���
�a�2]5�ҵ�j3m(&'�����A=H��dU��{,߹P��R�!��׈_CD9���c����1������H�w86�'8-4��KLd@@���o���R�,�jn���_{��{��t�]WS����!1�����{�ԳiK񘰜*#�~Q�l�]_W���p��e�\��Rf�B!�����bΞ
�##�W-a��|R]B��1��߫f(d�f��[:�cZ���J�
���R�9 �k� t�f+H��l��\͒<�+�lQ��(�eo��M�l��E���������e�ᬽ������r�7~f9�N�ᐍ�[ n�$A��mkl\����1F
Q[^�J�X�v�7&߬L����]�,q;�ћ��W֋�$�n'�qG:A��eУ��J�?��	��w+���	`W0-c��	�Cx��L�t.�'cu��j,��^Fi�G�0B�Kn���@f����d�XϨ�Wcvn?�O�������T�|v�:d�ć�N�G�A9"<��w��W�PQ��Y�{���8���'xq�w��{P�I��QBh��gFk"�쥖������YHC��G�@�8̘�dHG�UI�7��.��cWJ@�i��uq��^|��{aP�=�<q-��R��P��i��NR&=d1���t�>@c���7C7~���i����'��pȥ�t�-�=7���Ϯ��b/�g�c�S���Kx�� K�\��ȥ,��^���^���Q����C����ijI��Y��K�Ժ��l�*��S���8a\�������!I�x�6��bM�u^��D�o��jz��{���J[\O���j�ZAEIU�G�zb�u� |>���/��Aqc2��3сE:}���+�2u&O�G�!�~K"��^���rc��wX�]sU�'��+�x�d�$��i�a5#�)��k�Y�?�����}%g��;zZρw�Г�gX�~m	0�`�b�a�F�.����*4��]���q�k�O�s�%��ܞ�h��9l�A/Q]\��Dٷ��v��B���I!@(X#*:J1X�º��y*s�Q���2�Ϊ�j }�?���_�=����7ʬǿ����JUtb��G%�Am������զ��1n~U��f����j�	���ʪ:�w&W�@�c��e���=._�^m��G��``p��/�+�NL6ND�모th�7Ѕ8ˡ�0ّ�-O���!u��b_�䤈u��.XRW�������K��I��_�I�9���)Y�\fj�#^>Z�oƔ��MY���خ�Lk ��'���ߡ�IL�Z}��UH�L�`"H��ɜ +�yZĠhN�����雠0VչLң��ǔB�j����Џ�^k���#N����z��w�m����<�b����O �՝�[l ��Kꂜ���/�`^׉8UW�g%!|G���w�)�8[�A�B �@�����Q��0c޴; d�$�9Y03�+��e����K��L5lgks�!�9λa�,v&rG{��7����횁�z /��w�<UGZ�t�:��hK�hcW��D*�m�ɵ�ս���ɘ�w����'y4��iRn*�&��iZ&�g9.�E@TLl�ȿ`��Q�,+2>��:2���:����*0�m�S�,-Yį���.wy/	�P���{�G���2��C0%m��t_Ϳ����^OHEnI�U�j��d��*�r&����QV���u;EÛ��K�����<�ŭC6�ęϴ(�ɇwx�\��xOFcCI��i�e%��JX���9�61��a��gQWq�dg#����>��4����^j��|G�x�B���x��cX?9�:�w3B��Eֱ�Z�Mt֦��7+�Ϣy�U=��ڗ���3�WO�F^�:-�qT��B����r?I�x��u��*q�FZN��E��bS����͘��3�np�kn��\>�H�q�gg
����7~�����V�(����E�@kLA��B(%	,S{�H[�A��d�fx� BM-�T��2��l�Y���[�]8j�p�����(�
�����U|��g�O��I�It�Y/W��10���.��2U�ZC��Z�|����� {�[=�1�;?.;ꨳ&!%�sbf�(���<�I�Ż0�1�;U�p�����H��7%�7/��Ʌ�I�V`6��{c���a�B�F�q���>���5\]���;��w�����L���p*]���G���?����$�+�.��I0@G����T��*(�ؘQCL�=�$���<�z��LӨ�b�Z�^�6���-	ޜ;�@��_0)]w�X@$K��!.�S�f�6�~�m��3=�4��?��zǿ�~4ZY�-���j0	f���f�Uc[��3J5v��Cf�\>��B��W��d��$&D�����_�1��ah*ʩlAC\U����h�?h%�5�L���o�4��?���}bn_ʆ5�Fm�F�b!,��˘�Vye��҇�U&�<u��ǁK��sW�pc���4�Mn�)�����1xV�;���8s*�N��R�.����^<:lX>��l��s	}�&,�f_+�Ǣ>�9���nl �K3
�g���\�~����di��w��K4���N��\�}��#-�n�r�Q&/��^�J�����.%m����@K��������5g�8�h��X-���aV������ABbJ�?�X�^H���'��i���Ū0=>�G�������*ن9tՔ��#~c�~�B�}�b���W��7��8b.���"��� �0t\/�����XJc�)�$g,7J^)����U��ؖ���0d!
�f9���ߕ�aWvȧ�c܊��F�[�|�kC]H�rr:�G	�b����,�;��!5G|�W}QUU����X���C��v!8�s���bkU�W5�krQN!�7�����D��1ʧ?��E� �����}�W�*&'v�΅k��EQ,<iÎ��pܽ��6=כ ]���O�� ���Pk�� ���-l8�Ӽ\����և��Z�ln$�����L�8u�?W�KZ����k/o�[�8�r��P$n0ۨ�{-����}+�m-&=�-����l݇����G�Pp�Y#�6�.�mw�<�w2@N�o����W�f��>�d�0^
���Hɉ���w! X\	7�Ж���
 �T�І� ����I�J�^�mB�s�1l�\�t�<��5�1D�{�h��?��oy>��ȩ�=�'����ADs������(l���5��q�zCU�ܷ6�[�k	��4��B	
�,¥ߠl\5��j��)�Y͖,�)Y_;���:o�s.я�I����+���̀�Y7���C�~	�H��ϰ sT�m{��8�"���9�S:g��`�-X	��(1dOQ���e`����էU�jj��bR[R �Q�7��f'��yx����5������OM����~�)��O7�`W�Z�(��]V���x�B��BR���Ɩ�{�eY���Bj
(�R4U��ϔ�FXpsgs��Z����!!K��ӶO��ѹv����h��|����߫r�W$��*:��[��18B����i���#Z
b��8c��v�u'*�=������Ξ2� 9T�&�u�����@��|�;�B�Kpm�?�}�w ��GG�?�1�'x֮n/*&�5�Kl˟4A��a$����2N�-.[��RP2q0q�e���K�@Ds���F��n0<��Wys�=L�iX���Q��.}�t�|;�"#�x6�a�^ʯ)�T�Z�w��1�Gc���mU	�0���D��~�eL�蜩_��lo�w�56;3��V^�jrR�@�F𨓶*u��?��\�"Y��"��+���$R��צ(;��F/���x?�����;��@��ce���	B�c�l���r�U�ҽ20zT��%+^��,�o�뙿g�i���B�����]��]A�\���r��b�e9���1��{�dDg>�=!��ڒ��A��߳K���Iǝ�蛒���oSC���i��3hX�����{�y2�4G�d�6_�$��fھ���M�=�HR�ϕ��ڃz��S,Eͺ���,\�';�h�������W�Ҭ�/N�q���(�A�8�,QP*�K�'���0�3W�F��Z
Z�K�N�A�;#�p����x1:����R���R3ė����.45����'���R�TD�7�f�w���|������*���9��
�4�J)�'=�lۉ�� $Pw;��Y����\dp�3��S<��x�'�]�ԥ��Jj�dBꐥ�`J{/
��jzד�>���ӣ	� ǝ�$�_v�V�A�,#���Dn0Č[��+9GE
;Q�?����wArJ�� �g��
�6]�L�}w��Ѽ]S�D��]�<�P�Rea�q���U���b�y�ث�_�5>,;3H�#|!v�������:�H�7*޹�*<E�#����~���BC$�U�r���|q�~�Nz�qdNfS�
�*�W�+�T�H:����n�GU_4{�M�ipJ���0Pa&*�!��2"�Q-�B'0�"��ݦ���
\�#�{��</���;�Uz��«AA�~�;��"ӗ�`<�g)�zk&��S�U��C�ജ�\.d�TUp��K�+��o|a1�m��{�"@��	[��:��I.�W`��U�3eZ�IV�ԯk���@E_�To���	�U%����**_j��ƎG4���,�g�$�qgc;���Y����*ᯝ�5�6<h�ۏ\z���Ε���hX�Ĺ(���K���
���	�E�M,�YO��N�-J��'~#cT�^3�[��RT��N��-i�R@`�����W��>!�����L6O)��x�XI�aZ�r�y�m��V,g�i�'�t�wn/ӆQr��2��R�O�"��r�[��;��-X�����H"��2=):� u�$z�@f,$(*��3�ٱ���_T�]5زk��Z�I����?��鄳��I�4H!�v���+�+����qX]Xn�kCl]6������q��;�����H	AC�TE� ��삌n�1� ��� 7�Xgu���{K�������1pn^��S�Q��B�Q���O�r��*5h5^�:v6n�PҐ,���[��cW�"S̍��f���IJ7�#S�郄�Hog��6��בn��r۠�	�6��Y�p���Rtz,�3u�Ժ'y�C�23�ǔ����g ������L�I�dds�����.���U$@�]l=���]�L@����c6��`!ጙ�\�	�nZi�Fa)�_c�i+
Ś�G�p��--w��]�}�`� "�qKn��%��*�y��Hk®AS���M�:� '@�w�.rU�8b+3�/L��`�OǬیǺ��C�$���T�:�w���@�lO�)&Ѩ����2�v	��ij-	���Ukۖ_�ѽƵ��P~��X��X�.����z�(Ǝ�dR�JY��֠�I�GӲ}
f�)Ql@����R�&|kΏ�LC�뢖A�![G��`g��>��m����ϭ��H�>���}	X�^8�4�ܶ�ߩ3��ty��$O@��Z�:�g�������~Ӄc���X��f	�x�[��v����*�4���0X+���'��X<yeI�ۮ�Y�M>��Uǳv-�S��uSO�B�Ǿ?10b���75�2�����u����Vw�W��;mĜ9߄�L����/e�%��S<r�?b�-������Y���L�3�ks��"���5��4K��I����u��/�W屮�R�1垽�e<@^��q�+��ŋ rY*�2��k%������~��m^ � T���`*� >�?)��C˼@v��	p^c��[��z��ȤQy�J��׆�Lw�R-��<��A0� �U�|����O���<��G@�u���0�/(��k�^DՐ]4�i��=F;��H����� ��m�I��7���a��F#��E>�k>U�8�����wU��1�C5':}���4_���Lemp4�MKz�Ê04��7����b���=��/
jU�~QFz�8�O�F$�W�@Ѽ9�I�A�3�Lī�;�%M��5?$��P��jT-��#�c���7�ͺ3�m��I�ʊ�Ş�fϹ!>�������7�"��J��
����
8l�^d<�N�>|O�N���sT���%�W-�����,X֜�bD�n���<�@{~��zV����딳��񀑿{Ep�-`����A�s�9�ϯ�����+�?����х���՚-Ơ͎�B��/D�a��� غ,aW��Vjx�v��2,����Ctʉu���R8�`h<���5�fCi.�Ji�v�+u��e���$%��Er�D��S�kf�����Sʅ�#i�����;�#��ެu�LClS����Mu\'�vٸ�� ިyBY�R'���~SO6R�8Ǭarα���FB30�j��>kc�r�C�a{ZP�J6�v�l��D�+�����n_8D���.��U�08	б�-��Q�4e�V������@�*�(���B�A2:����x��73�Q.�³3���O�%��2Js����֌Yj6Ev�M�Hm�az�8��jMn�&��|\��n��	���Y�{�l��6G�T,?B��-03�N>j�`��=��g�]+,�+#��-�����$;��W+iH���k��_��׿g�ñ��b?�Y$oRM_�MFj��(���Q,fz��͛�OX!��D�|��T�"�/k�j�t�-ݍcES�͙Y�2��������Iڒ�T����)��a��*v�^�"&1��A�7�T�Y����h�#x�>7t3�x�b���ݾ�1��{�]�nO�����U�_)�����O���J7榄�v�A5z��O�WTi@U���j9�|��OBf���yXe��p�;Yn#�U���W�+�`p���nd����䋾:��}����'�OT�B�u���uNlY�9	���V*@����u8]W�42�!R����jt�q�x���O��$s�rf�Mu΁��XvL�q�K��.�V���~x����� �&e���h���8��I!�3�˴M���?Y�����gQ���f�@�/�0��f��e�cRE�t�X h"FJ�J�=�b&�Q�tS������W���~MVtc�V�G�T/�DIq����U�h���L�0����NZQ��.޼��:®*=��f'��"�Ny�id�Ľ�4^�����kEE8n�BpY����@������$�q�Ъ@T����\�&��r�s��{�B�fk�c�5 �i�J����ng��~��� �5�5pk����7ʢKFN	y�U��D���R�8)b�1�'*S���#]�����������F��~�B����9L��9lƑ�.�h)�	�F������w��N;��<������gQ|�/�3��p��� ;��-�o�)uN�{ZCm�paq�p'��]�@*����S`���V����@����l2�p�}��߱�k#{0)��&C1|-b��{��:�J�g΋c�{�x-�.���-���OwV$フ���B�J��U{50�塅����A%��t�H�"�/!�6�}6�+[L975v��X���/00�I�p\׼�}\T�Jqr�YtfG�5\������˼�t�S��ge�>���V�.���f� �m-��Io>��ˎM���- <oMˊn%��.I�`�|(aYx��RKw�.�����Ȁ6����gX�X0��L�ے�	�ʂг����w
�Q�]�Q4ևj�4�%�Y�ЦgH}nm���`��*����Ŝs�Ka��/����PJ��-�Ȕ-j�j(����}.'�a�ɖ	`��H���m觋E�Ϛ���~O�p�A�"ؗ��!��QE6;�E����@��5|BwgI�?�q���(�\5�#h-��p�8F�)�l��J~-E,8����w��ɼ�5L�4Z5�?W�@����+$܍�|�+��d����A��Ù/!���"����[wa�߂���T���1Ylµl�/g�Ǝ`K��i�١��Ϳ�+-�	O��Q�1`�6�9ubT��I)qS=?�����b�^-�7BzL��<���`����E��3�@��|�g@�r��
�����Y>nI��O�U���_'h{q�؟H9���^ �9��s�}j%����(��A�.���#ǲ�?�J�Ť�#0����5k���?�"'����)�5��fZ��K��j��A�X���Q�(Cp�6�qȞ��'��1 ��x�p�zx����f/=�B,@Xf��Z�I���M�;F_�O���x�cg,҄

֑z����"�]l�H��U��p},}�|C��h3��dXK��1tK�j�ԁb��(D7�Xa�삯�p@��\?vPW�J�L�܀��F����f���6�(�/��e���l�SKF�d�����������$	k�uB���X�u���'�A������x���nV�6�֗Md`%+�"�΍���E��-�G���dM�8��窘HW�Gu�3<��m���i:UMԨ>C�y�Q'���Q������S��F��#K~�̰ �d���ä@/OLjȫ�-줟bߙN�g��=�۹�a��i��(^�ђ:Ms�&a��H�|J-Jս�����,d��`$���������$��7������d�$,�nhi�m�L��r��T�8T\Q�^y�,���,�0�tmݹwLJ�f�pݛ����V�R�����m�I�f�Ƞ�S�~���%�e^F*��o�x\w��I�Da�����j����������<���2��K���A6pJ��v���Z��{�B`����f�tَ�`Bp��g��zƁ��]��|���0�0k_�W���Z�dϾܻ'�\-�Q�Ϛ4����X���O�©T��q,ZD"�ECV5����8�gL0�3t���D����ö���ÿ#:q?
�z���A0���E��$���9��G;쪳�H���{"X1�	�¾��HZ*��>�D!(R�F�ñR�.W�w$5�b�[G��<k�Y���h�d��S~8����C
��ŀՈ����B��*�2����~��aq�� ��5��.s�,��>JA�"����W��s�<�Q�i�D<%�Kg%.J�U�= �HÂ['܃�A�ߎ���I���b}M[�Y�ܺ��J-���J�+���1�
/��Z�� �%�|�kM~?���<K,�7�ܐ�Up�jo��ӳ}�{6tv`���s۫ZN��XG��![䔼�h�Ct蟯��c	w�Ml�2��z����̗�[��[]�4�V�?P�K�A"�̞_>΅`�w����˨~��7T�<0��j@A�����-e�R��#VMe�;ǯeO&e��lN�T����Y+;�Ӷ���%!�);���!*×<�Or�Q ������Oz �'��҉�\�g����I@w�L���t�u���$/r���Ew��>r�ٚ��]0���!��ٺ-h2z� ꀍ^�ş1m��n	 [�"z�QR
lF�cv��:cm��ZG�˅*�X(��ǘB9U�N�8<��.Jk��& �5b>K(2+4�nf���X=g�Y����Vg_'�>��'�ʦYM8� �׭�^�� W��_I��?;�	wތ�<��\ω6T�C5%#��E��:�mx���?Vv��A�m���p��[OS'O�Q��������k�|�ZF�Z�{`A�r��9�ʴr0�kh���W͈k�ւvB�j<NF�W�$,j����څ��u������5ٚ$\(Nt3ܡ"�Ɔp��1��ү��p��^k���C�u�&��s��l:T_��{y�4��<*������5ZOY�p0A��F��ϝ���(�n8,���v?$�iu��JR���_�v8�~1O���)0_X�GrF*���I0	��6,�%�o��=i�=q��R4���fnYm��q���a~��~6Bcn�l��J�^ш�9��	�PpP�t�uL.��w���"C���B�x�K�E��O|��,�ܥdTJ�u��)W��=�|���ĘL����[_��]�e _|mR�W?Y`�(�E��3��$�Ԛڿ�jj>�)�s�5���D1���:��{n���1�v��d���MX���b�`��:�V�n�F�m�J��c����9�ع���8���v�A[`j����J��D�:�򁓘���o\��Iu��Tŵ��yc9Ѭ�Da�;hc�.�o��~��|��e�X'ʄ��Si_�	����W��0i4��Ƣð ��0����3�c���z���lO����5�,�'3�Y=���t��L"� ��$8�N����l�s/x��DZ�[��Z1�E��ۮ/���R��V{򅲜�F�p��+3�����G���΂	�"V����pdZ���(c���`UR�L���|Y��>a�R? �1�����Wн��U�%�Q���n���^~����b��S�?��}��T�=�O�C�]�q;��ݘӜ��Im����E�q!� ���D+��f�j���U�Nc�!�+��I�7f�GQ�H~��'����C?oD����nc�H��?��j���U��_a���np�á�� '�̵��C�����J:`c��+R���xd�t����Dq�7eU�RsĶ_W-~�L ��%s)X7g:0
����`�U�t7�+�w���*�0��{sn4%$i,���Ca8a�?%�SF�Ц��.&���JQ%:V���6�(���$�߁��֙��m�D� \�Ԃ�2Sj��Ey�k�Zh^B���<zKS;uk���0'DYU��&++�gC���g^�Ib�M�<�4���1s¾Zh��@t�#�:w�B�B��d.\����jhxKRe(�D�L.���Do�=��m�K��Z��@���P^��;����N�6>'�ȢUv�۽Q��^>��{��owU�Z]�����8�8�����O5ҩ��C��~�ߢp� r�8{�Gg�`b� u;Y��q����(os�}(!�x�=ô���z�e��]�G ����3'���+ө�촎���60��Tr�A�<�J����wvF��5��ҧBҝ�Ը��ja�m'ˤ>#���"��[��)��m�}Q6ײ�
K0f$���\BKg*�jm�9�,����AiI��I���{��щV������+��l�"�
��q���6��e�K㆏_%XP��a��/���1�b<����8A�t(,h�hټ}�A�'��QT���P����`���4jų���׏<Q����~2ʆ!�q2o������J%��]���~���N��d�"�����9�SZfMp��v;
��+qf�Jj"��c��H�V�2}G>� k�8��z܆M}��m�^�t0}N�3��N�
\R��r2�ݠ�k�G�������6i�h��8c�$&� O�(�)i��%���&���}�Vf�XP���B��>8��'��S��4���@;v�(鸩�*�-U)��8�/�!a7�7=�nJ��*������`*�Zz�e��nݭ�0��Ss7)�w�.6~z�HT�~*��L/}����eN��\O�^'a����Y��)K��2�\�Q'��DGA(5g�,�[ՖD[�(���+�ɻ��:�Y$�x?��u��{�sUֱg`N8�CG]������N@cx�����<C0I�O� �/y��d����b��a�ꃖ�"�oyv�[fM�&�<5�π�B�^EB�9����5s�֣�!�T����é'"���g���Ͼ��E�C����(���1x�/�F�0�N ��]I|��BT��Ω�c�%�m����]��Sm`��k���/���,�i��yDqG��m̙���F��GC0��U�����&��X1DK���<��zC�>�/wؚ�>���iZ�*Z���`nnz��\`�@M
�0��^��4���A]H�+B��3}d�p�Z����@϶�u�$��%��?�h�|�#�El��=qnq�F_0I:G�:旀�G 3N~�f�#��"� ���E0�8:_��މ,u#դ{���h��(�*5e/���%9�~�f�H�
�׸����]��˲}��O��FS�Q���X�L�58�l$��7`RX0_V��٦�I����ns��/�6�O�~��*55�_&�p.�n�����H0�GYl��_�8	"���
[�w�o���I���%�|ѶpQ��ַ�q�GF=)~$���B(^� ���4��zJ��:��G�A����b��
���	?v~{�tS�k��mK�!�P@W�+ϭg��%?�GY^��#���caz��B�'�Ě����o�X4,��	S�A�h1�+�I)�Έv��L�����1Ҹ��G��(VO���8�A��/���=�@�F�Px��ܧM�Y5����,����<�q����h՗�)�<��S�f���p��|�yyGH/����qty&H�z+��\��I��<��l���d��N���"��}�CB�	�^��y�E_w̕��>��i���!	EU{�/"��Z*����k&��1ZR^�`�bV�?u�-�]�9IÖ�ξ�q����\U��ٯn}x���+'E��ỷ�Jr<Q���T[�7O��m`��d�
�9Z(���j5&�bَ�1�?�ϕ���d���Z9CQ6gh<�t|n`�W�FHUΫz���Zd�����!��鵼���Qrg���^�}<A#;�sI��������Ĝ�����q��;BՓ�V.��2������;���+H7GJ������ O=���ibw}���1*&�Qƺ�_��v�H�sn�<��l��@C�#�@$��X
���$�X�����`@����#���$	���v��کS��M#�i�ZKyĺu�L�߳��\b �GT�Y�ن>,�;S�d=s� 8JJ��g����r�� i�'����"NA(�M4f���j4u�g۹���4��h�{&�@�b�n���m�T��R�Y�lK�@��"⯦5q?MW�][�c5隽o
���d�~�	�ں��+�KR \�|�/����f�zy&ݫ�\��Xf���ߦ3�'��W�[�e˝�E
�^@*4�~/4֧
���2�́8��ș�¯2G,��������FU��������RհdճNA �O���<Ӎ����7i�����C�t$���LS���?��d��=h�����ȡҡdK��f1��|�L�8��d��,������|[�r�ʜ�� �kTڸr>Q]fNY-�a��}cbS����q.u������q�,��������~A@%
�tא�o��:�'d4W	 �M�|��}Bww�����@��]Q���n�gō�޿0��G������( �D�]us<�D�S�[\�[BkLQ�L����"h��	�P����̚V\�'�󓿇4l�`�Xh�4h���ۄ쀄�q�\5���|�k:�m	��;O��@�g)��R��+x����Ε�����x����1�=��G��{w�T�y�:�N�����C�8t}�e�T&s�I�wԣ��M�n�t�ag+��z벇2���4�c-���T���F�%�n`�4	�*��)��/eӾ�"��Tg9T�oS
z)L���E�/�M�R�����ё� ^�������$2tB�Yo��(�d�eE 9%��m>���dwR�|W�7��� ��l�o���b@H��㓈�b>9c
�00E���$Z��%���������V~ɬ�w��&��W��Ԉ�0����	�+q�NUw1��jp�ʎR�d�v��JTs9j�c����̆V���@Ao��<��	�.]P��D�q����H��%�M`X������`����4���WIZZ�+���م}|�9�&�0�Vr*
(�
�H�>������rI3!���{p�I9)B���L�(� ��;�[��)f�Dh�=��/�xr�S�n[Q� J�|�=9�	���<O���2����9�E:����0ϋ5K���#�/~k�9�ud/��	W}N������dx2�"����p<�|��W�ę��{��C�E����A�-��]:���R*b�˗��t_����x��V���K�G���ӭ�SsJ:���	bf,�3▷�����5{���VW��mm������b�u���a�<��>���K����gI��'>S��ci\�[�4�nY䇱1۪�((a?.�Գ��b��\���!��a��C���ʰ�>& ��7�p���{1�w���~S���
�&BW���k?
ɚ��2;���^��tֿh�k�0%@)M�|����z�vu�bC&�\<��@�N���1U^U)#��ф�,[�9�jJJ�?)���J�xM:�7N�=~>�n�d.�7zI�d��i{�����������)��pe�k��W%BKv������b.�!<�MA-S�J���ñx�e�<ᾰ�畺36o,ox��v��͸ׅ��8
g ��dJ�t��i�b4Ü�c��x4Cߝ�+WKy��9.�$�6����r�X���q�j�z���B�?X*�T-a.R^��� �dUu�֭#�-F'�2�~�N�(�)�e�qzt}SQ���YS�꧋t8�
��<#�7�	�l��0FSԠ�4���h�\h���(�y	�ȭ�"w�XիҚ�ހ���r���F��Zh'��u�y�u܅B��l�qg��H��`���f��1?�+)`�F��9q�+���u:3U|��Ȅ5��FV�b /A`��4W�ĸ��n��x�X��q��>�+�Qwۈ���Z�0?0�5b.	����R�9��vm�$�&>���_�!��/|�фp��u6PiXǠY��������Wj�& ,so�����5o����D�o�ʄ]ȫg�7���="\���S㓙�!,���Y,9��K�WQF��+��9d���',2��	�Ɠ����)��f��bI�h�B��^L#MW]�A���W���UK�мн-�fD:S�?F�]�X�Yȉc$,������M%bi��s՗��b�F��9"��������F�~��o�t�=���8���D|Hx�Ӣkv����87��C�q����bDL�"����������E��{?h-l���/,��h}lY��WXo�_��0E�U�"�)6"U$�6I�ȶ��gߊ����v����)h�B�d�l�-��������K�+栦�.���b�=Q����4��ۜ���(Н�	��?W=IA��D�M�SA�GF��N�?nB�\�x�
��MmP��ɃүǿV]7�j�t�)L�^#�qP4���Fn���l�7�+����7{��M,P$}��O�y1\e8z��R�s�x�Ňj�`�I4��ç���v&�#�h�I��ޔ�03�CQeG]z�c�r6�q���>���pq���hDG�8���J&�4:�����{�!C�?a:Fl����QX�=cX���^�XG��m�:�d��Aۀ�Z���VP!�6�3�K��P���sݦn�����F-�L���aG�Za���E`{�.�c��%mX*�w������p�F���3��n1ӽ/}@�'�c���x���L��J!�c�;v�K4aqJ��"hx��j���\7g�4��K����|�scQ[#���ĺY��>6����"d�d�y�8�~WѡP�/}���o�q'�p �/XsRf�NA+|
��
)�(z�wB���ȏ�b>�ۮ��2�:'���f�Ń{��W�ʣ8�mP�N����u���>&��+Nn�{c��&���������B��9k���_����rD��������;�wG��u�F����s�~�� YZ͕�_Y_���#� "����:D�����I��䈍�&\<��a�'��񼹌���T<]�oE-n����ﻉ~[w��e��=?���ȝ�y�嵽����6���EF\f���Ϟ�B!{��]�+֦����sb�k�M��Ov@>*9D���z2f��{�)��S$�mfߘ@�P9�v���i4� ���,^,���jKD�O%�%ۻ����a��0�qc�2xb������`�Pl�`�+m?�XL`W��2P�����Ƒ�DN��Po�_Xu=v���-,�m?�[u��[3�)_��2�{�	m�IL�ÉH'mZIi�G>��������c-&��,mE��Ǔ�u��G�{�B4��/{�6p�{�{j���H}��XfD}>����2d�M_��uR�a���:<~��i�	@���5�B��+<"[���5��]#� �:�b� Ieg+�ɀ
�e'��;;K�aJ���H�Y�h���ǀ�\Ƀ�I��;�R4��'46D/c�v@ʵ�?��r� v7���0@���_�͡�*��X���o��9��:�T�37��r�8��< �Hf�`bO�A�bp�\>����H�炻J��֪xj �^�:�.C&�A��^���&��k[�K� ��IOR�w?��k�X�g���m�ڠ:w�-��h�����8^��?N!Z=T���n!`�>@�}C�<�q��j�v)�)�L����o|hҡDS�~����zU��ۡ�Q]�(j��h��V�}5��ı�O����zs�d�;�_�`}k���VQO����usz�4�-�s���.�Z���2"/O��Q�M��Ő{2�㸠��]bmX���-ozM�4��Ѫ�|�|�E���Dr)��!�m4k�6����YC?SQ��#���� \2��| �6�)])��!A����z<�$�ĕ��cdD̗�����S��z�
����t�X��҉U�ٚ&��w��`� ��t�X-c�<���'���mk�'wf�t�yU-�f$�^����Kf�cM�p���5�Ò��~�(�ր
8���0��y%~R�����eVGLh�&�? *$�. �De�4l�J��\ɔ����j*�99�|�Q�\ \�C6ܳ;<+a2x�E������ʏ^sF�2��If�.Z�z��@6�Gl�+�N:������Py�ND&�`g��FAm�n5���&�`����;���8Ptk��v�m�ٗ���ϫV�xDp,Y�jl�6��U���<�<�V(���pM�����z-C�PO�`c�m0Ţ N�&���������.� 9����6
."o��\��5"���z�A�i�K���H �o�B��7$}��U����&�+΍z�<:O��΋d��6���a<�|�:B#j[��K&�#"d�=�]��VpnEݶ:���owZ�#z'��R��S�8"0�i�����R�s��.E1�F�bM�=ŵ��?�i���q�1E��pp
IDv��9D����7.���V6.=Ȍm_��s�&:�o�c��7v!�D�����1��J�������m͡QX�E���h���pL[G���ȷ�O����rKht�4���l#e��5f� f�)ԡ�t��O�ld�o�*�'i몧'f�N,7YA�g�U|yQ_�&w8<8����^>�ꃥ��n��!�� ߤ�.�cz��Bԕ��K��dߞ����&ڎ�I8[�  :v@I?e�>��z��],�����=�9����J\�Ƅ�0�	��O*(~��s��n��Q-6�/�1Eq��	����csB;f�f ����]։�g�I�$x����ݼj@amg48U%���K��s�$�q�QE��8y�r�c�o�$��^M*�ܯz|S�O��9�%�;��:c_S.�Եc�<j&08�h�7�S�n�;�pf�0F^�� M�A�r����Ըtb.]W�������,�:9����#ǀ.��o���^��X�պ��X�ͯ���v��p��W��./u,�HBɲ�\�g?���F_�Gw�l�V��H �����U���OM�+��e�~FtK���܌��gu�Y�:,�����v��M���X� �ՓE@W��� -�r�h��n?�z.a�]��t]C��_ëg���꒰�3�Y@���HZ�^%��QP�4_N�TU�_��\�1�Pʒ�+��!�T��4A�����1]y�ʬǯ<��t8��GЋ� ��7Ke�դ�
(�Aa|('[w{�{�I8�OS7���y�E�7
a�]-�;�
�<�T�T+r�U�X�z!_�_����������]��L�����z�d�� YHi�7-H���)�C�`B^T�[��J��h��5�������ôC�3M^[�ǣPP��h�,!,�O���#����cAB��}!s\C8r�K%�%���KRz
��	��]YN��X����� ���ɜ�s�~nP���וnf�m���Z@^�i�W��¹�jL�^ʶ�UwzV�5�nD$�*4��u��X>/>B�j(�5�J��(]O%���[����;���0��,g�؅����d $ �!k���bE+a�l��� t^ꌣ���3�y����a����:���0��(�DsgT�$"Q��Ӹ���a�;L��j�����}��k�3��h@����[��n{�������}��D�\���u�[��#��a\�Q��^#�ZE<z+�\��<�e)q���ny_$�F����W�#�<�S��@�5r$oS�b�! iuc�@h�-ǭ(��z,ը�3�������W��ڄ�������VL���Hz�ٔC���2|Ģ��,^K��E���S��=�O��q`Za�T���J)_[�!"�@�)��)'�faa_u�<��L�d��c���z����Db����4)�3s����c���o�4O����e�=�?呀�f��|�t_�/-��b{"�sh�'�3M��:�Ww~z��`��ZK��p������Ђ�B����7Ҝߎ���f�k5����PTV}�AwbV�ds��(�2?�=:;e��;Ut�1ro���� ��P��w�<�(ȥ*$����(�ɷ�2������z�t�%9�r4�7ׂ&��)�r��Iڷ�s"��/�I��!���3X�TN
�fI�ؕ�����Y������V�E"���p���S�T�����2)�nS���#{A�JXT��N�P�9�9>��hQ7��|��8�.�� ��5��_���4\.Xi�&�{f++����)�|�2A����ƅLr��I��P��,�V�W�Hr�A$C{�h�}i�5|v��	�B�b�"��m�V�黺`T�-�D�.�k+��9���)���A��	��@u@���Y4�8��Q,	��_�v$�X�������"�Sn�]v*<���=�� -μ1in.?�%�Y���~:ȗ���k������=W#��l&��C���#_f��Ҕ�N�bG���/J�P����:"���?���R�P�:�2�	�<[M0t`\��=	ԴsVCԠ���1��iY����N�����p����r�E-
.���?<�x;�^�H��۱d��&�=�D;K�7Ò�{{-H~�61o򪟌JT��j�ͨ�t��]Dݱ����:2�GA��sؗ(����2�-��ߤ�����u�N
7���y�9Y�]����Sad���:~U��t�BU?�Un��\)���6+��|����"��YNح��^}>���rJ��O�{�4��oG}�JW鬪 ��aC����Fq��י��`[���'2C�W���)>Q)�Kr�o�s���%���E"5RI5�r�傟PۦvAu�9��Rϡ��䙖�fVaEV��l�ǧ�fnq���E*��a9Q)�]PFb�}�o����	�
���W'u	h�YJ3ƈ-a��P�9;Ir,���Y�(I���p:*��붷�	�b(F�����~���RF�\���+�ß�4���#ti�2����^�د��靄��Wa�J�]�vp!�S8��)V$m��F���� $��vh��0"e�{t@ڇ��D���I���"biP@�N#�&P]��KAz��:�R:"���QW3$����_>�Dy�=����6��_�V�>J�`�ڀ�tp����K���Jh��_1L��m!�o.�B��J����b����8�v,g詏{U�x��Hb@��_X]��G��e�����|��'nt
61�'��	������|#W�v8و'S����1"]8"�Y��88<�Z��_��)є�3��t����$���\
Na�/���x֤ڥ� ��A$�S
��F�Dl�����V.!j��/q����ґ�i)�mo2y���B�1e��6���򧴇���m�Co���QGC��%���Ԭ��d��*M��o��F�#��;�	�<��*����v[	�y-��� 7ޑoS.S>Ѭ�7���wY�Gu��.��e����fH�/	S	1zչ@�Xm@�+����3՝����2l�ݜ��1�Pc&�U�$}�\)wp�lW���U�
����u�Z�2�����>΁�jS�'ob��G�z��"���6/�gS(��"�7t�٢��S߾�p�EOyN �E�ov���,��8��a�a�F�Rû�v\D@���-�������W��t�L'~.@v�p��j�&z�%�?�eZ�^��U�m?�;Tv��E�+���h8l��evu��DU�3tֶ�^sTjk�or��p �[	�j��M�L�jWfv�h\��w'9�~�e]��j�7�Jk�1;�R��s\�0l/��(��̬�w��.�~=3�d>�v���"ۀ���_�e>�zډs	�h�j�+#�3�33���'��6'��e�)n�L?�D'�t��v�����#E�8�2�4/����VC�㍹{� �^�Y��QbzD1��L&?���_����[�)Cz3�ߠ��&�L��Vҧ�/�����O�1�T�������S��u?���"y�V��㨕��%���5�H-��BR�	�b��\�ĝ�U�����=4��{�e��g;V?~܉�N<]�\�GZ��3�a��$����z' d��F)��~���v�"prTy�DXk�v�pW�k(O��+\�Nzh�@�N����ID��6"l�s�Y��;&`�D>?�x�үK��;Q�_v��2w�o���+]�sa��x�ePQ��V��Mܚ��k���m��N��l��j?L-�O4����T�k�C����f))�bm��Qt����6.HK�1@�������f�?=_bU���u:�YL{���4�� "� "A�hRpKOq�VR ���a���3��y��׎o	ccy�����V���Vս���R��$3*D�j�`x{��Mt�2iJx紨�46ʄ(�*��c�i.��1>������Ά�n_�Q�7��zF��#_UŜ��HL��~7����D����N��9��f[�ɏf�w��)��Z3W��ܿ镚@��q�N�>3�)ӺtVw��h����ub*@�p*LO�[cD$�@kh+������9N�7�~�È���byw�\<�I��~[�̙�Q��WT���g���.�DðK�'��*���%$��yO)���m*�W;�M嬬��>��̲�$�������,2���1��`&T)�h��EgbY����I���t �����e�M��[��V�Uf�U�6��f-5m�$x��=��.،����}��	���������W����B8J�^_i�Ui��R��˻Mq�E�}�D�\꿸�i���8�p�Fۺo���P��p-��$�Ƀk+wBB������)
������$c\������rooEn�C��f�I|��.j��Ѿ�q�%�y�d�Ƒ�<�F�C���'�<I���
���tD���n}7�*�
��gΌEb�_�BXzMܚFB�dh5`Ȼ�B`U-=�'���d�~�O�eF���K�VK
�R����>Mi�� H3*0�~E��:�|��Y9~����"���l�����g��ɴ9֪�h�f� ��&`V%ux\o��Yp�adQٸ��>�x�eG�Z?W0���wŘm4�#�9���}��K�x���1D�3��� IS0�b��|W��9�B�$`�/j��n.���{(����E�.J�"��N-8Q������¦0	�'4�����:���U�bC˩��+�^���@�x�f�i�X��Д�^�zj��8�'�d\-��jf዁��:�2BS��|�P�e�H��A�MJ���@j�S1^CH^i"K������#�[\~Zlk|�ړ�J:$��,Z�a "��g��N_����ѝ�B7 �Qsf]��?�J3��z����ъ�'&�Q8P@l.�-�T��2m6!�+qQړ���Kj{�fi�W���Z���4���2����-�>��*���@���DO���� ��eak3,�3��u �P�u|r���g쫸�I�\� �Ϻ�l�V��ŕ, ��
	�j�����л�?��b����W�������+��A�l=��svc*^	f#��Q6 Lz�؀1	L��|��v�@��i@?��\t]/9d��$'���m�F�{� ׻�A�����gz"��E���	�#��+>�$@5�I�˨~��;=G�v]����}��d��-`кh�t��sH��`ҕ�oL���f?��AF�nK��N���=�&�)�y<^����-��2�q�x;�����<4�k�=�k�K<����_,ɠ[���ȯ�+�aP,`���P��j�K�)yf�0�~P�D��������}�����]�J� ��(����/|���P��~ b<�j�b��q�&��'; �{���^��$޻�)�P.�]y`�s}����}�X�L���F"	`x�o�m���\һP�@�r�1�vwLg��6$X	 ]2@;G�Ɓ�Ι	�ߋ4@�U+�``og(�y'qȾe�t��{��X'5qQ��(���ĽK�i&Z%3����%��~�I��H��T"�WD��5�_�$JA�+nsQ��-K�˝c�XP�����x�h�ZȲ�x\����� ����G�.���W_�"����q�gȘM��*�,? �532L���[ED�/-��C�Ðl����� �Y�Vu�3�;�d�FkB74��s����~͠��ٹ�}��{xkJZ��xRo�I�U[�O�h���^Z� ���a&.1�
�a�m����S�����X%O�%$z�eQ��$�墕��̑��d�n&B�e[:��V��i�2DA�V��V�i	/��y���'5�G�,��f=pg�w�|�n�����T�{�x�;����5�7`�G	�؆�+�*D}zϡ��2�j�5{�aK�{�%f0���a袍$Ljm��z� ��H'��P#(7"叩�/z�yj��b���V38bk�U�:����~��::}x����A��9ֻ���]8�NKA�9��_��=����]V^
��=1�gGw���\���P,T�ȓ�o�}�Ko�GDJsS�Ũ��®���*CI�����B~��{}��ޘ+�؆�U9� PuH
���θ{1�S��ؿm�����o.�+_�V�n֘�"�%EV#U߃v;+�1�F*�_�<'*�zWv��TU���zz�1/�z��-WhfT�]*����=87?.�(y�c�6�.E:39�H�G�)�s K�� �;�R�>�;��R�)m�j̫�W���wh�����%J$ټ���	+���B|:��7T��n��l�%�23�|��G����Gka5b�*�v���'̢��	GF��;j�À�P�s������z<�c+�K�[�����!��MI�#V�29^E����=�'�9���Lƿ�8��a���P�/���˸�RTi�D�
K��p�Db�=�������s�ŧ�2"~�&N�9�Zu�x�|�Ƕ�X��S��cFGaJ���|�k��Od��(�A�(�69�wb�ǼX���4��^1.���cvp����Ko�.���D��	�V��Yui�'������UK-�/�kN�D��jm���Z||���وW�*0����׌���#�~���'9)�����4>����<1U~�,j�b���hi�����B�
���¤ѭ.����)׸�RH-���6�,,�ʻ�6��'�S������[���?M�0��S���%�ΰ��Pr�{@G�j�[Ik��*���jzw:�*V}��]?��j3H~�o�́��n"\�a�E~��t[��] jt"��rf������g>#K��ʹ����w/��A_6��Dċ�+n�?���,�+v��Q�/l�1;�v�s���>��V#��yQF]!N� �8F������ěr|�'��g��hȯ|s�u�q&�~u������t���~ E�E�Z��K�k�?4�6}������;宱^�;�m�dę���3��$��Y����ȇP�HW���z�;B����C���V� )�S�J��Y�o|��/<���G��t�gj�K�p���0I���ݵ�*�<��ic,�n��B�BcR玀+pj̦�d?� .��e���#��>R?HE�Vw=2EԨ������g�����n�^�+M&��' �s�B�Y�qg.���MH>�Rӽ�+���Μ���5�;�`�R���R��5GD��Y~p��� ҫiG���[t����	`�y�3]9VXmbɐ.u�^���.�R��Ѱ��Չ��l�9��|���d�֢ hv�SҠfI l��3���C��/UJ�����5��y�Ҍ'�\�/�tS]��}l�Rx���<w�ػ�_�E�L����u�.���j921���Q��5��U���E!��h�X�}� 8��mD�����	�K�M
"B�u<D�t�IJ}���ju�x˞&������e����R�(���=
�>5��s��\���ތ3���/�4�� �?t��pcF��7I���T}��J���8�aY��w�Nmm�-'S�na�����}�6�d��]�G�d	W��^\��<:�"#���B���'V#���qe3g�0R�y�C�Td�߶��}��w̥[�@��Fv.d��;;�EX��R��bWVo5��h��A���L$zYP���u��S-��Y�[d`�S���+Hca���Q��׺Z�Qi�<p���Z�(���C��r��_Z+:f��E�@H�X��ގp�)���P^]ߦ��ۺ!�6-�Ci�v��">[@�����Z�f/|^!c#�%ż�xB�H����sAT�Π�q���z��G{B�\����3�	
���	l�$ţ�ؾ��U�Lw[�W�.G{��o��Ԭ�`�֓u�!���P�dԘ�r��Xl�[��Z��e�F\ܜ70�~>^�mY�h�D���R�Q�����ʽ�BSD��ȧ��Ŷ���&WA;�����(l���Uu>��QkZ�&�>��Å��'�&C�����1^&z1�f<7��f�����#׫c���BB�O^K��!�%l�1���l�ȝ����w5� X���@m|-Ƞ'ǃL�9���[���簢U�R��:?���A9��R��9�ߺS��6��^����U�V�I��`�d�U=�}�ߑ���Pc_S�%��[���K�\nn��y
Q������L�������w�~Y��6�!�e�ڈ-Bl��{TD<���Ȍ�H1C����sV������n(��9��vծ���Ƿ,v�n'k��D�2^~�O�T�h�:�c��5���>��*��Eo�Y�P>^&�������^�Yb�Dra�L����E�����Q��7t��Uz��b��D"\ܜidd��1[Z��A�7���.6Q"P�? "���D��HHX=���C,:��Z��I	Q�"R	P%������{��'JyS|h$��v��<VާZ��
���(@��1>�7F�X�ƿ�$�1[����/s:~���@B�%)�NW��97�Q>{T���#yȓ,��1=��W�2��њ_0n�}��
j�e�;X�E�g�
�C�2��dG��yT�}�ɬ��+��S_}�W�P�z�N��
RW@���ߛ��bAÍRKY��0ז6R�R�f�SѦb	e�r��~��I>W(�"S��`x�m�S3L��yD����;�e�a9�[=8lz�r�)�[
20���E�tGI͹��=��/~nX�?m�����1�:�S�t��g�jP��:('f.Mõw\��U=8��J�'P������-c�I��[�g��>=oŵ��,{&	����~c��t���K��;�ok��襵��ʮ��/�z=��:Y�fT��_���4l-]��ACCּ:�K>9�"Ƃ��P!��π�g�gI<ĵ�������j8(�Qԡ�TyĩT��8�<��}����r=�a��V�#�E����s4�#=��KMbU�/����5�?*���(۸>D��Q�2�o�P��Y�K�0t��+�}NQѷ�[�Y�=�{W��zSX����!��C��
;/�l��nR�);�k���'�ɣ.��&�I��Db�>�� �T���_y'�0_�3gq1l�����H,�3���H�z��07�D����#��%��Ȩ�l�jRt������t�h>�p��K����G��u{à�1����Qz�% �/pNQ(�Nf��{՞��D�w+y����9��a�����P~��JX�D^��7���KŘ)f|��:w�D�b���R�呱�]���I�HƗb���������F��?șwo�(�I�=Fd�t�v��B2���u7ε]��y�;�����ŵ�����h<?I���I��8��qʔ��g&���｝T��?7��P�1�e�B�:砰��{��H
<��ˈ�p�b�^�r{M��|[:�QDADj�`��섞^� �l"�p��:ԦEqD%ۉ�� w&��*���>�4����\��=i�گkk\-�v��>ʝ��+�<.I����*?���(ؾ�����pg	�$�w�A;*u��
�z��mHܒT�ęı����e�iلl��ȶ�>?��j�"lQ%��o���%r�t;8ʛ��xT�(W��Gr�f�� �Ȯ���j$=�'3V;c�z�I��<f���
���U�C���ۂ�+d�Pp�b��]O^5���
�=�b�&CQ[��b���t$A�&t|��Su
��SgoΑ �v�(Ģ2OLT�#k�s��#}��"l����%d����69�W��t�*&�����h�>���o$L"_�ﯖ;������]����jn����"H�[�ҋ�թ��Csˑ�x����P�� �9-[�u.�s?W_u���r�B22c�#���_������� �=�o�v�!��h���Ld�a��wɱ�Zv����QI{�\���E�/�c�z��mS?a�Ѱ2xt`�\�g-:��c"��"`�Z�^���~�]Ӊ�|x��N����E-L���;���l��w7-�L	�=�Ar��pߗg���(t��,��*�@��zpizʪGd?�'3֞�X�q��ƹ�:-Nc�%�S�|C�Ӫy�eH���5�A��E
S$,N��B8������8��:>��O�X }�����2��*X`~a��`��࢜�U�
yk���vi�4V
]M�,����_1&J�0);w��y�8qY����,�Z��Cq�"�# �`�\���o����R���U���Gԁn�&�򫮍��4&����@��F�oA�E,h��E�z=�Y��7� C�}�:���~4l:���U\`�n��ݱ��z�:c/���)�J�������-�D[�Q)�F�e�c�d���Jed��^>���
����g"\x bߣJB�	����^��	?�6<���������J��д��"f���h�`��%��נ~Y�ڠ!�z�Mw���0;g3�  D>v{F��n�tu�e��ı��n赛w�s<#E�� � r�́^P[�|qJQ,^#����0@)���1��Vg0�(��n`��[���[T�C�(ZO�+<!��%	#`x��b��y��0��|Y}O�V�}+ܟFn���2z8��i����@�CV�|������� b]���?W��ߨzĳX����J��vP���W���,�u���wA<�%�K�����a�Y	��E�ynXe;��Vd���$L�>ԗ\2��RC���8�;���¢^�]����W�vO=�0��[��v�й5����@�h��~������ �h��q�L��[-u�E2��W�?��!}�e�Y�)M%i��j���[9�,)F�ÜǸ��� w��IU���X���b��KXAL{�Ņ��T�����'�����@4�(�&a�'�~_��? �9*n��&��&�+�K���"��S����y�����}qL����������F��:6@;����d~#fj��4���j��Fd�$1�l`4�xH{�S��	�����l��VG�k����V�f�Y�E�w�d07�0�r���Ĳb���4I*�d=����b�RU�R��ڥ�.^ḯ���O�89�_������;����������kR�1�&��;�Q��vT@�X���1%�{W�0�J���� ��k�{I�5}����������dV$��vo-q���Zz��~.�N(��l��;ӬM,<h��O�`���3p�!�o��`�ʣP��PW��5�s����|�ߛ\�I 12�I~���n>��m'�$od��{=^�p�ɞA �tQSk�;�:��#O-p!�/�hE�Rm��d��CS_����4b�|�X���w��Y�$��V�U�=!kJlx���]5�p����%��M!~� �(Xz���'E$V�\�Ԑ�|��lwM�+}V:��M��~
�1���qJBy�*oV��1��F)�P�%p*��j%�]��L�}�:X/j-�g9���������S˧�/~�`;U����� ����K��mMГ��������L�)��}�A������Q�[1������-��Q�6��~7����J�����Qv���,����X�����
��n�gM2�ӑ�-%�Cʫ@���D".�uK;�ĩ�#́w��(�:��g�{�M��#����*��Q���'��)�C���*���B�i�J3�yqB� �|Gmy�O��{@~�M�5�Gӻ+�[��~AL���h��8Ύ
���r^W��_�YY+��s���A.r��U8��r��<��RzÏc�
��挗|UF�Ȼ����|?�1�p�� ,w��߸-��k�����f��Ӈ5��grd_�H��ؙ��u�n0�ZYV9���;�Q���R�}�Pj8L��6��XM�%�61�$�E7��5ԩ7aB����]�]w�^K�i��b���]_�6�)pۓ?^��:n���w&��h�/�)����%�����*ƌ~o�(���C��H�H���L�4�p��*�ҝ�J�@_<��h��:��*W��
�T,�.����b�7�-�!ߞ@��D)�{��f�Ew~󵙻�\�gr�h��p��6/l�~,�!�D�� ow`�\e=�]�S={�-=[�x�P�H���\�ӟ���1��b`�x����С��[�n��<��f������Q���Ƙ�uy?�)�"������H���+�^�_��=�sn�,Ԏ�W��G7�^X�<〈q��92�9����[[,ĈEGLh*K�T�F�KVf�S>�S�l�hW>,n 3��q�e��0a�_mAw��f`3d7ɳ~~
��:���C)^�ߘ�q)=@k��5�B �j�/DDe��Ds�� �6�M+g������l�[W��-N�H�x�^+�RRUPo`y#���C#�ݜtE�a0���4���9ld��3� �����<1,����^�I�H�� �%k\n0�2��Wd�?Ֆw~����-	iD.�ћ��_s8�is��"|�J��$IwQ�;�Y�]�@i�U #�kB�%�p���бr��XM��X���j�&���Ω�Ǵ�'q��m���9����%�r:�(5�!L�r�G4��&��s �]yC�Pq�����+��H�������o�$��g�a������g�);g��I&I���ƒ-"8	�?jo��$,�v�_�b�Y��$�ɞ��>�;�N!׹�1R��%4��7o�CҪ��'c���	.InC��f�#��GA���L�pgf�p���wb�G[�b�K��oo���2@|(e�E��R��4��hP�&�y'�c.$����%����\�T$I���쾈�3��,=���{�Q���+��V���:��;eR����mᴚ����;8���1ILs>drȶ�_������co�tj�MF�2�F7�9_�q�ۥF��\{��}۞
�f�'V�k�l�E��:�jvh�M��γ4�3mR��_��M"O�b��4���W�h|��yٞTfu�����q��V:���*u���'�Hf��.J�u�|څMt�u�j��О�$*7%~�9(df�^��9)w��B�k�"u����!_Z]}�ѥg��UX�L�$�S���]�K\�f0��3|�h�:
<^���㑑ٴ�r��/D� ��M���`Ip�Kc4�M�'����}Ґ�$b-Ҡb`S5�Ht�ʺh<� �Sgux�9'��8;u��$4X�
��t�xz��E�mԷ�Up¤���-��w6�n:Ѵ�	���vo���0�ݹo���nص���4�M��Vn�axiQ��;�^�S?�nik����,`���K8�xB&�i� �I��B��}�p��"�x̉�2v���I���Uu�h�G�G�)�OxE���Jx�Dk����ʦ�F�$H>go�k�UX}��'�$v�`-��z�Sg7��9�v�F�u0�$	Bivr�M�(y6S!�\�C�����pd�r�s;Q�����t*\��\��?��l�����(]'C��m2Щ�!A�����x��@r̮����.�M�6Lx�b�F�X�[r���]�yѳT���SЪ����l@�%�
C ���m\"��ŨI�G�Ц�}�o[Y>d�Y#/�+sA� ;�!��'�6��3���p6NCyk��^��A~C��\�^�4.���ve9��0���I{"ó������BDI�\xAD\�Q�nx�����"��orX�g���Țv��D�[#��iDPF�\���i���w�J���}�9�#�Xs v��2\�;����εF�ga5P�z���6�n����mS��QnO�ờ9z�Ӿx�]���Z䮡&��`�����E�� B��,�-�3�P7Z�V:wsa�*7߾
�K�Ѧ�-M�Pŭ�RwgvI��V7l
�Is���"�z&~Pr(�c�f��}�İ�f���D���U���4�k4�l���l,���M�(5�\���<*w���:2��ބ+-��~
�8���}���P7`:[]�i�^qg�Oܨ���;Y|��!��;���Ї���;8���Di�p$&G6�L��o�����<��I����ӽ�����}�^�����o9K�<�*�W
�aK��E� �D`�'G _��E� ���Ju6�g���{dR��1�7�3�Y��K����k-�х�!��@���&�-��#�깍fm0-������Q�'�8�*�A
v/��{�"� f��^�E�i�]75V�ba	�/(�hj�e�V�7��P�%�~'�G����ʿ�^��H����./
��:��s��U���b�@��=*,}\��!B} ۆ��mQ˺��������NWS*a�Us���oCyN�ږ������J2~^��
*T4�EX�&�n\�p^xB�Y^�cP��jyf���D�0�=�W����E:#��,$��ی��Y|ԋn��A(�O��Y�Ua���<`��m_huR�$���Nך��^��U������Ok������.���,���&<�h�2�V��	W�HJb0?�C�o���ș���r4����(y��j���ig�d/<��6~��Ԙz	k�٦�ŵ���=zZ �Bn �֯fa(ֶ�},����f�	�����x��ׂ�7�������������Z��#��Aڰ�e�<�w ̣�2Ye��G[�/�K���#[=��_ŵJ��vo��5�˾�Pj���Z\��U���M�C�YD��FE[�>^
Gꕫ��8�#²C6�l�~�M�(/t��T�	9�"3X�E��i�2jl�=�!:�	|�A�����O����L �
3r'���X�F�k�'�W����`Idq!獮Xz�����`
�qf�>#�ңaq'�g$����s~C9�+��~��.g5�RʇB�]���}�tg� �%`���$-�@PP�F[EpI��4�*�������͑mz&�dS��Qu2�R~#j��(�O���4*4e��rC:i0S�Ql�Q���(�;�%s� �$�Ϣ%̛�V�E'�9�ĝR�j�"�8�XW�S
�[ ��!����!�Ǒ�V�k�.��l�����S�([��_/W�olg�@xm_k$����Gc���Ԏtq�p�2"bf��3�#B׋�mwh P��$hV�h:����rn�TF�jt��/�e���o!���7!���h0�X��!S�܅�ٲ(��b�(Ý{A�(�Gj/f�"b����7���o��WSb*�l�-1FxO�Zh7�N��5ё�]E�/���d+Y೯��;�N�E�S`��8T���{����HA,���Z�u��<�t���Q�C��NQ�Hf��UYy|�e�!~SA��3���<�����9�ˬm�9�2�uT�6�(H4w��ŀ��|�d�ⱀB�]HS�����|D�׃w���*�M���9�%W���,ɋm�rdǳ�����H{��Z���S5�ڂ>�^X,��l$�S�,[���4᜜ɛ�l�,0�!�Ԧ�4���FVn�������^$
����C�,��0)����YZG\��>�� {�^����X)�2q���(��[O���w�����Ȉ��S��7�h�����$�_!�(�q����R](�η��*�����:+��qV{��A���2������"�#d[ĺ�2}�q����dƆ!k�Hb.�.��M&5Y��\,�!��G�m�B�im�%	2~<��l�"�<<mO~P=�w����`ko�̮������K���07}x�yM;|DԎ���������ɀ�r��e^Υ�n�2��]������!.��/�k��D�x��������������
^^�t�� {�B�G�3��,��MOy�n�a��MbāEc��#�+�qj~
Ȃ��Y�R|�s�wv5�B���.]�p
�@����l�΅�����"*˚/_i|��;1����Ĩ�pJa�F�<��b�u4TZ�lQk�H6��Hu�r)���JZe\���o��K)��PÜ��ד�tE����/�Y1��+�ͼ�*� @_�DT�Ye���>�٣�>4c�%�z�����ґ�{\h�Ls�L/a� *�w+�<"�c*�-�K��f��)��"�|���>�m�N ��O �Y������Ky.z��8
��Q#���5E�5l��'�2�C?�T�z��^���&���n�0���f3<ܿ3����v�KW)�|�_�R�'�-���m-�w��v���uO�t�l��.7���[[�0(w��%�@�iI��`V���k�JdTz�<���q�o��nF�PoONM�Ho	��,L�%�6T�l]��U����|'���³��m:�h\�AG��td�Í�~�C�b�ˢ�֌0�v�A�	�~O޲�ޞ��>S�Ȗ��R�MT�9�!6D}�2��E; �dЉ��gss�O���]2�Vhj���7�8�<��Pw����������6ް[I	�|{k-��Z�"҂����5�_�Z�`X&o?i���!h
��4��ɏ蝹Eo4z` �(�K#hP�fv�Qѷ*?m۶�����*Ů�����w���r���P�PX� �قc���|2I���K:�*挀�Y��N= �.����@���`�"wg��3��anlCS��Hov�et;Aҥ��N�,�Z8�����x g[��ߚa����]�S�b`�^J�1ݼ,<�B��bV�h ��p�bҷ]�ƸY��#t�3h�� ��u`�s�] ����*A������IT�M��\+Ks�dEK�j�e�NѷЩʐ1bX���/�#�pM�sy�����M.-^��%A�-լ�^���g-�x�Ef)��"	9#��쎮k+��M�ӹtss��􊘜�k����rɑڊ輋�m��g����3 
����sR�P�DX�f�7QG�7��#u+xoЭ�����q���YKzE�;��C�⢊H���R��찚�)��)<��,�l��׷ZtzGV��T�b�D9������N׆M"m��W>Az)�M��0i�!�x"ɵ%<���aX��C]@f1 V%x�(L�ch�pMۼԪi��&���OP_�Ű�[�X��׈�/ClD�l#.�V
���ut:�
�u���
遖Y�?���,�x�w�%�� �9�Y�F��!��]9��uhU�v,�<qv71�_�7QAW�R3>>rbi�gxL�9��
'Zz�g'����q1JSA���~+N�]���ʶ��B���3��ܫ6Hԥ4���%ɤC�w��4�.��R��i*d���D?��S�d����M�%�/T
ʍ����u�ȵ�{BHXb(��ũ�����#��<��;C���}�c����$�ϥx���f�j/w.LuyXQ��rC����Y��'�%��Rg�~D�_��I�	�V��%��-�!� {V����H#��t�t�+s�������φd!'P�l�3����0N!�g���"z�5��䑩Ώaxi�F<a8�lTҵ�����:�hq�"+9�>Ǥ�ī�']NX�,}/'��\�`��r��4�9�xz��ܿ%ygl�&5	ח��k��
M24���O��	��dܕԙ/|�^�/�7_������+R�L�O��kCcB������9-l~�/�P�c E�,�ue�� Q���r�>-_��CbJ";�{���?J'O��-��E5�)�z�+N����罥>z�jsY�#�,�~��k�E8;{{���y'm��Q��B�)��2R��B}y�����j��&Vn�i\��
]f�xx�[�!:ڡ0EUM �	��7�.6�u�v"�����y�02��e0 �;z����΄k�y�D�c���-����"lO�.�oA�~�Er�+�a���w'�T���b��\�)$_��uq������+�S�u�+��\K�"�d |%c_A�ӟ�	�ى=�^�ե���̚�'�a�{��E��O8H�5�3�b�g��p��ԃ��~zl\V�]&A��{C�J����Ed�ءz������mD��3K�u�e}�S@lkMbT�Ǩ���7��>��5-k=��B	�z�NM��{�e�k�hj���S���@~0���4]E�aTOCv��,�#��H�3�����LXi:��j��S����a-h� ��č��(�{B�<�D)Q�Rm�D�@�̊�a/�8�d�/�D�[�Z ���zZte lm�-�����B�i����6�O���c�����Co�i��Oð�9��H�I-$��E�3řj_x��������\�����T�n���$||1�A.>Ĭ�й�G�Q��v?�G�5>7`r��?�ya�Q�$��%��Ks�[�x�=���gJc#�R�o�{�ϗ���]V�^�ZP�^̅��UC:��=��9B:2�+'w��Exiȫ�Cu~6K`��E�܋���u�F~���d�?���U��G�悜�IF+��(^:���`���,�ZM!C��\R~����8^���3�j")���$�~.ѾG٫a�vyd��2�Y���L"Oo�%'X;x��x�<���\N�QR��Xfi��Ǹ���j~��rt�}Wq7�F�����.��� �䌥�b��[��I��:��Ur�fxH���(k���û�A��.�5��U6l;m�(f sȭ+T�W����c�~�N�G��O�,��@�_��5U,�'G�Nɠߥ��A���2���x�E�_�S����߾
�O�x;��lR�c^�-�p�AM�ɡVl*�D��\zP�QC��/pf��_�U'6,��}4�B���(�g�=�����L�Ʈc�#L��괢�a�i� z�$��Nݠ�o�nf,v�G2��#=��P���he6a�i��;,ۗSL�]|iP��M���43��=R|
��/P���<��a�ᳮu�~2��g�� B���b��^����C��y4��	�;54k�b�����)q���1]h,Q�c���q�ե�P|F|sB0�'�(\�v��3��%�o���{�`*M���u7%#3����]cu��2�*M	|t�h|d��z����h�"��Z�%z`��I(�S��5ٶ$6�8l�i�o&�Ƃ�u��_A�op���9m�0�5�����L�6;�۶D��2"����M�P9n���C����/]��Y�P������=�1�,�#%�i��� ��ɂ`�:w�r��4��n����	��q��|QuT�����;�&!��+$��*u���N?	;'9S�Æ!M\y
*B�Ҧ�i��/�!��<�Pu���i��z#7���҂	�g߻M.�/p��4��wޓ��!�bS>��6���I��"��"|���YL�`'�1�1Q�-���⻉nK;�[9���yG���9Ba�1~'m�}�oX����<�HW��%C�*;A�b��p����zبvW,y:J��8uI?
Lu��&�Uc�؞K�!����B����.ҿ�FmtYd�S��3��[���&�������~CN��z�y�tm����Ysg��=�ت��^��/;|ҰR}%�(	.�����ƾ���Yu���dXy�hl� ��}Ϋ,M�f� �$�;�D5���?����n�V+J��uGZަUM�~W��BQ��ˮwCO*_'�S���T�S*�u�uzH}�^�k��ۯ&�o�`ˠ >7��֣5��7*&(㵦-2>��tW���}�3��$�l�$㑩C$����zN�+>؋>�sa�w�����|�B��Μ�G�#t~%ҠQ��/Q\�p|��'��QΪ��R�7x�Z�s�6|��Bae�c����Cض��qO��ſ�-�Z�a�JXe��zSܾ^=3�5
�W�Ě���o���뭜z�H
S��O߀��~�!�I-߇^<&�V�T|{�����d�>	_܍ ���$U�M���������y� �x��ޗ����X�A�ӋSޅ�Vd)	.0�@�ߣG����Q1���-F�f�5�ż����nf��1p��:��_Ԋ~4�b�V͕���U���so a��Q�W3��$[xŅ��v�TW��u\ʬ��T�*�x'ǹS�^kA0����Wd������-�E�
�_�T\8G�P�mf�%�p�;rk&����>�ex�+ �W� ƫ���}�I+�(���"�=݌9�p��+l���Me
�������t5�9�{�3�(ӏ��Cs�R�x���1&٪ HYW�\A!] KC0��y/��x� ��7��H���r��"�ii��Y~���5�f`-s=1+�a��6��>�8��b�����±ea�kf�Y������Y�r�������z��z���C�m�X��Ͷ�0�A�dA��3{
���h�U��blu3�텄��"	��-���(�T�!�D`�-�[�Qw�����f�~��>��Ń��o�E���	�bv/�|SD3�kbs ��/�p�P!�u=18d'OJ�.DNM���5g_�I1z�����/��,���ĀO�V�T[W.؝��<Z�����C����u�#��PS��Y�q,F����٠A����9(B�n�+F���E%8ʆ�v�/:QdJ��Ȳu���!!c�-rM���ք�+��g�VgY�&a�؏�7m�F��� ��R��6\)�nz�l�>kT��M�Fม9�E/&�2��W���B���=Z��A���2�>:�%�X�kZ\6v2�%��+yX+^@Tj.�˯����\�XZ�BS~�n�p��v9쫐�˙�ɻ!� W�� ��|p�M�)ͼ���m>��5�A(7]!Y�ʈY����o�R|�H��>^�U`ԔJڟߎ����|��fk�D-[�g�����X��k�T����{z��p�����l�����6?{^K�_�����X��.���U�x���L�/qj�P���W� ̜�z~������9��^�0����2~#�cnm�}|����T�D��C'w2���wb��O�dB����nnD��w{
�o�]�_�\�AKy�X��V�)�h-��5,��Х_]���ӢK����V�!u7-A8Q���>7��L�p__X���up��L�Ѩ׌y�5ʂMd�R���LE����n6����g�+`˴�~>�T�/x�&�`����M���H��\��=��G�tk�dk:�C0rU6�&d��|���]�,o\�	���վkRY�Le��YoM��>,+X�)�[ ���A'"��N��3GG����4ED�,�FʥɳN���-�q(�0Z8Y���%A�_x8�"���j@�P���z~9�$����
E�J2��Zw�ż�8�:bV���(���2�j�]$\��]vʊٽ�DV.� � {WQB�-�~7�߱�<���I(\��-u�����ђ�1���@Nu��e)s��P����?r�}-�p��'G�ŔD�����!�x��^(�z��d�0��U6����O�hC�j�֮9ZE���0yݼ;�f�]\�˿q�:�<ס��@)|H9�@�,-�l�_�`�e�7���s+���r���L=7��M���� r��xsr�Q�S����^t���������� �{�G'�QTp�ͯp�쭢�́�@��T=B�D�u��(��`���nk��k�\��Q����������V*Q ���kMʳ�:w�A�o��nnbϒ�{��65v"?���Z��Ƙ���w����Ni�@G���.�7OU��x{����;�B:�[�O6<ә��#�H�*%s&5$�Z��ë#V��{��٪٠ـ���9�����
�r��VҨ{��{AK7Mղ�u�\;Mtr��Ϗ	WS��O2�*ncʝ���Pԝ}�����!���[�#W���}��<V�r	���nx��ݠ�j�L�c-b�[݆<E_�U�gM���oJ�7��B���Xú�8�E��X]� ʧ�l^��)��؃�npY��Gvl_��Db�~4~�.e��!Gh�a���.Z��{躗���5��7��1��uq&ݍ�0l��{�-� z	Ax��@ǯt��Q�N@���n8ދ8%���y
i?{l���3[-��շ�����}�>���ށ�̉3دM����+��	�ej!��-1	��	���h���.D-��]�C�$��Uh�I[�>�ФhU�w%,.�|��Vn�P/�&���6Ց������<�t����L0I�NO[�0��(/���ݽ��8̌t��x=��������᾽M�T���>o�߳�=��^�[Y�KQ��s}��tA����իڽ�dF{?�i� �_=��q}8l�=�
+�&���8�Ȓ���lݜ����k�ϭ$����Io��J�&�K��71�������<~<�I:�"���N�]D��0M膚��u:r�7q�0���0x'��4c�0N���6:��X&��}�|���/9ߩp4N�����Lm�	�!�CT̻bU.�*6��*���03;�x�앓pE��f�����q3���bZk�	��$ͅ,f��;&o	^ݘ9�z�>]V���钛��g�P!�U$���c�'{zZ]�r�!��w\��]L�Ra]���� o4U`�E�s����lO�F/t[�0k�2&�]m��{�r��Cb/r���<xm�Q�y-i3�Lq�S�90�4`_�+�W�\w�QN��d3a����/��3<�`���N�^Ob 7��L����C��u%�����q�.h&�x��H����VV�z����k��`9�8�Xx���'�TNt��yڛ��s��w^�X	"T&#�����o��܅�����Ay��{V�z���-���[��������J�x-��]���w�h/�qI�w:���m7�B��������A4Xp����4��y��]�K�t��-����qw�W���j�2܈��ݸ�5��[��*/����M}GD@��%�`a��[jHy2Ɔ�*є��x�g��Z����K��׏��SQ�b��1F�piI#��hESJͺ�0��c8Ue.Q��I#�#��҃8��� ��1�&��m�j�cr�ߌ�' JϻW= ̬��VJ֘>�g!6�-5�zj���a]�Po����{�f�W%�t\$��Z����^����{,I�w؍�0,C��x��f*|F��w�fzxf���z̫�����2%�6F��m�+1�i��[g�w lNEYF�fvYL���q����eE����g`�8b�ں8it��%���	�UnÞ�\}>Վ�Un���v�ݸM[$L(�$��20�.�ı�J�~W7�kY@�>ƣe�Q��uG$!��+>�#����2rjx���;�+��jB[y�\�c�VM�P|F%�!�BZ� j������0�3��LxS�e/����(�쌣}����t�.��C�k- ����i'|>�1�7�je��$����ΑG�D�V�?zf�ܝ%�9�{)QG!�)=&)�=�2�[!��g�ƀ̓P�?D�S�1�zE�@*���:.���EU� x�%v��99R�gs��@�J��V)�S���
>+����Kͼ����8���݆;��DZ��z�9t[l�����h�_;�|�A�3��]��
��	Wt����E�h�_3$�ͤb�qQ�����h��L�91�x�fǵ�z�{�C�#��=�*�JVfs
m�C�^,��ޓ�;Sj(�/�;��4w1W̛-� � @
��@�>5��:��Q�Qbmo���`sp��g��� R5Z^.�y5h& 0��J�+'��JS+��)�ҒT^�=�8x�+�<��đ���,T�!���2|����1��3���ό������C���T�
��E�9����ˢ[�`n�r����R���H���4h9
�_=(-An;���M�z��@��ײ}��[۪
L�P��h��Mݭyo��/X��oz��e����/�ZJG$�?9r����f��D���4K|$��E�l�*ڙ�nR�h�s���V	I�~����*�.$�Syp�50I�"Q^.[<>�����C���C�4z�Qn���Ոٕ��<��x�"g��	�|�ꖵ��c�F�o� Ә���:�׉�����м
L�T��a�����x�h�7�TV�Fk�8��د�DQ��Ba�1Wi�%;�:,���b)3Cp� '#�d�����3��;8D4(�GB�Α�gC��O�u����`��6|{͡�"[�;�������QE�]$����fLJ�����Z�9j����*�A'~B�پ�;h��O��h�����n�u�jVw�l�v�*�[����G_
�]�S�+7��/@$����M�zᖚ��6i6v���`���)�~��SRɢ�|��$�z[U� ����CӅC�/�l�'݅g���+[�����st����_��i&��bj^F���}�O�]����fJa�nYw��`
o�@�x�D݋�d���;�b�-;a���e�G��
BaP���:�t��\T�z̈��n}#q�B���tϡK�(�����?i{u-ַ�}�˳���!c���'�Ҩ6��iI�^:�|�5��G�ue:�4�5u��TA��ΒoaF���Z���\��;�(���v$	,��HI���XD�q� �f/�0O_2��ZD�t�ft�������)���������Ezd�,}�Y����m�#����u��E���݅��m;�E�k耂0�O>2W�H�� ������+��XAХSt�F&;$$����qB�y��s����h�� Ip|ժ��
5�=>���a�]��Vˇ�.ƒRP�R���/P�v���h�:�0����#n*v	�B1��7�
�j8p�s����ߵ!l���S�Y�˰p�<G�٭��jl�O���&�z�-!5�*l���!G]���ۃ1����1�c�$�U+��tW�,qR�_�kea�f�f6!&%+MɌj�V�^�XgY��!(z4�%u�M�e�u����ف�A=h��CokN)j5�=�M���\��gt-J"�D�XC�/�4�!� 5�Kq�k��y�����T7�u���^e"9e�)��� �W���R�]�\M|,� 7��h�>V�5)�D���pb��#�1E��� 6�V)�>'8x�e�f�����Hn�u�Ak9"V�=��$A�J��S~�1Zc�#r�4�����Q�]�Q��Q�V��m�������tdlR��k)�Ɓ簍eZ+�eK��-�C��!��vD�&R
n���%贘��G�s��,Ѥ3�^��\ۙ��D�0=��eu�t��~l�1�� dԣ7�} ��T�i�ԧ�����<\��uI���~�{����K�ǹ��]��%��r�,�рK	l~֎���e�H��*A�U9>�p�P�۳�d�+�*~�}���
VQS����!��3�	Ռ�}�#��۵�URf*}�{hH��������IY�5��L� �J	^�L9OJ�3�25�|V0�|t�vA�����c6��FҨH�uf	�J9K�ԁUm<W�6��Q0:��v���o6����:����r+)uyŻT����3�����
�ַ��G��:9L8��X��"�V6��kB�"���J�(�$��ϝW�OoO��v������v}�ɣ'\˴L'��X���O�(@��\d�pS/,�GI{��C���!`v��Ҳ1d����_խ	d�� �7�!�I�\U�݌�S)�o������C��ر��C��K!����i���}h�DǸ����"S�ܛ�����`����=�5\d{'~\�#��f��������wY��	�1�="篔�k�\f_�^�um��a�Yz�#�>& L& ���(N7�3~�e�u�vqE�"1�A/�]�T��y�-0�v���˭�'�eR���B�ȱ%@j:-2�E뮒8s�	�i|�$V��0���2�7�e8� B3��j9�w
z�?�]�r��`��B�Ku+̋���R�X5=�ra����'�(�I�<p���1a��|�ͺ��M���:�������RƓ�$��#�o�rd~�r_b���1V����FP� �Ѽz�8�˼�ZW(@�9P`Y��A�Uy��0����Y'�
�l�E*c��=�u��P����F������$��oiGw�u��a�	]a;��?�?��(�v<��`g�X�1���6��$wS�l��\�R���ed[��3jr���U�2	�g�LHt�/� lCT�+,�ӥ՟����c��#��+^����������t�>�5��.�~��m�=��࿁��}{�R��APM�d�N�m	�����'>�P���Ef��AJ�aCos�Y�n��=�kK���5��Z�0��}��n��3c7CQ'�V��~<�:%%g('7�3̪C믜Nh��&�FQ��-DJO���x��z��N���	;0�1�P߈cn݌��0��,���$��S��ChnU�j�ebhq�U�?�k��(G�3�z&�Ҹ��bNg��K$�5�p�����Ǿ�x���Z�ֈ���H�%"au4	6��}���Joy#�ș��9��Ek��gXc��KE��'׼�ÌǏy�X����\�?��գX�9	�k�^Ԃ��Ń �U@�Qei6i�?{����nd�m��f�CKۅ�/n`p,ϧ���RC��%�H�C��]�Th���������'h7��I��A���ŕb:&�SQ���+*��q�S4A!�]�T?�8�sʳh4xK�(O7G�"��/r-����([f�x�3���_�=�\A���c2�������ƉQ��Ǩ�k{T�2�Dp}�J[�-0���$��x��º�ݪ,��]�B~���"SY|N-An������Ό�ԕ���C!ct{���%oT�,�����o�=��gΩ����_6j6���\ԩqpxWRF:v��"�ao^��G�$7�k���$��}C������7fwAR8��[��.�����KR���M##���� ���^fO�>�����^]�ij�^<���π�n]˶8sD#s���zʢD%��9�%CۿM�s?y�!��'�G�I���Md�����o��Q�A,;"��2k	�-�������X�F<��d𕱍}�V��49̚��#Ӽ]�^y9qrqg��qh�I�Ć�vj	J]���^YD�'�N����ј>j-�{�2�7m�`K�O1��QJ�v\1c��;G�"^S�i&y������Ă3x�|;�:��h��-��{��FEM��������m��`j6�C�bN���cgx��֊t|em�s۝�d����c�Ju�1=6�"��64~}Q~�y�/�sB�ky[X�]5�Z̧���!���eQ�� Ʈp#4b#ʻ�i��9q�rG̨}��E��&��>kl�՝���A&_ż����$��"��x�s���{�9���=������%�:����J�5�L٨ȶ08��5�B�r+���[_�Dc\sH��_k�sa�#^? G헅���������?�$<�&���R�9	/c��vG��}yO�ּ��'��c9\�3��H����^!D�O)P B��Z*�����QL�{\����,��ǥ�f}J��d��.��-ݧ�ճ���?�d�>�5{��ۢû����'T��(���MD���:�}] �&�n��@�]E��m�1�s�a�Y֎�)��{ ��I��7\/)XrZ� ����O_��0�g/}R������q�:�'�@��3�	�LT���Ze�Z�i�(��E������(Xkt�*�@�pĎ#�&��c�3ۅ�PSo�c:|J����I�v4��4��8�	y�|ZA��`��{�����(�ܳ
�8�hry�v9��R�P�JgQ��� e>�C	���� ����YZ�B2���ڗ�vN��>�i����8��E}��6�B�k�����;<�<�|%Dvn�hj�ۢ(q[���w��&�,��uI�ԋ �Nr�"�I������kd�����Nc׎,>��;��K@���X@&ݹ���&[eȎH.>��M|��T�@��؉��c�M��I`-xLA3>�M��S=��q�q[n;���W��<����,��yPl�Q�r��#k�F>�Tr���X��FJ�I��Hr�x")�<@��K�2Od�J	�bG�̈́���+��P��xف�V>�]��1��*�!Bjn]ᵪ!�X��\~�6��@�����s'�^����_����~�=��zl��<�NI�
~�Y$MԖL���-1`�s������9�[w���ƒU?!�&^1ve�1=,[���(c�sW�r"WA�21��6��a���h��"`�E���t��K0S6�6�
��!�rG���1�(��JS���)���B���V�kOl��GO ������!��B~���>F� @V���ѸyP����a�k���p�}��Z��0�r�7Ɠ5�"��h�K�ņځ3�z>-y��b��)BҦ�\Bc���
J�����ˠ��qt_t�X�8C���uW{~}mBQ$���-��LG��jV��{$�#�8Y�}�^U�9��9z/P��ֳ8?��Q��{u�X+E�>��oꄝߏ�4徟����=�i>ݤ��5�+��J� ��N�ե����M��2��N@�Z�0G���n�����qB�K"��GT1�5k��>5M�Ks���yW8q�+��d�ˎ����τ�/BD�)<��K� ��+w٩�ٌQ����h��:��E��{��ak+�Nχ�2�î,{w�y���7e��Դxk�㵞��LW��8��G��w�KY��F�ղJ���]D�Bc+;Ȧ�{!G]j4≥ֳ3�����m��b3������d�py�r�m�����Zg�%�c��͍ʈ�̖T��494e��Σ���.e�{����u�k�b��ȉ���Ӵ�-ie{��ŵ4��B���ž��R�gB�4O	)�Xț��t�
DFG DNU�c��������~'I܄m�C����!�^�m�����Q�v mGJ7��~� X�g_�H��e�*ɘ��7d}F�O)���-�$t֠�)��>U�#����Nx�9���WaT�g�5�o�ڙ<����4q^H��}}��']��ƃykQ�����a^��m�5�/K��_�M�r�o�"� ���7X�Shx��ke��}6ے/��6x,}Qb��"��
�� d�'jz�2SNl�QL�F�,�
\�z�	��J���k<H?�D�M����`Ǌ8�ma��7��%���J���"�2x- E_��m#I卮�c r���Ϗ��Yw%�0�N\v3��.��to�R\)�� �v��������3H��|�DK���Rӵ�9N���D�ܻ �W�9Z�RT���w!�#6�w����Z�y�b� ���xxI͚���
�Vؓ"�1�ΠC���gcH-�635�a\6yeZ���{~�"���{j�����̍ݢ�bq���P�2c_-�D� ��f�v�1�O �[�j~d�-��^�jF�.$�]�N#k�M��-��n��莗�gs��A����e�=7V�	�I�[�sIJ@'��w�k&$
7n�@��w�	����wp���~c�c�G@fMS�e��7��*�S}*�p7c�&f�w���0W��~ݾ�8��'�^�ھ�0��s�v1��N�u�|S�7��:����9w��V����A@Z�*��hw�=^0|���채#� ������K>�-B"��E�k� "n� ��2v�^��r��P�f���[�����{x.�f��*�Vp�~*� �)]���~#h[�H��jx
_?����A\�83�.��Ā{l
�jw+�uA�/JP4�(GY�$z�x�hN
�h��-.���N�TP�����-���Z�J��$�g|�~K픉S��1��V�7hp���%��O(����2%XD쭛d*�L0k� Յn��]���f��������HH�i��m���Z����W 
�-�)4�h�d�@tqI���O�����ԅV�H����0FS�,���@2�����D�?J�c����d��{x�NՊ��9���ТѪ9�+��7��C��쇞X(�Ԣ4,���?9YV'ʔ(s�jp��?g~����)\\�<G���� ;�����J,K�QV�m���V>����\^��7)���y24�e�f�r�p��ئ���}i�p	����G.)��u�j<�(��T4,8��GO���Ӥ79��+	���`���1P�*�"�u�V*��������Q�p���ue� �������e��+;�V���
d4��QM��E��Y��JH[_;} �H4���bF�~�n���BJ�du1�5\��)��L��@t�ƥ&2�7�w�|�K8��Cb]�il�Ò�h���?�Ha!iG�<�!C�2�
.廁 �#���=��uV���N=�k[�0d[��2.�$\B�ߝ�(��BYE���G8 �}�7�ϛ	(�#�z���W��b7�h�.�6�;{0B�pt^X�.H�59M#�<w)g9m#�N8�@Z?��� ��^r,�y}Ru%���,X�{���VGOY�������y3J���\" +d�
ڳ��pAy�3Ťh�H��,l��� ����#"XV��"���U��!���A���RQJ"�ز�d�$�����_LÍ_2�'"���yj����>�ه���lj�TS'z�� � ����@�S���R��6�����4A�dN����	<�\��`S��h��������v�8�@HLv]�k��vHy:q;=���6����祥�9�f!����Z9����ֲˁR��Q��I����]'5X4���ow��b�&K��9�ʜ~����j,>�;\q�Q*�Aw��ڄk�+B�HXZ�T���@� 7������Ҵ�E�{sdǦĎ�PP,+�����;��K}�*��"6���8T%ZC��������3���u�|����*?��G-���sZ]��Pc�t���<F�B�R%Q�r17
�4���T��^��gi���Dl�+��-�x{H�./� \5��`�0ne��� Q�&By���dj9�0�-m���8"XHm�3F'ܫ�M��T �2|p&��[��ke��y�0']�:r�`q�7��HX�d��}F[��ǥ~J���q��2�F�q�?rt}�(��!�%��
�Mn�Q��O*,G&�X�/bdd��,R:�BN_�v1���m4��`��4��=�n��܅H�';� ����)���'9C��}ֵ/
D�l ��ת+~�Z�� �_A��2`�ci�)��v�)������s|��OƳ̴ͭ��KMP�U�bǲ1m�c��;dd�h�#��B���1�B�š����҆��4��'�P����Aӷ@���z�;�~�PH9O��R4�G�0��#2z7���/#8@w�K%P�r	�<~�>��]���;A{5d�f�R�mL��K���ď��i��t��"�S�,���'ND�Bs.�-\p��U֛J���99���j�h����0�`��a������偯���?��K��7�s��V�"Q*�2�l�v7Y,����Km�dCc�,����p��5
<�������*۹��r������5�����G�fٽ&M�B������U�]p��%?�n2����P娤8�x2=ʹ���j��4��L� �q+�_-���ra�D����/�@12���/�)��m����'�F��ӰY��V��{꠳t	���F.先�<�o��~y�v2��Fa<TT�I?D6WFC�t�JNd	��a�N:��9EM'�P�q<.Y�qy؋b�@>&�2��f�n��筈����K<�L�	aq�z��#d���:Ч< t���fH�ݟ�b�����"jL2�g/�?�Q6Ni�(�EN�h;͟Y��W3	"@�ˈ/��$	�����.�"3�r\��?Ѹ�aȿ�ߔ��1���5Vr���D�o��Ο�K��sbMM�k�t��jA��5[�N`�u���'�A��HO���6�lC`�t�\`
F�ɖp6����U�����ˮ�Q�ُRA���˦;h=��ٖ��f�Ҿ�"���:K��m�oU9�G��
#�FMP���.�!�� �����ӏ�)I9"�t3i��:�ߙ��F�pj�����b����x4,��w���ȳUpT�R��e��w��z��$�oG^%g��Φ�e�0�QƓ�H~��iS�\�&ݍ^t�҇��7�!C����߰d�	���b���rƆuMP`{�ͥ'�Q�|���+M���e�=�w�r92����|�/��R6�7TyX�kw1��"\v#tC�@������M���E�;.��`�6�[��1}Ut� ��s��-Mp��M���� �f���4�n��6v�S���<������%`G����\޺�P���Eҵ�� ��F�n��l�aB�]�S��Db�O$�Kr+@(� {����o��1a-�zj�h���H?D�4���iWqFq��#���i�K~���tS�f����n~b�Qb�o�^�e��fZ���Zk|������ ؕ�Z掙q�}c�>�]Ǐő�>=~�P:rFM�mͯ�$��?��Ț�G��=͛ϖ*��6,�}����IF�6��(Br���m�zc��Y���OY���Z���o��O�t@"��������CN�Oy���>��R�E��!'&�f���h�~9?�{�
�P��̴��o��`9g��.�pm�-9�X�Zq(�E�S�������'E{������h��r'���~`A���`��P3_[��!׽W�κ��PZ6�ի"��=\ ��G�����u�zي����o�
<�u��%�z�Ly>9��Kq��1���������VϠ�y��h�.��X0�?�y�*\g�a<ؕA�ˆ	�i5;��U�"���#">�����qd��"�>ݢ��cZG0pa�ı�u�-ɦ�!C�?�M�����U�Q럊m�����=M��Ǔ�0�*��
�yD�0��Q2�5����j��|�R��M�S�� :u�����"u��U�p�һ��Kq��6�{R�:9h�b-2�͛�r��J����sڱ� ]Ǫ�e���v�@
T])�ʼYI�L���S<'���%Ÿ��g�Lg^ ��]"δAO0�
���{Ls���M[2-)��@�L�;x0�/���~���̔�L.I�-��/LJmf�s��{g�@�zO�_����~,ϝHj�[7�cCXS}��'�6�>�C�Z�I�h�K3�5�XL ��AT+is㎷;� F�g+G,j�L<�C�BW|ƫ��Y���8j����{�C��J��`��}S�A�WE�͖��zѭWM���<��A��@��&b�%���6��]�Lw3n;�]��pXY�����x��8�(d�0�|`)�� O2[ʠ0{Y	,�M=IGr0�����U�т"P��zg���̓4g�f�3���&U*]�
�Hp���z�HN�l��i�w�,k�A����g�/�R�lb/�:�K�6:Jm��o?g:��(*h��وx�0{��X��GrE��_���"�\�����r��0�TAU'����P�7*h�n��m�Ù��3c��vtq����U��V��Z���1zLLGj��%�O����# �4"T*��_RvHGYZ����Ҁd2��#�g��x�[X ��j��8�^UK{Q��5">~�|�X&��.����\�*z�/��r�W�܍���!8S�[3���k��l�K��nL�_���|�W8��Ih�ɪ���1�-���}~M���v\J��O�hj����/�T1�Fe�M�SK�KΗ�֤-��f-D�)���f�Y��0��/ )�J�]��PFa�������H]P(Gl�}��<�W��>�zL�ӄ��ͣ�l#��>�%�iӽ2�l�����e��ͪp]O��rDt�su���s����2i	X��D摖ޢ��0�
���"�� ��ޡL�p�j
�3�	��LT	�xj�B�}�Iu͔G��pK�O�t'2YS֦O��AO�𼑮���1�$^]���r��+�d#��#�Z���� n0���Ŵ�������e������^F|�"ޛ�| �OIF��}�E�U#�,��֧���
>�ؤ�&p2�	�h����xQmV��Wǁ���_5<�}*X���X���f��f��"ŭO{Nj�V�Auo^տ�nj쒆�D�A	TT%e�v�2~�taV|��V���t7Q��i�44�=I��Q)d���Ub2�V]e V��x#t>U��F�j�#l(D�h�*�S*�T`����k��=:�?��m�C?	vG61�V�0i2>`�oy����v��f�m��]���]��_��m����l��H��~�W�K�H�;��qw����G#�Y#]C	D�-<ߘ1A&1|RƆ5x��+wr��Y�y�O2BM�g����ɍ^�A�]֗r�1�<�X项}���DNș�`.���d�߳�}QD�_" :��ųN�T��r)�t�+k15�ˮ*α��aŲ̽Q�����S�aA����v��׌�qVK޳�0փ���^>�M�m� �F�[��a����mxt��DՃMFrof�bA�6�TiPF�3W�eH�vu��ɤKv�F�)�K"��_�����;����ki�n�	tu�ͲJy��g��u�xz��h�A�"�����aEZ���c����0��B����e���;a�j�/گ7m5U:q$���F�3=��u9�)���2���W�GX
;3C%=���3�6B�έ�����+΍R�nt�0��5_�qԛ�r���t�m�e�;��-a����TEn��b5S;[�5+&���2Qth���8����(oސK�x����N���P!��?�o�������P���*�a�"j,~߷��
�bL�1�� .�.�ϝ�ǜJ�jbm�w�O�+�<�����9V�+tZ�j�%�p�����F(��E��*t��h�}|aO �
����N���I;�L^\�Cdd�"�׾>�GR�i�-�X>���^xj	itDm��$�ffU�m�ЍA��[ҹ��ʿУ��L��g���F��GEP<b�(y��Q�yX���?��w�	�m"�hN_|Dv<⇞��TF=��;��i,�X���Awr����J�%U�)d���:s:eM�蹡��9USd���w�0̌��xd2ࡣ�`��p�,�b7���{�t_)������O ���cz:���A�X�:f^背>�ӟ'�`~���S�p�zG=����w�j�~��B6T���<~@.�|�ެ�o�3�Y2���\m�Y�m��Z"ݹqi{*�"+�ҌĒO�.���+PX�����b(��;�7�RX�� <�K��uQT�f��F����U�Dx�e��[��Z�E�'�YD�`��i= �Ք��;hTT����2p�����To��mZ���'-uu�Eʣ��K4�������sA�o]�j/%���q�B1�l���D|�����\�dgY�sPA��W���nrW
�@�,��V�R�+�It�~�{�M)Uh��)8��/�ГϏ�R�	����C�Sgp�W����S8{*49H�T"����OM���U��?�Y2�3����َ�fO���yg�z�tR��H�Ǻ�P�E�AS��y������3x�_y��5Hû����u��j0�k����8�O�9'n��Կ+'�d<3���I}e�����~Q�D�Uȍ����iJ{�B�U����G�(���A��͑��-YO��j��������7(C-×��4�;�&�����V��O#"� ҪJ���D�a�OdR��p�e���s���%+�h	;wӚ�b�G�b��ԩ�F�o�VRΩj+ل�;�%��L�3�_i��9ZQ��Pl��ཛྷ�*�~�:|���y+���z9r��Ax�l`���d�#�H���c�D2H���Y[]��/i'�OVL~sZU7�uCdY�Z�P�4��@v���{���mi}������*	�sy*Vs(?�W�}�v�J�eg��~,3ܢ!��Ӯ5��OÐe+|������ѹ�>��W鳥�y�M�c��g���P�Q��l�C�	�� �W)Ϗ`L��_��z'(+���e��������\�t�(]6O�����)�@x�C�o�.�kB�`��u�B�?�N !��&9��L�6��x0k�րp�H�%:^�:�X�F��˴x
OCڷ��zf'�q�y��QS���a�Sl�� ��kj�5q�6db_�O���$^z��]-�KZ%Ϣ����c����m�^0���ꠢ��� ZHK�+:ZS�S�,l���5ysx�t�g�/�h��P���$z.��ώ����Y�v�<�_�j`�V|����3J�X3�sD�g;	�^B�!�A�W�r�L����Qҿ�����ӡ[�q2\9[ֹ��̠������He���h��%H�Yt�F6�����>�hY�I�a���;#`�wfj����=�Z�S��m	���ľ|��z��_I�׿iz�̏7���ŁUi���x+��xQ(B�J��k��G
z�-I�,�q���ś�j������k]���6��|����WU#���H�A"9����)���GHw�pҝ�8}��0:��F#�$�ר��H"�0����ѡz�E9p$=;>828����WS�]��:�E�I�WkpH�WN�Vq����c�UM&�G��btI�^]�7ּ���9�VC����~��$/g�y
�;��n/������zfb[��ZL�F5d�����p��*<~��+��'��h�S���ہ݄��4+�� V���)j��M���\QE����#�W���y`�{�0�e�����9/^��b[��b<&Z���a��Ǒx�����p������s	oo���1Q�[m���o�� �����tz��Jd�l8��!�+�>½�%��g��L�F�!66�z�|O�)�����ğ��>~�m��H�%�ZF��Za�`ʓ�房\����ʧ'O�@�j�b�n�X�:3�������A�|@@���ħx����D�p$u��>&"�`?=�T ��ثɈ`0*��.@�(J�&�1A�����'��.���9�1�Y��Ps�:!gv5[� JC���9��]rhC������R�:�Gz��$�O�1����㞌��z�Í�՞`!'���!���ذD�'���B~bl���������V�-67��g�gmv�ڒi Ř~�Z�<�W�E^Pdѝ��"(n��舒F2.��B�R����|��Ӎ���� �oM�$�Seg���C������h�
C���d^����&he���ȥ�́A��K	P]�/��h������lD6gY���ĨӮƫeG�7�.�0ߵB?��M�V��lk=g�{V^q`�U^�[&��W߉J�='�(3:6��'�MCm�i���֭2�^�T)���U#�.��ȗ�֬>���[���d�D���Eo��5H֛z��n��x��ʬ�hsLx28nb�d��V���h���!`���z5l40K��Rn�V�������hC�{fw�1�{*��{�gGv(�[��ʠ��"{T���q���o�����w5�$�EK��/dz�	��/o+q�I�f�0M�����?j�|c�-��b����P���(��Ց�@q�ӫ`%7<S���_��U��3%����-���a7[Ő�g����~5���D�#=�F%���Y���!�4-f|�Mbs1:U��W3��n-���+�ڲ���]r���	�+�D��\����G&h�d���Ѡ�8J�l���g�n��?#9�]�z;�'���&��#r���y�X�oq����qѐ��պ=Ԃ������sR�����~@��O�����ړ�����u��E_��uH���a�2�{�BFv��J-=�Me%��p�f!��-�
���n�ģ���q��@Y�M��NՅ�f��&�¹m�$]��h���|�/��}��W�m���t��$��b�zs!9���!������^� �)(xV���+}�l�]��1����պ��T�Êo��Y�!p��Alڐ��Y��,3%���%�U�ǭ������l�f쬣N�nw)�����X�M�Rl�f�#8<����XAt�V���7bc�����k|b�l:��@���c�n�=�8�m�׈���4h�3���b:���.@D��E5�ѨV�,v떍Ќ��ksݖ�r����͜�*��H������8�~�=�����4N�Y1�Q�p'�M��SLl����݇�����Ȯ֣�Lm՚~$UoDo��TmTnt��o��H,(?ٺ���D��j#�h��Y�ǽ������>
�e��\�8��t�m�B|����3/���W��)��?��Tu�D��p8����V�a�K:���?�^?d`�Ŝ��AOL�.���Q�,��H�c�PԀ����"v; ���1���
�0p�Э|yX�E1�x�I�s��9��W9C�r��w@<���F�+��	�U
*��X��h�zx���mR��t���}�v�v1�R����/���ӻ��`�Ԕ\_�S\�Z��|kt�( L?H�!gV��57��2F���6�K���[�>m���3_���'O�����N���~}x8"��C���5��o�r�/^�Fx�C#Ot�-�Y�a���C�Kwl�_��Ӌ>��{q�+%M���üL��e}/a6BI�6j?}+������H����C���N+B���>?~��Mp9u�
���̰/T����Hs�V$򪹁�Mr���	�M�c~��u��{%0�N1TK����7o!Z����J���N̛gk'�x\�8qE����r��4r��X/D���"�
X	��ݍ#P�`� ��U�$~z�X����&��s���*i�2��~v��;��bPl/��xaqݰ5�V��]��<:bĬ���Ci��*���0�J�dcĩU�7��]�ݷŌ�X١���L�-\��W`CR�":��"�f�>��})z%1��֌e��ozKR˚.��xed/�S�$:ȰD����@�O7������ͪ�����2�~����ʉ/*܎��6��i�tɻiJ��U�V�~��"�-1)V�gQ	�h5����u&�`:v�,�~:K�}c�5גhx��0IY#��v8ݮ��|;8+O�#�\�Ke���j�{]�B���.�N��MZmT���=�j>�?�3��%*r�\8�������ܿQ1c�|�a���\܉ً޽�mg�l9|kL$��b�e �
�X��Ѡ�y��[�a����Ǒ*����m�u���bO�P�+?�%��O�9�\���e�N�9��!�{tG�F�He�bU�g�9{������;��+���H"�8�V��Tu�̒aQ	霴�5;CU/K����K���8�P��ۏ�)�M2�3�S[�Z;#����?�Q'&�������? �$�ʉ7�R(� #�G�::�W�=d<e�r�"�����q�/��D��)��Q�2u������p�-^�o��%=7�)y���́:���c����TN*��,����,���u�{�ܜ�����f�-ȠM�˻�4��|K��W�e��1%�kю�l�H̊"��i>�����t`�3N[�-5�?g�"Y�X
l�W� �\��_�#�j��קd�
3.?�M8ƃ�,fg�Jg��b%����J��<�Wkz�����s1��j��v�ۘ�zI�5���|O�`�*��� �����U���q�*B�6������V1�Nŷބ�cؓU��e�ㄽ��]+@)XN�ڴ(cwôgף��~_B�8�G,�؄���֤Dlm0ǜ CٗšƮ�����7���1�� �>�2#u��V�Y!}�%��T]���Hԛ3W᣽9��Ĺ��s�a����;�����`��z�W�q�3:]�2��,iX�2�]�G�|���d{Y�5Qm�b�O)ZX���!L���r��n�)��(�M���7�����;1_��ʢ �2(�'�8Drg��x��Vm���RȲR3a��v��ľ�2�'�6�31��g��EuV[����T�̠�-�jI5&ܑ>#j��xů���+�*�M��1�H�k��S�{z�!��͸Ί#��@⁜��Ot�*�)��S�"_4��ȠL���`Q�R�	M0g#b�`j�.0]�+��湰�"�8�M#doq}�w%f��s�
N�f�idB��~���W��@r��ċ1�5��ˆ�,�>p��q���pr���sUv�cz�C�H�kQ��S Ğ"p�Q��[�sT���	(' ��ݨ;�牀JQ��6dw�G+d���pZe�2�o��Z���|5M���i�r��=N&����/0�1��<��f �yF�6+��oIF��/J��Q�dAh}�YX�&��#랖�G�Y���m��nsF�ѡ��\�w��yG�s�f w����Vq�/�Ym+�����R����W��k�OO��N�m���o�[�<F$O�A����z|��vF��q�Ii��i�N�鑷=Ѝ�߫���^�b^���N��)H/�*�ά�U�۸�(2fr�ƭ�|n�D>ÞR�"���*�Uo��xR;\�*F���iKF��q�{���T	>U��O0ϙ���0��9=��� *�~.c����peW�׸�����p ��� #*T6^kQ��D��䕯��8�bsɞ��%�{���{�70m���2�~X�� *�8lB�:#��#��u�L�rb�^�a'�N�r�f*��pK����_��� -&ubɀ��0���支*�� a���%�x���D}��/![��щ��s� �}��$5I�U��tz�6#E�����<(f��~1��� �d�=�e0fn��#��[��I8Y�ܤ�C��+�h4Ɣ��n_F�P��)|k�0�:�T�&m#1oV��t���KGC�#݉��>�����i�L�.ӽ���L�����@��3�<j���ו H�f̜j��F�{�	�>57֡f���'.*�������4��?�[����U^@�vì䅩P�=B�ɆSR���_�](�%}�Q�y�K�M���̤����y��?�UL����	�[���&"|c��`��C�>m�RMN�5���!h����l16�����x��̳�b�4��� ����"嗅Ə�
�3v��O�J���K����7�XˊX�~_U�T7!��[� �D5F���2Nԅ�����v�x�J��v�hE֧"����4/ċ�S�l��Ր�FaF-d���l$�H���(r�R^L�=�Tޣ]�?��sƞk)Rn�}�Jϱi�K��!�\�� ���,���g����9�za��eI�ʋ��dR���ya
}��Oh��V�"fF��W��d�՟!�܋���>��<1A��cl��QޭO�4A X�S���giP�^���ʬ��*�푲�X��=u8�?	�GZ(+%'�mS�ؘ&�98�A�Ѐ�p�nL�ݺp�Y�߁\�	��%8g��u��pA{>b��v��cg�}�?�5�_���1�Bk�[Qs�{}�NC	<�?�W�����}˺�J�$az�H�W<w��[-A��j�y���M�(|�rn��S��N�ۍ�[�Rl2U� �����o"Q��g7E�.8>�3��>���\jO�9�~�+̜�n~ڡ� �������:<a׻���W���nܸ�� ��+6_�c,�)\�.wXԪ�k�\롻hP��?���D�=S/%��Aw��Vz�M�m*���'�Vb�b�����z��h8�%�\!�I����.3h�t{�	��6|QV('d�O�b�yE�8��eM;�@Pb?@����tWb�O|�
��l�>!٦�$�2�$C��*����8���K�H�,�1o !"tf|g���w��4��M�V��F9/9�[�����vۙx��4d�נ'^�k^C�)��. Y�xpu�{U����R	0L��I�d*�ð��h!h�zXI#�?z� .��l(���?��Y��Z۔��-�F��O ����\4����J�[I��y��8յ{F?��K'W^b.
�����آ:mؗ�SqF� �%[S�,q�DMo��.d������[.bV̳��h���ߺq��� K���.�ȑ���ӽ�AƐDbIJt�y�N���/u~�2���f��t,�����u	P]����1�tA���X�n�RB��'vs;!{Չ�n��<�d�o��􄮓�jRm'�O��ETvW�\����X��L�],P8��GjF)o8fwÎ�fB4m�v� 廓����Z[@��n>
d��r��)�JF�3��_���ϥTI�=pɷo�H�U ��a�;�[.왎}�-������A6�>��̐�����A�ѭe��@�??���A&�Q���]��M�GH��'�@�t��}�8�D`��%��i>�px��~�0��c7�H�m��y?���Am��8��}a�I�(09d��a�N@P�}���Iz(�>��4���d㈢��TFg=�uL
l���4��EW`'!��]�bN͕$"c(�e�Ow�0��4��_�\��X�\�t"q��с2�a�L�?�剬���A���iOL�ǈ���=�J�� f�0��T���cE������=J���rd�T�laV�۽vY�_},���7��I�5� ���Q:C&�J<�(�xS��%D�p.��&��K�șIÏY�^�<EEH&�p$�{pH��Zd�$�kx�
�F��Kfe��̉�R��0��P|6����%Ƽ0�d��,c�~3�=���@�&�Я��s`<-X�
���-'8_ͥr˽;���"� ���_�	�ߧ��'mj��1�"�e~N7.��G%q�ܾ|�G!|}Lӄ�S1�A]=W�Y懸�U��U{ͻ��3�RDy�;���.;S|��ݞ=���P�+>e9]�Όj�Ґ�O�����*n�Օ�M�9�v�S����CmӐ�|Z!FS߫�2@^�3��i�V{��d�Pj���(O�ڈ�ѝ_*xf��䪠��!�MY����-Qf�'���
s]�fkG&ڨ���^���LK�� X #(��ť�h] �O��5]Y����LȑZx�)�$֠Ʉ
"�}�~�8�xF��ȋu��*/G��>^˼��� d�\Pq`f��3�G�cqc��1%�4˭ð�2�i������KO��M�˖\'\l���2s"�I�b��`/�T�=iS���Fu��tEz}����l�smI��Owa���pٮB��89ͮ����8{��	��������Hyb�4�q������E�演����E����O��D���A�B�:t��%���.Q[h>YFbG7�0%�'Z)s=
d�kTMg�3Ҫ�.�����DZ�n���$�O:<�a �["�v��E��n$�-)����(�nV��6��!�_�"���lz(Z`��!�Ŭ@r\@J�(�
�օ$YPs� ��Ć��Bb4N�X������ܸ��\T��C��zQ���{�@�J*�E�����c����������vġ:����v�]�������#)����xb*����� �K0���b��ۺ��7�v������2�:�e�����u��XF��鰿����pb(��H� �
�x�7K��h}{�?}%"��h|悷��=˕,�T��}D�y���H3��d��3�R�#8ĄPw���E��R���l>G4Q5XmV���~�@�b%�d�p^�P���Ñ��k4�4 ���a@㡠NwᅕI��ԧ.�06���iNpn/�y^�.a��r�b8k~P�FM��>�JV�+>�������ޙUH$b�@��y�������<?
�]v�~1��Ք��T�$�^�ʈ|�3�ʶ{es.�C���C���6�R��:��p�]F�M��p���N�\&V7��N:�A�X�����#�;�Q]�wp��$L�� b@�e.w%�IO�7>vZO[�a�+�<�oE��C�����}9'�a���Jr���0u]Kv�cJ��ܪI���j��#��b+y2a��9���K�� ��K/�b����;���AY�\)|k�%��/�r��-�� �-���K���ަ�E��&�����VI���2&�}D��@K"�
c�Ę#�v^�z��mcle�A>5 �f�I䭋�)��-h��,��b���7�_��I���Jg��;�RŅ����xr���b����b]��eM��hF�tV�B�`6�@�T�SԹc���� 2� iNmH������m^����b���(���:4� ,���B����13+-���z��_���-ƿj�z%�7oG�Ȋ�#f	��FU}ӂ�<�/�:�wݏ (�5��+���㯱��J�!W�ot�<���-[��\c柇��X����d�;7�9�,��:
:��bPx�����1j=������J�wp���$7������0]�*j�hg��b��C/n��3�*�/G]�c���:Ɵ}�%�u�����9i�}*�6������i�,0�t�P	c���P�0��D��fgs�@����p�!2o�$g�wqD+� a�7VԔ��;��������󸷝��V�:��J� gIL���$`x䤩*J��j$<�E�g��a�rPaJJ1�u�7*�{Ȑ&�ru���|�̕�,2ů�]ܵ	���ώg3�7��_e?�%Q�#����i_��ok�!��P��r���v�z����A��$Ͱc�k�~7����8Ղ���*����uMLO���XW{$�?�����>���	�*��DpԔr�b~��[9b��g���ﾢ2S�-S}Φ��bP�����J��u��B}���e���9$0m3oĔ�y�`�P�|��<P)�_J�]�:����J���k?vg[���:<|`�upRI��P��8���zy���& \֧V���!��C(���C;��E����q�	�g ��o���<|�8�]� ���I̅M){}�79�f�t�Ds�zVFD$g�4�L���^�ۮCΘ	{��]K�xf=�RS��r���p��sy�`���ƹ��^=?�=�������rĉ=�v��w&hJ˙�����H+�.�SGP��M����Ŏ�P?6a�����d���U��)�}Fr�=�]���h@LE�)y
i0�^s�%�7�;��b<I��rV�8QP$p;#e:�r��ש��$�DD�(:���,��P"ؗ�F���+�f��qP#(����Z���ҲN���͵��(ź���y��e�M�xz�\�v�y�H~�xI��C
��Mp-�Q�=�cMsZt����w��?A͎rMx�GE�fC�łe���e�Y� ߅ ЀJ��z)�}Pvt�|�ؒ��{�}��/Vivc�C��l��K�Ң��n[��U ���/�;I-	�dj���@�(QE���σ�^��-G�rL���v`����iN&�5�d��n��V9#kt����)��(Q(�y��Q�gR��@�t�%�7v���J�:�1Jd|�hk�b������a⭯�c"<Nt�n|2_f@qaX�g\��^c��A/��L�%s�9�d���a�����eϾU�2��LnV4�q@�h��E��3a�69��J�2�Uns��m����c��$��G���=�S���yw�2'o4Yavb�(�G����H}/��ͨǕ�Dm��J�XJ��j�/�ۻ�w��
�������hS��5!���s�n"oh��
���N��8�fߩ�-D/�U�N�8�H3@�Hͤ2q�tne��ʩsrLsB������*������;.cV@�I��1!�c��7)z����\�ň�04&����	�}�o���m���÷T�گS���%�eAnMx��*j��O^�E�h��UF�:8z�%�oBs�X�<���aH�xsji�r�~E�����_���)F���-���w�n�O�ol����S�4n���Nt*�Ao3������_�~��T��k�����5�f�Ŋ^%|�}�ܻ�<w�r�|O�kX�i#��a ^�=�zm�Mp؇ =l3�������|��閍Ӓ��b�!�.�K2���&� )H��K��������hB"����z��-L��	Ϯ3=�����E�j�>]�-�ِ@��c���˂��gi���,3����Z	�� ��%�8-�k��}�x��C8����/7C�5]"�h~O��	��堗'�]��6�rj5��7��f3 ���W�΋��mrɢI��`ύ�a�+ʝ�@�~��Ǝ��_���+�/(������%��
���k[����2�o��\%�#bю�X� ��Z���J��Nv�����H��G�����#���=�&�&ל`�,L������WZ��o�R�	�E㲼���3�����uV�;�����i�b��#���~����������i�v�Er�Q4Y-o���iO2�I�+]�\0�����HDK*e�\��Š�%��ţE|\���r�� ,�:b��`�|KO!8^��П��a�%�&�^(|u/�j��8����t-b�<�p'�'zӢ_)�r��Q��p#�/��m�k�%��H�[Rau�w�_-,m%I��1����g�"XP=�mь�"D3*b3�q��o���x-j�R����Ό�6[�	��(��Xn����N�]��P�D�f@��!$�gC-`����VV����T磠Lf��+ql3�zHv�|�%V��vj $��Eմ�c���[L}S_�M�-|]+2,+a��O���;�qȑ����Q/�(�OΎ�z#����V6�缟�ۮH�SC�?�d�{R��lK�q���L��3�5Z���y}�p��G����XL\�w@+�<xW�ڴp:'��}��/��q�x6}>f�Q�vR�I.���Ez�U������tB�a��>Q�Ә<?�@�xk	gMi@|9M<:����،�uۻ�V;,�r
X`��i�����ʤ����Z�x/�W�s�T����K�°� �����X���0w�B��h�%p �,���Nq0����v���|Ub�Хo��q#ET�0^#� ��_G#M�"��2-S�9��Ƀ\��u}�Jnƕ_�yo1b�$_ȅH��dP&�g!m��/�ɑO�_��ed�I.������pS���1������/������?T��VWc�֩���*,�<Y��jK��͇D��VHs�G�r�zڎ����WIBH8bW� �8@9�FíTԕ�V�ŁLx�tT���J�O���¥5~��$�|�����2W���^�]%�����4���<���n�A�&1�- ���s$S
�R;�1�g���5�8/��l�|h�TŎnex'��� R�9S�<���N��M��ЈL��˟��V��$}�4�]�A�SD�6��$6*�^(�p�݁wC�cR��d�o*�o7�]j@_��{�O}tN�e>|m$/��WieF�ʜ���Z�Z��7c� J��c�Ij�!5�M�l!�p!��]��g���`�4Z�����a��ǰ����W�3���_$��v����j��$��w2,�*�'Mo�C(�ʵ�,A�P��|% ���;ԛ�ɨX�H�`M�G?殯���Y�yW���sqim��D�57�Ta
%xV�������.��C�����4a�6P^631sq�a觔n��7��%�bU�6���O��d����9K�S*k���P�u#Ԋ\,�A2`�(H�H�ꬻ~�W|�����܏�qnZ<��x8zv����I��}�� ɟ훴�S�׋:�<ELA2���OJs$�UB�N�U�P�q�0�)�}�`ס�!��hQ�^l���?E�ߖ/����:Y��a�������֝9�xBJ�_��nV"n���E�(|��m@"����o��4~# ������b1T�����2ꑅ�`�O�Yn��7�f��ﴄJ*ag�����o�!�i�`Ŕb�����]�,���4�£�/~���1/���B	LUc�7��1��n[�0Q^��b��!C�f��k�qWaÊ\��Ƶ͋�������,�ϓ�G�OSH�9�7�2�����k��?r*6�J��b�R��<X��NX3�Y�om�fC%[T������r��7�׎��ۭ'OT>�j%��2r@*rl�� ��7l2���^���P��r�s���w����WJ�$L M *� 
������{��x*n�ٲOЊ�v�NR��}�ԧ��h���}��ys�ǎ�p��s��k��0�q1��4��)���V��$[�Ɯ>6&�ib y�����bn��
k��Q'Sם_H�Οx�J_�T�i��֭�j�ύ�F�[��A=A�|���(&�i[�V{�Jm3�����,�!�Q��W�L_N����������:6&zU(�8stx�^b{��&*ӱ�J]Ȑ����ꑷ�F)�Ύ�] V���x$vr��O��c�8Fu�P	���)(�6Yl� ��"���t$�nM@���0.!�!)�^�}���r�^�]�bG����s�|�a�U"e]Q�� JŃ®��z�W�����+%��Da�W����ts^����Njē���H�V �M�T���\����Ɂ~$���(���Ʒx����{17lKܻ(��&��Y"X�_�>�/g7�J�R�N����N�gJ��	�م�K�$���� P}���sA(u�Hӧ�c��������xO~M�w;9�0eu���X��B�n��%V�i�#b���)~���&��@�̝�6��B���'�h�;�XOE��a1�}�sf�	'm��-%_����	�����c�M,�ٵ�F���j�D�o3�{�Fˌ.h�F>�O���xDM�]/x@�<	Q���imH�����}����3IG:��'ݩUy��RNJ�C���@��;\�߾�m����!�g���ןy�T!N�@��23پM���z�`9⡶0���U����E��-�E	�5j��}�� �>�"�!�^n����*�lJ��X�������=��^���L�����F����GZ�2��X�  3�Dr��K�kj�{#=t��G����<+b��
��F5B��d�&�E]��N�!#jW񀽀�&�.N��U߼��ܗ�fL��#?u�	.�kn�ﮟ|!�_�q���J��
엎�U�c"�|H�~7� I��ۓ�����(w��[� q^�+ul���#_�a���5jf�Q��Wm�2娪�'k`K��!~
��{��	��;ʱ��54�&������X�\]�՗�%�M�A�7a���C�*�S|����� H�Ï�4��ik� ��NM�'�,ա�1R�Q�p�ԢoEd��׈@8���Q�T�ެQ���W��zx>�'�'U�O�zf�  0�:�Cѹ�UvW�ݑ��;Q��P!���Dd��܍��B����n��Y0�{�do�����r��)��=������2L9�{�01X�u7��|���𵣆�3�K/�ڭ��������#.ݱ)I�#Z7�|�~,� �>R<YpK��V�G"j���!�ˆ`�1�눁�
!߽ Ղ���4��؜S�畛�ֳ�2�^sKC5�'�����)+��{pH�~���;��J�צ�
���݂/+����;w�IE |Z_�+�Ԝ��|�u[l�gBmXt�����6�co���q��\P����E�=�Rq[�)}*�9Ӄt�a�b�Ϲ��H��}5��,�uy�*� �E�S�nӖT��H��Z��� e0T�>X�	�I�Z�QQ�0�p�k��nt��Q�Ű���gHaoK�i�F%��zh�oWXT:��2~�����t�[����BxN�� ���/x�������`s"��?�r��
��W��~ɏ�4�ݴ�c	���)'�a�6�x5E����8��a�t{	�����st${�-���!7����	m?K�*V3�:���+v�i��@�7����]�D��ù����n��{�cPk��"dJ"_}�cvՔ?����ݧW���s�K�$�^(o���#\%CH�$����/�2���9(�
��9��(S�zɈE�Mݪ�������#	z�/���6�2�^�:�.��x�� )�sM�mK]̿	ݖ�9��
3U\ԲJ���=��}X6���{-쟼��>ר^�1w�z�� Р��t��r�M���еo�=�����N.���R+GJ�Z�>C"Y�:d𤻟cv췌�������U�2����9Λ�G��5�8���N�5��_-�5m�^K=Q�W=zl�ts�c����i�͜1�Ƌho*�y��=	8���o����!��BK+���_��E�(�Mz� �o�F�	w+`O#טژ�<�2�[�� 1{�l��1�H��Bd��������F�RH)��·��s6�q�y�I���
�һ[�}� =�"�F^@
��ەD7I�<f�9��g[2��a����x��W�VC=�����n��ry!��s�V���Z��<���CU^0�dyf6z�9��*W��d�(ɯ������|�[e������}!����`�$EL�a��!'O��y�=C������Gg��vk}�k�4{�a<{}�=��	]�����$��C��g��k�RN�R��T��2�������Z��~��ЀSXh23�$�|���%e{�����#)0��Uf�9�^л��l�Д��� �O�{�O�� PB��*և�p /xc�K��*j��}�!ƞ��Yӧ LedO��-x.�v�����tg��>NC6�q�Y-�t���':�9i� Pɐ K�O<�|3����5w�͓�N���(��\������%����y�_���{��o�,L��PcL��q���\U ����ɒ_��=v��i��֣v��EN�2�,�r��BA�vY�hpB�BV
��V [N~��x��qx�Qӗ�5��-S�:G�dZ�����N�Q��i����Ԭ��"�����$���%6��s��G4����B��o 8�Ne�TQ��'�������G�)FZs[5�'&0θ��w\�)��SG��jpL�D���&�$�XNtP�׃�]��z����w��~$L]��?Y��P?��xu�U<�{�R�wF�v�� ��+T�S�Ws�K��.�\Y�0gL3<%��K��Sh��4�=o�e��(��"�kt�g��Z��� g/5���j�U�*|�p�҂�ó���gJY_�8�����{-pH�Ru���x�}�0ʩԮ�^G�G�a��=O
!���R�lr��R��s-� �5+��
2nV��	�Ľ�>y��޳G)��=1ԖQ"(Yt��ٖ��u��}{s�k���:{��#ޢ��İ�s}�+&�h�}bd*�I7�XvEhkMb�|�}�8lkiq"Ah�p���X�qYg�Vӕ����s2��W���!�a@���Lc��ȡT�CGH��j��ŝnR�b� .�ϩ������)��YP���d/,�\��E�}�������_L���3#�rTC��SY]���[�'��.�S�_,ȥ�L��p����W`��J�y�i��A��W�i'RA��ؽ�d-gn���AE�$<|��������o���=$���Ͻ��ZO�hY*�����D���e#���.��������{{�ے٪i�V����
���ߜ%���
��..K�qp����i�5������R	��saA%]Ί���$Ʌމ��pn�=B���-�����L`Ϛ�
D����V}�������I���e��u�C
u�z��SL�o�Cc�|;-U~�,��5,_`L��%�r	�dn�����o�Kxṯ�Ν@��.�K]h��Ēj@O�J�w�m����Ku�oB�U�K�Nb�|=f2��(d3E���+�]�kn�����Cr�qP��r�x��CBQ�Ȫ�(����nP�+Z�3
*׻�4��e�������wc����{+7�'��H[)�8��_F�N.�߼J�[-�M���G`GO';�0�duqM�gHEEw'$a4�}��f����j9�4��ofƦ���1�'*r#�\��Q%�,a��F<}��u�TT��vl��q�-�M`#tI`ףgF��m����<��%�"$[�P�%��{QQ�Yq����~-�[���}$G�	����:#zX������'�7��/�������F=�
���4�����;c�߫����ސkWvz^��,��6�Q�Ā��|6�����slc����@���{����
V@�,�d�mg�Vc�����Ֆ�bO>�'�s�H�{�\�ߐ���s6����ĺ�H��x����(ÐBoE��)���A�1d`{C�
�B�$���ϥ��w �����d����64K�N�{/Ѣ9_�����Z�9��fb��n���@
xҠ)�|������� %T�oW`�l�f��;8�;�*�(�H���-.�����{�O����>���snɅ@����^��P4�+v���9bq�Q�������Ai�}>�є&|z݃s3��ԉ�nw�4%r��c��{oᧂ���/Q-)PqF�1���O�~��M�=�������Y���͌����C�-���Q-��sV�2�3�3�����^kd0(�H����;���Y�x������@�Oֱl�N���/�V���9\(���ˡ�f8�}5��o�b^�f|jI��+�D���Y�
·�Pdc.��u�~9;^t��eQ<n��c;H�ϗ:P�9Z�k@w�)v��.jR+(p����d$ ���Qj��x�O��F-5�GHF*�j�+IIŁ-u�%����3������=o�C�iz[d?��Q(��jӴ�%���n���ΒLS�d���F���ü�O�F�uG[��/�az'v�o'C��6�%S)^!`��]@ڈ0;�)�F���_�_u;�i䰄h�[�Z�^ŸW$P��4����Gg���������W��������%��W�V*?y�l"�v*L���SȐ`<q]��(��r#�����jc�D�ŧ%����SN
�������W��B�E.�/)�m����e�g{hIq�\��'��F��,�(y�����{�ˇY�a��,��$��"�>�� �)�򞺍`�f�-����,ly�BJZlz�#'���V[)�Z���\�Q���D鶂O���@�>�bOw#xCpA���?�2�A̡�[�n��Ϟ�H�s�H��
fG�*H"�-������-�_x��w�a�=N�=��������-�c�/�ʣ���I+�Li�X�i"���t�B��0R�uFV���7�DC�X�_�n{%k�}�n�MƇ�8Jvڀ�8l$��
��u�U�mE�M��5�ٿ%�ul1i�+E�Ǥ�<T���̂��>�Ҡ�����FQ���ԕ����͇�p�&�Y�=���j�V�YIm��Kg�j;���'�34⠚1	f-���9�+���ӷ�f�H�#�
y�e,�q��d�&\۫��Kdy��)�����6i�Ѡ2����U���M�1���$��n+��sY�t@��9�	F%ã|QR`�T��S{��A��Ԯn������1��}��>=Ƞ��1aiN�S�g\߀��iJ�.�k�P $ůKٖw��`�
�i�|S<taR>wZ�J��Iy[A�P��˒0�����T�OǙ�͖yБ�N3uk7��T�� |��=�Xu�Lȩ\0�J����b�2HP<A'�qդ�/��\��k�tOe/����R�m�*���=hP7�+��͡@)��y{�F�y��?�ͯ�!v8�{���{��[�5���t�%��������闃b��y����=:�|$[ �Y���k5[[Bu�!"a>]��j/�����$�NZ�'hH�]���yE�y��������z驧5����L��6��:|�0�9���YJ�$��~���	�:�M0�dg'5���v`�˘���S�=lf�b=���N򔀂,g�l�M���ƺ�QY�/}Ó� �L��t�cH/'�Wu���DX��[�A�x�4��N%���ǻ��.�`0��l�K88�Ί��u���.�G�kX��>��PV<���Ը��� z)�{i�>�?��G����j������h�j'IB������/�j��(�~��K\q���<�A����@������Co���z!5tV\*3�[!l�\bn� "��bZLè�s�����Vw�����sm2Y��F���o`�a�H�P�рڄ�N�y|�H�}M�'���̦Jۅ��I��S��L��8"A/���Z�2��gkfQoq��\~��[XDY�W�8Y�%��u]�Z)$���wǿ�*܈Ubf�k"n]n�#;b�bC�~��@Ց���Z�&���[�����x��ƺ�Z�+27��!���v�_���;��2֤�z��|lc!6Dp܍Ph7��M50[�S���	���"z��ו A��T�e`4R��<7JA��� ��Xr�\LQ������|J��Ȳ�����p��u����M3��#9G~q1�>���+�V��K��zղn�P���Y�i�(Ow�Y|2��jq&,��X��w(x�2n��45�ޖ���:��;����2�	ӣ���μ�2y!��ֳ�jv������
,�B�֪D��ɴ�b.w�<�pI�ȯ\��i=�6�h\d\�鿂�3��}(�p[@�v�h�WX4���ql���^��<ha��.l����1�P��)�Ε�\��$ ,F��9�����R��SY����_m�lx64���k��	Wz]�M�,[Z�,L�7�$O4m7��1[^]X�7��A�r V/����I�|���PbO>������K��t1�W�ޫj�ZoY\u=�+LeX�7Jެ�h=Y�����1���̘&��6N��v2�^��?�p���!�_X�zI�r��/�����s�6���pF���1A�ץ�L9%<̙�p-��ޣ[�L����)���r�F�������� ڑ�Q�C�w}z�z1�A�ju@fY��6�N�{��IT6��ֈ��O�Ӌw�������8^M�d5�g�`�����k�)Sa�0��g>��*�j�.ԣன��`�X��-�d^����~�1`HE�Y��Q�
2W�)!�|0캎�*w'#U��Fa���s��vq���
c�����9s��K{��86�9O��\(��z����W�Rf�>}fN�*��P���{�<i(�>��e�[|��<f1�#-�;��E)+�:W�G��$���5�V|��+��q:�]��`�BZ�7��S&q)��N�3!�˕4%�Y��uÜjX�*۷T�q�Rv̳�Lb�_L�{��F�M[��y���x�Z��QV(Zyʞ��י��csF�;�n��Um@N@^��3qݚc�Ƭ�L�g4��~���#B]>k���d[��x&c;��4a�Of�b��"�n�ah�.��@2�H7���x�$QЇ��A�B�Sm)�aʟ�s��Dz���1I9������jևK�t���]�RY��
��<<�Zkل����Aa���cՂlƩ��M�:}ͥ���R�s8���/����|ou�7���%��.-��}kTW_��v��q����`��6�m�Sl�P{\s�O���w�b�i4�9���(qM�u��c5 ?)�*����nUi,D}Q{Ef��=r�o���HH�{�1�Nn�v�$M'�(R�q�z� :J��`u�H5�mD�=Hl�㎝ᘢ�~��o��������`p_���\�73�F�SNt$�j����T\�����aQ�����}I�VA�Dy���&a֘�~�n���2e��"-�
��+���vB&�<���pK7�������@%|�J��A"�y��ҵ5*%G�|�������r����+�����ڴ�ǅ�A����eq���R���2!�k�rGL�Xt�]F�T���恓�r��_�1R�E��Q���e��{ly��b�]�.*��ـ �����_9��gr�R�JE��vw�m�b�2Ǥ8;��{|I��@�x�Q�E5Y5���?�u����V��U�=���68ܚxge�E�y=?5�vraM@z�W�u�p9[Iv�TU?�^/	ӭ2�.�����5=B��+`7�/1@~Lٴ��w ��׌msT��1�kS��֛�����qW0��,���67l�b��ݞ��{x�Y=�d��s�˧�SZ#xb��D�"��X��c�2�]2����e�3hV`��^����4%%A��6���	�el/\8���zbl+mN��R*�Ɯi�=[ͪ�,Z��v�cn��GLʿ��L�!�m�Cf9��&�,���-E�zkW^t��Vg۳(��Q0�j�����n�cf��i��z	���o���O�S���Ä�^v_!�^kg�c�P�c���>��h�2��(�5�uGK�p��I�'>eP�[��C{/J� e�h+]7�!BTKy�i�:�\�$��M"�5����Ip�y>"!,�i�T�v�d���EC��OoNs�z�"�o6�B>�7�y��eac�����xl�l$�1���ٵ1ۖ��*8�B�T�2��	��A��)��k�O+V�x�v��}��,H�5�f����^�
29]|t7o(Ke�!�%\@��2AXqpE����l��:Ry�W}W��hz�������?�'��q�q��^��藨hm�pn۽�ܠm�V�,�%�6@��j�D3x�������-ԲR�a��J�T)�A���3>ZC�s�c���f�^�/0���=��ʃ��yp�X�[�$�f�J"sw
��[���Za��e"ҵ��E`ԣ?�K��2	����A���Q�����G-�u%�
� 	�8��	U�-+6w�Y'*F�%�w[Č�^��yΚs)mS���"�\�����qMVB�Z9�f�%�e��an��'�\�*�;���0�r�rա���2�!�_�}9z�߅���l>Ȝ*$��"���W�Y@?�Êx3�w���%?d�~Q��!0�4��9�v���6���޵�(��������N#^583,�[
���u�o�ŝn�kK�3�A��k���H3V�t�"��K�2�X��e�p��4�TF����d�h�-��{��g�#j�X	�Ɲ"���2�K��ioU�C������=h�*D8�ԭ$�i�+NH*���"�_�h8´5z�����m�1��Z22����N�p< d�����Mr7��Ew��<�[�)����%Q�x5`��6��K\l(lJ�sj���(e��i����&$����?lҞ����b�;�|���&�8+�kd}��Qw�G�W@ߋ���rz�S+*s7M�8w���S�߸���Zuq��M�׌�[l��]��!Vv�V\���&��7�w�B�@ʬ�`c��>���8��S�d�����S	}�%0�ݦ�Ghp5p��ٿ�^T"Һ�!��,W��U�Į�Z��x\��b�F��5*J��`��t�|�<ؘ������nJ'���,��2Tq`�+I(p�Ͳ��}����0u!�������Q���-iO���צv�	�ꉬ��c�,3�$Qb��5��� G��?����/�T��xr���>1�3q���D2^���G�����Y��4����[+Rt��L�bʫ�g!��7���RZ/J%�� ��5�#�}D��V��{��+ ��c�<�4s~�0�:Bg��h�W��Z�أ ✀���E�����I��`���M^�LԖa�#.����!�e�/@..y�B��e�%o�tٳ#���3���࿑��=��h�]��D�h6�
-!�"[���������~�B����,���~�J����J~���Rȋa�]�TQB������B���W@9	��~#.y���`�������,yڧf[�ى���DA��:5.�!����a32�+���vzWtc`h��L���g��!r���k�iB�>|�]�����;�� ��Y1c1=��B���֥�81�[��4(29&Nj����mWi�̈g�j��6.�=l��z����ʍ���rV�\GC[���/�G����I{����H�2�s��ޒ8e�bՈ�P	�z�9c[4'��4u�r��6\!�����U)[Y��5���xUu8�Xk R%���k�k��}�_��)��O�&��~��@�^�xa�C�E��B"7p]W%Б;p����o�$7	o�̞�"81P�¯�Kv/f���[i3��uBk�F�!�
���ɲ�v�� ���_�^@>a�ٱJo����ڗ���:��%�3PgdC�.����S�T���T�q
=������M�����~�llj'm�w���a)�u/����+��{�#�������
}��;Fr2l�LR�y�>��x��/��2"�#'��G�M~�'�$px_�y�A����Ӊ h@������k�.���&���� F66-�&����>��=��s��Xw����^F���/-��һ��pӖ�qqP��f����޾r�'!�v}hM[����y�z���XiN�M�8��0��'O�r���|���"���%��gj�����e4lͅ��hy�R����X~|������[a+�όG��7\���B�/w.:�s�k��]9xs&X@��=6������@����A�^������+�E��)��r�AV��}�W���A�>,�p+��z���D_M`�o [���5��._ݜ�l����2;���~���Z�kX�5F@�9�3��)��:�:Q�/ox71g(Y�Ijuν��X�- ��{ _��4���&Y*��ɕ�i�Jѱ*)��uB�گ���ӵcYs����Z��a#�gHx[ZS�:#N��/H�g�Y�{꧰���%�8��g�0m�̷e@dOP�.u,S��o0�y)}�z"MLRH�xO�H�z�(ͥ��ؙ�}!'�Q>���;�4i������*��9�� ���ΐyK䦹��_�LH��1����_��
�\��K�����:�:(\q�D�\!U�șك-Z�"Ҡ��y�-+�(���Ay쩶r|�Y��uQzG��L��!͏�g^�%��`�p �y�x.��6_��9O��N�A�X��+N���&B�'�U�Wm�m<���t��}o]�Re5�OC:T�V9���jv-�ٳƈ'K�Q��y?�	 vae�#�O��g��W�U9�Đ�f�{�,I�W�q�GR(y�(�q�5�"/�~�ɐA�Ӈ�u篻�fw� Y����GI���`�Rޔ�W���k��Å���5X��H�J��F����)0��Z9a#�%ZqҐ���5����j�����c�����g��ZT�P���x\�ԈF���DF����= �sZ���d�&&�/v[��iq�F�o��=V�� ��}�tJ�վiۛ5�I?�}d!H�$9��lw�(�y���0����Ef1�<p{t���+�p·��H|��r�H|��S���,.v��:j:^��X������j�+zнa��<�`lb��-�+��{Kf��(ULm�����!$�5mk�8��`�!�ͺo�%O�%��67�(^��@Rs��E�H����cp�S����o�}5h�f</*'Z�B H�s��G�.�����j�6�*�+y��{����	�C}Z�i�9�t�T7�i�D}�5�S�E���r_��/���#�c�ql��n�U�m1����w&�3:oC��C��8,��e�va��YFg��!Ͽ�~ē��yWK���EO����'��۫)�U�b8��L�p�W�KG:��3�`����-x�\���~�y�U�S__��Tk�M��9H��X�"PS���}�3K�z���P�.Z��RK�In�w^\^�v��Bʑ>�C�#T���"��g0{]���Z�5Nʳ��4���P)�ܨp�Pk.i���c_ �[�Y�
϶
�#�KM�S�b��I��7�Gy��dT.݈ �5�B�(�!�&^!y}��Zn������	�7*�E��I�gb�P]?V	�MDq����+	.�����qK�g�V�n>���!���a:Û��	{+������֑0g���Lʗ <w��o��2��5�i{̪I"�[��Q~�2P�b�=v�$oD��sj�� Z�qEC�f�
ה�R9o�S1�dĔ�*6�CN��JJR���,�w�N��:%S��IL4Y�`��Ҹ���l�C���t�ě�(�v��l��ڌ�+x��qfh^�5���9��������ui�p�m�۫d�?UI�#�������4{��^�٠�>rw9��~٪����r�o�M�P	�s�1��U��`�ݏ3=��&��Ys�γ��u�U�Ia����8à�l���H��	�4{��ܯC���V���m��I-c$jGaWئiw8���������:an�}?��a�N�q�ub�:�5N�3zE�^�ʪ�
	C��b�;[�X`��tc8M�o�Τ'ih�%�z!�x�;E.Ȍ� XV��Ǐ�2J�Re
6v&��ܭe��(#&����Ԧ� ��u��mƶ��36�8p�d�Q;�F�d�ńs߇I��n������H��UD���&b�]��΅�{Tg����=[�=-y�f�#�R#�RR�g�s)'��Kx^��F���0A��V�	ݙ�J��N��n�L#���QR��/0�.�BC �����r'�X��9��52#�X�'؎!�k��:oa�$��?���u~[�Ai�vro���!,��y��y���A�T�rj�O�V���ݔ�PL� �5��T��r��zn�_�/oQ�[�������w
&��.�2	�|{a��.Ϋ���z÷D L��fz���
�uo@`Zh�x5g�K��a*�+��C��䮷�t�����@	0cA�U5�7���W��uf�
-J��2}J/�P*qm51n��|������I�2���e\��&�#��q��/�Ϊ�V���tncM'���G�n gˬ����BF0/����k޴wK$,@��/��:��߫C��*t�&�O�d_:k�R���v�H�>.;Ղ�iXh��Qn��9��B�S��y�!��QA�Q|��ru������QU�;�A���f�������B*vb6P�:�����x����Δ�*����K��5�M��E��S0�R��������Sk�����ٮ�
&�@�9�(g�M�z�k.~jb�:��q�	�?�Y@�BV�C}n�	:V2�2�D�5�A�8����H��v��z���L�H��*R"퀞8G��`S�����*�!������G�^�#3܊����Z�;MM���2��0L�<ےW��A������Q��&�m��.�����L��B�V1�#�x���ǻ�%F�YI5N���lpveXss�]��{��6JDZ|o>hw��=6oU�l�2*��XeO�5��X��4�FiL~���ߖ�
%)�/'tn;�@���m�~R�L!���4IY;㛢;�؍!�J�k|D�H㳔m'���zG�"$O ���&f��Ҽ~x�����ӏs�����Wj&Ŀ�L_L� ��TkQ���0�wp�V��7�S��C�4�-<G�6����|a91n��7ɖe�ߠ]����g�����x�� r'�Li<���
��? �	�3�a���#=E�� �6�N���)��4e`,���� Y��0����,0M9hΕϘ1"��m�hD����-;�c�#�HV�[�;���f�����|c�,'X�h���l�HI�d3'�C���Y�z�'P�Z}'O�;-4�Rژc�K�p�L/NW)�'��+YCr���������.����cf�uK����۲3�z�(8Uۙ|0%���P-�3UF����4���d	�+���ǎ7��VZ�nj4���.�b�~aa���"ԋޕgjc�^���p���6/;�4����|��v�Yc&g�x���2|�#~َ}�ʗ���̯��'��w����}-;����ػ6O͔��Se�����)����6_D'�^������z�N!�aS̍?�R�>���<S~���9
cھՏ��������b�;=F|O�L�T�wQ\S�J
L��$ެ��ɧMe�R!�S��kmRP�x��K �$�^<r�8?����Ј|���*׭JM��"R�a@Mo���ʀ?)� G�n�����)�q8����g�������ë��ܮDe�_����7��Q�C pjB�T�"�ѥFC��Ů�q�$^1��t/N�pp����������-\�#a�#�C�S��_I�,�H����c���i��;�]]c����c;�meJ��ɖk5��%\���P�;(��K"�T.ӏ�QF/�����@2%���7���
���{Rx~�p�

B�FuSv+[�O�핍�!ZO�jugv�{V�_w7�bc�r�r� ����6�O(b]h4��𡥀�Gzi)�[	���H`?�#<