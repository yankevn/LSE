��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2X~�*���O���k�<Ζ�?
J��I���iR��eϴ�J�Ij�Je�V�e��JB^ �9�E�|�h,����� �������c���k�zbr���A�5b���J�f�"UP��"� ^$wW�1�t�Ў��	�/G>�ڇ�[mȺ��j���K�_���)ϕ��4�����k-�mVs/��͆Cw�$U؇�/4dY���J�=������ ��e[M����
㌞c��|?vNqs	U�{)�i��D五��*�|!���,:��q�A-*��aW����w�	N�5%�5�2{�.7P�K�s?�dэ��t���x<Ӹ1J�H��=�Q��Ud��k�I�k�j�C�v�ԉg��u���ѵpq�U|���̳]�ޚ���j# 

U�;%��St��-a��&-�%�c��m\"x���.�ON�ް�X�,��* ��?v �.S-�����=��=	�c�/c:��4L;�IZ�/۪ӨB�w�xei���J+|�_	�2�m��NqB޷K��ѯT���\0�w�3�3G�a�1��0��m��jѱ��ͽ��j=w��gR��*Ӯ>-vP����ͩ�RQ�i�W ���%#����&_�r���6bm�b�_:�}1.�r_U6���<�fZO$�}v$�je@�<�Ho�t���G����� ���3:K2H�y'&�г�pL�̎��D����u`7k�O��(���S��ӽdU��yTֻr���H�ҥ���aFu��ZWK��}n,��o��UZKH�,� G��(4��i,}�f�x|���%hHa�X�Th�;9�a�<����f��My�c�c�C�{#��9�9ô������8+S��I	�aҼ���u�Bf�v"r�PD��z�M+>�XU+�iP�J�<0W!�C�ǋ���e,G�.�<�E�6�ث~�>�H9>�F����*
�_%�Z�>�I?�f���{��sPk����.v����؜�a���7H`�R*�LɏM������<{���&�ڼ��%0\[㻔�C��~ȷ�˝�S�W�� �Fþ��"���)5�垡�
���Kl��lgl�{-����,E3�0q�zZ_�9՟X�ē~���%J����!T�셑X������R��uQI�s6�����q�Vy�O�K��3�@	Z��V���#\M}�v)�7�ZO$l��6=ҙ�&��)�aR���Ji4��r˖gIn��G�t���Xj�.Τ�&���m���ʋ����_�x5���ؤ����l/"�j�(�Mk�.!=d���z���(��m֓�B�5���Ð^� ��S���J�[Hi�3�$Q�RI�=�)���66��9����wV�m'�pTH�g�;�F��@V;�1��M8{m�S���PO}�,��+m&�/��})w��6�y+ȅ],��MMw(��X�D�lxO�����8^}�ㇰu0�.\��O��"p���Eɣ���e!�.B=3�����㴶i�;%�o�[SA�d�n�ʨ�F�8@t�0y-А��z��6�N���tO���)��c��0�ou��gÚ'���r�QN�&��$���>U�\�O��8&+��o�j"�ʁe�t�ҩԼ��oCH�G���p.���w١dHC�(��-��q �Ҁ���ȌA��I�o�2�D	� a��u4��=����g�{(����9$�7��<��#db��A�Qz� T_�����A��8�;�I����SdeV��g��癊����t��6:�(�z�c�ؤ5�Un"e�R`�}\?2��wM���M���*yw���[�� L'�z��Z�U߲L�8�ᜩ�`����"gl���s7��7+'�>'��3�J��a���o��!�w("ߛ�h�0�;9*/��U�� �A\�~a�.���$`d���5�N�y����?փ�F���'��j�#�"!��Pu+6�`G�F0��(���o���6	�*f����PKu��<$[��b�b
�j,���ϼۭ^��Z�0�Y�
A>�~���ǖ�ȫ���1f,�.��؍(���ƾ�fCzə�t@�"��WpM�,@)�"�i�騪�;�-u/��~�"��������څ�@צ�	M��S�Y��riZrE�Y�J�w9S�J�	#�F��kG��0u&����㆓�d�Sg1x	 `
���1VDxj�����x�p/��h�9ճ�̊�ge/�,p��;���w�X���0f�_���^P��g��g\��^��S���5Q�$�h%��!�ʵ��jƀ�F٫s���jS z	�%P��J�8�gWN�(-v�`>"p�ۣ��b�:��3���dZ�}=��w��V�@^ /F�t$�O��Mw߄��'�h$H���apϜ'eFN��~H� �j!�A�y�q�n˹v�Ӆ�0`Hh����$�K}@���=��1�9��|���/�Ц���'�%�ZgT&to�̄�>^�`����q������i78^7����΅�pP�w��3�^�-w�.�$�'t�n��q���nj�BL~�0S� ��{����5%&�~�^x.Q�X9X�V���H��#���ʸ��^o�9�E���(�qdT�$��OUzۈ9V�`�H��v��{�=̳�+^�BI�-j�eVn��E�������A��Ng�����#Y�yﯪ��ރ�1] k0 h
	��(����[Z;��zÀo�u�E:�?��|<������{�$m������Gv�r�0����8�?�+��RWG����&W
��~�v�j|T5�0uh6fڍ��K�Q��?����)!��W�ט/���ޖ�^��O����^�Hc3��m6&�Uw��g��d�{���
a�9
i���k�	K+Z���_����.h�܃bt���)�]�[��l��"A�c�\UR�z �H�Y�5[Ǘa�ۛ�@�Q�\a\_������-H߹qU���.[��F�h�N,=��G��~��[�(�Yf�p��z�z��%�Icd�Ҏ�[�
(B؂�v�d1�9E�m m�����w�L���n�3�V'���]^�s�Y$�_��c)�\�.w��j���s�ṷ�$Gk����C���(�H;6���W\)<�����:oE�[�׶za�:��Qu����^�y����(�T=¡���Z\��,��T>���t�L��D����ߵ/X>$�_�R�l��d�_�a�� qG'�:����0���z����m��m,̩��'%̤:�M�&c�nE~wߤ�	X�z���N���l�AO�a8S�"����L����Ϝm��+_N���dA�6��˻��%m����za�uL���YIӟ�^n��������b?E<8|���$J��b��Xn��1�&�H��¢����w*�Ԡ����NS[l��i����F��H����%xS�qۥr}�+�����"Cp��H��t��[R��Q�lQɘ$��oŬ�i��\�4&���!���yn�l�x�{�"�.qb�kw
��U�$��=��E�{�I�+�13�Q)�,\��y#q4#m���N�~���>�V�(N��젏���K�k&�G(7�M!�b�;Ie��PS�Φ��+L�r�T\��fA�>ɵ���v�̆�)����#�#L�
�T������8850��8<Hm�o�����gy<�{��oU�?�l�m7�|���������感Şt����x_ʥ(TQ%V�|��3�f��'�J��m$Ο����-���)��)�m��$[?��6N�T�Է���P%}�Z�ǬJA\���b�ye%�SǊ���q��Sɢ�<f^-�&��G�y���'�Jt�s]��*�M*M�F,�����!�L�16�[���Q)������C!(EH��ښ�R�M�����'�9��2l ͢]�pd�S�x1j���ٗ�b�E��?o����{d�<�=<z�ڣ�Dlro��#�n\���3{[;�ly^�u:�&�sl�W>�I|�T�
:�W���͟����`�͋p](hO�%>{D崼���K�A��������g��$�3G���D�o�KI�M�ЫCH@��
��ݳ���d��	٤v<����ѹ�+ߦ�����0�p�܆Nz��Ǡ�p:X]�Ո�x?L!�$t�T��u�}Bצ��-g���(
��J	�":uR(��K;O�T kg�O�hɲ���,��!��5a%)3/Di�.^M�u�v>��K���+0�]~ [�V��}�n�#��V��ɾX�G*��dQ��ݷM��џG��+��&��ي7��0����*��ɐu�0b��
�-�ۑm��p�`%#�`�5���tږ�+Q��4F��,-�[R.%:;[��߾���sq�o�ݝ�!"�� �rnXK���7uZ��f��%�5��Qj.Q��M����]��g4�U���b�>>���@q/�����CC�G�~�w��"k�������̨�>��t5|O�V�O��|�p'g��W�Ku��c��U�@_����ܔ��˘0���z���I2���V�Х��u�h��Ǔa�!�F��|֞Yvg��7̺�ȓ�FK�h\Y+�Fql�q)U�c��*
.)C)lP����N�{I��5����M����vf��#�##߳<U����Ho}@9�ⶵ�6�B��+E`��3K\$����������c�j���h������/�C��@D>
>ڜp�!�`������s(�?B]���`��VV"Y��/[��-YE�Ϛ荜����/��$�y�����Ƈ���G�Ɛ��}W�~�jE9�|�͖�.p��O-�@�1����f�?��yLI'���]3��0�T��o��^������R���#=ς���:��)�X�7�7� �?}�����U#6b"���n5]��M���~��1�si$+e/�ɴ����Ǹ�F��<!�3y�P�W�%+��)�����_c2_�t���s:����Y����=�v��Т��9,�Q ����=�S�J�Ǫ��%����d�3�Y��Q�v�%z3/��.�����d���2g��P�6������$�D��q�9!׊��a�U��B�N"����!�>i�	᨟����h�����a!���p
�G�/���f�r�/���Ŝ	�}�0��BŊ���C�6{��?jw@�Q@_����r���s�0]]2�?�sh��\�+,S���w��l���1+���6��4ܨYM߮��K䣣П���mq�R�59�@wn���u=�|b�<K����	=�]�<��c�ƣV�8_��d���0k���l�\�E���o��,��<_c�#�ٲ�E�gN�-o}��ea<d\{�X�j��^kCVaeˍ0
U�3�Q�.��R�יuǼ�B�[qS������؊j\_��d��EA�G:|��=��H�wę���e�ܷ�up6���7�3��7�<j��2z��|�J��u��I�ו��D�׏�F�� 9����ʊ��T��nU�a��
Y�6�͝�Z�<���j���4�	�O =8�z
)�P��7zJK��M��"X'>�.{�ǝ_Z��\e��4�� �^�1u{���O�����q��m�iy�u1�D�{_� r	d�|)U:o9�,�a��cٹ�h�m�/�akG�Y���/� ZI�B�X�^�]�:�͘�I4yd�_ɑ��Ds�6� @�xN�����1l�8�-Q�]8�<��Z3��G��l�͇/da�B���i�+��: ^߁�4BH���ۛ8 �/?Pp�d9�:<^�#'D�w���P6Ī�����c`��k��{=O�oTLˍ�=��d�q�b�Bj���Z�A� �J���y�p��Qq�����N����F��eX6���|�o��6��;b�
zC�ꐖ��P������pw����5�i�dٶ��ɸ��u�3  ��ʌo �v���V��H�W_D�����r�#�M�g Pa�h(	_z��7Ľ*������2�ؔ��E�[��� �O��u��o�X6�#�TW4�˅�6�Y��R⌠�Ŗ���A!��m��°��]VĐ�ȯn��7��  ��g�`�<|�ܒ�^�1�5n�#a�����/��{�l{�
�`"�߽[��=^l����8c��<�J̝�I��7fӃ�2'�����Co�d��q�Z��v��)�*�7���b���A�x䞳ޅ�!�M.)�&80s��p���x��:�yw�R���.Æ��Qiډ����ڞ��.�	�Y�M��͚Tgȫ	�pf�.zc��!BsT�|���HRtr8�����Q�B9����@w[�痓b��>Q�#��i.pG`mNF�a���Y�����H#E*��(�<��:���hd�V�/���0"�]��o�3��ֹ�7��8���	� ��{q���'�,���=Ԫ�����B�)�Z)�#^f.$t�mv���"�Z��܌µ,>lPfK�_����ꁾ󌱲z�?;j֎��z5��˕� qE��i_T^
TS3�	Z3�ϽW8�inTX_��v��b5���1{�Ͱ,�^�������c��Bl��;�='�`�/�<ɛ���Ĵ�골ZE�����>O�(5�Muw*�4 ����s����p�4���1/����97l�|~����7���i��H��按'm'��*�.%����M�@�7GV��+T�2��\��� ���a*ֿ�Bj�S��L��[ .��0�a����3 Ї�{'l�a���i,WX�\3M�K��@�=�h������/~��d�Zt!|���\�!���/#�խ鼂�EPd��<�F�Ws�@"��Vi3Y>���T�W	
�^n���D/�vm�t��o�-�	Lg�d���3&�wAHLE�Rs�+�K�ӫ�5�$��	�;T��4�EZ3ьeJX4<8+�L���)2��>�W�@(	����"5c8Z��˔�͸�FbYy�����,v������#/Z/�z��|ۜ����?Vw��p/�kH.<�% y|��T\�:K?��L����]Af�MTV��Q�dz����|q���G;�s��E_�aZ@5º<uk�Ueb@�-eD_5�8���1֙��mZ�-��[�i}� JG#d�^:�a�ە]��+􏌤&*~U��lW/$XbS��m�n�Jv���w��ɬ���o�T�����C��l/�&�,����d���54�ě�&��D��J�	g�F�Z�`	,mǥ�W��(NCF��}��&�s���_:��xi� %���+�cBL�-0�}]����}� =�r�z�n�פ�x�"4�.�e����*�5W(��cC����J$�Q��Ž�ړ�A�_����3��F�ר��|>��H�xh�f���Z�-ڕK�ɐ��͹ٽ������E|w����')|�h���o�
�*�@����&X������`K�۸�%|�+LF��)uVa���V�_��&J^�@<��f�u$�N�@��� R������;�*�6SY5�d*f\ �_�7�I�v�����}�ӭy�r���\S�*^AB֘�ɬ�kd-	�ڹ����B�����ɬ�(c|����� W��tN1��-E?��iޔE��.ă@���_{�U��L���Q�Z�Ax-\��Xj`g�5��W Ș|�/P;ı�6����
H�[3?q�g�[���Q�%9�]!ً�Ɲv*{�7$=�#�۹lcm:��� �V6:�	�$R�Wd"�P��~�_���T_E^'��|1����� ������)1�5�!����|Gڜ\qt<V�������EoHWHJ# ,�J�N����,�+I�!� ������TI#���LP���Ag�Qtګ�R��3kӵ۳�Q
����7�GsMa�c��Mi��Y�w�]!�t���1O��P�8��#^�J|6�A�ܔ��ปc��L$��Dp:����`h�R�L&Z�sϟԸ5�"x�q��{hY�-����<L=��Rƛϐl�)Ø��8OA��je2��9NaU1 d�2.*�o���-!�����/����b4$�#W�c�����SU���X��(<�p���~W�iQ�祅G&/"t1�h{2��Es�����};����f	?Q[��m��ym;���؂(W�m����DѨ�](�d��R�B7�+��oO�;aN
>�\�������8�����e���4�`��e�[�!�OLo"�)l�b��{�|��/)_9#���6����9J�v�*Dm�k9*5+�c~��Ϳ�([X�Rܦ��,��E��怃��=����=
7HJ\,Nծ���"'���E�8mU~�o�$-M�M�<ex�cv�;�FM��J"#�X��4�j�3DE���=�L��4�g�M�4��RO�g�i�LsJSKZ�q�[��5��[�&cqcf+�&���Ȝ�Q�7�,7���@s�O>�^�`΂͈=J%ۜ��tx?w��:�-W�̠u��hs��nl��G�U�JC�qva��iI~ۗJd"�=��B�2�|�r ��+紙�w�I����h (�G���Ĭ)�X�S\gZ�C0�^�g0��2�˟B5"īLA�e���F��?e��Ċҭ�|���
U:<��������P�jKS�����
K�v#�leЊ�&*�m�^�/�����{Rp9~ ff��l�\��xƀ�)8<H4��9�}.g.l�V�;Gջ���m�P�����`�KS8��+~� ��$eۣ�+g�����֔h�{=�&��1��E�����ja�����w�o�0�*�	�7�3B�WM%w�W�PK�� (:�l�;q����=;�*����([R�2��\�.n�G�U/�L��k�R�b]�����M���/^&�͗�,A·�U|\��ϐ�����C)���k����X5ɸ�G��dGc���fJ'�3�x`�#Q�' ��{л�S�x蔈����͐�n��8��Z��������݆6��T��i����W�
�H���IA��k����<��'���"2�#,�Е%�4�^�怭=B�jBZ�7�46��- l�Z��˯5�T8}fGv�!gɫ��OE�b:����i^ {�ȁYo�QV�^p"��x7KI"{'�p�	-�	��o�+�#�<�q�d�y1�+�{�����C�휺�#�z��Fq��)�����:r�P�[/���f��@F&�@h�>�4�^↻��(�&:�)�?�>��d�U���\���6:�L�^�Ȟ FE솉�����P�q��	v�4e����m�v��a����L�U�����Qj���?cM}e2X��8��feFn(]�<�,v���)Uk����W�ՌRU��2���U%�r�_���u�y^����`�$�T)1&�IuN�JK������l���~�����v���D�#�/Y��*�̓SM��mJ��W4j��w+Q����2�����ڠ]�O�Kz?܂<ϳ�E;�J��L�������Ftۑ��f	Q]0�1��d���֬SDM?C}I§��K��o�$�T�Kj5�������]2�R� ����a���j�X1Ѱ7_��"m�����!C���Q�oܬ#2!���^�<2,?�zn��W�j���1:0��̜˔�-�~���t��s�[ ��O���!��h�h���l�����D8
ц�ȿC���u��Pg]�|�_ݸ����7������񞐴wP���T��^���젱��} � v���<�Xg�������+���&:�\�H�Q_��"���y�8Q��\B��M��fíI���"�	��v2�#}Q�e=,��^��7Bf����ӜV��-3�:[��&�����J�N8���w�>K���d�#���;c��^�3bP��%��4v�&������d{)���F�:��W�(��Ϥ�?ϣ,W�s~$|V� h�qU�$����� &%3I\*��~���uHQo���u:������fI�D_6���<�3�k0odΏU*~�./����r���!H1�|&\�`�pGM�13�0Y�Fu�`uX����XX/��uJ3c_2_.��id:��b7��k�/��9������O�F2�+��02bS�d��2�	m��Q`�����:KuǪ�h�[��t�K�o=�0n�E�ɵ��#���*j݉���R_��ԢE�����6X�� 
�Ŗ�=���ȁo,��~9>��������H�
7�!�|!���v�'�=>��4���[��V����LU�:���?;��>���G,JO:0�o��Oy���H�T�d��S^���̙VE��Y��:~q�H���l!"'�DY>^1��4%.�f��������d�Cx4u+%9[�&󾥊��9S����I{�x�S�|8� �tg��pB�K�ɥy�kM�E��3Ғk[�a.�����g6ߺ� lwϝ�Y�:iCW$�A�_��-v���
:�na̾:���nQu�h�?���4���^��l�~#ws��b���(�1o;����2�^>��W�Q��P/��eY�d�l2��Ry",
/�5��!VjA��`�!�?�b�7 V_`7;"(��׆�+����;]��w	|���?g�ηs�&<���o�4L�ᔶ���Lb�_����|�����L�9:��@!zlQCU��?�KԿ1ܰ볟����s&W�F�2�ѽ��FX{�~�u%��u,
l���q(��㛊�,w�2��7�a�V�w�eb��\1::�d\�o���~0~1���Y�SM��w �y��Yԩ덴۰�,��tR��tfy����������(��Fc�)�-PL�Q�ut�eU��p��d�����A�8暂��Ԟ�>#.J���?�Z�!�̰�\oĞ�rm�k��m]����^K^�1V{3��ȫgR?�{
�7�&l���8F���!���ɈM1x�I�2ۺ�G�n� ��7��<`[l�Y
�KE9�UF���V�d�sx�e��ͨa��0eL�� ���q���Cgp(���炢6�E6��	�#�0�#=�b�4�έI�]���!:{vķ�-�m�x`�6iI�r T�!?�9DO�ǖ2�(k޶�ﵾ�-��¦�0��:��; U����R�����\���BPލ��D��=��H�;2��"�y|��y��;��hU�%+�CNt��-�/m�:��i =~`�j<=o/�ۍ��J�������YU4���:�DO�$�d���`v��LJ�pM��Nm�u�k���=f<�$�zg�˪��x�/�_Xv��=\� ����b��	)خ�N��(�� =')�:�zx�@���|Q��{��u�KAg�}�6�,s�_�[윝D��F��������n �R� ?��J���_��_K����W��di*-���{�gS%�oS��O�`�R�K�t `a�e�Pi�8�����@+��lC�(Ҕ�s��� ���	GE}�Q��M���������5d˅��u�:[AK	u
�*����D��!�Fw~_�iB�k~B22�/,\��%�(���QP���x�K$����5i�c[tMJ|��J�'�
?�0|�|Ff��,>&�%mɽ�.v.�e_�f�]��N���l\��$�܂�g��=�$MJ��B_�8_��U��T��I� 8ɳ���9 ¶'��Z�h�qH��H+!�W���7YXwu�2�4�_�����m�x@c���[9��-��S��=�n7fcdq��D�˛d�}��F�*���|����!Q6����4(p{��[B�[k���,��X�Y v���"z��x��f�]zjPӓ��:�c��[��b��~W���z�V�XR2��EOc7��jbT���k��@K|U����P2O�u����Ղ+���ԙ��d"�~tU��-5#�ht$Hh��E���MK��l���Ş��mA=Ĭ�EmBL5���pN{�}���;{lu7_y#�U��T����mˤ��ڥ�^YD�3N^��V���~/����F'ڼ�cO�Q�u\er�!"w�����`$[tt����lg�~�S��zh�FE��0��0�����D��3�G4G\(�d��2XO^!��(*}�p�/������&eZt�9��j�C%�~��3�dϤ��u\��?z��yY5]D(�������va^�9�DV�y�g�O4�M�di?l]A*U�F\0�k3-OD��)ޒ3�`�O���팀`)}4���h�$�ٗ�|Kj��9�_����N�����͇���yJ��*�8��釒5A^7��FW����U�L��T�7�oxl�c�7.S��Ӧp�k����B�./Pa���d���.��
iajS.�"�t�3%j��I�g����ת��J#�<����"}�t�ڵ���\�ks�C?�\=VX��V� &���m�Y�"�������|n��-�אp{-%,jЅ�0@W�G"�W��[�;�ތG��χ�c���#x'��=�&�uqR�f���㴡�/����O��_����X�(�}o��0g.�ߚp�H��Xw؟���+:��գ�X�T���������4�`��Yp�᱋M.c���y�5rS?_",�+��/S�z��8ͧ;��w�?M�z>�m�DhR�XPt�'�^��&�����&l:�v��ן��k�N� ���I�M8�� =�����x���cF���E��/5.5/�'�O'� Ag�ey�]��O�e$�ʗ|���2'�{��TΧ�K��b�<��-�߂0nX����6�.��~��ᦌ�6n���:�_?��J����/�� ��' N�{p>����nQ-��\X�����=� 	D�:ʄcA�-3�op��}��7�<,�#�/Ueȏ���I\��	��.'���o����ڀ���+�q���/�`����YhE��S�'�wƁM����)q�8�U ?nsQ�S"<��=�S�-+�H������򤋥Ws�'M�<�"!��6V�Dm��y��)B����&��걑��m�Y�����x�t:���M�sxH���z�Lg������ĖiG��E��l�@�;r�|0�߅�;ȧb'�޹.�r'R�X���R��V�ǽN��DL�*��A
ޯ^�z�#\���o��~tಽ#8�\V�� �F�	ﭹ�z��6�E> ����6.����o#f�ӽ TL�On@HU�ǜ��K�}����ٲH����>_,��n�B���[��̈́���c���(���j�����l���hm>}PU&�88r6�!���!�<���gaԵ�S��MMt��U��ȱ7�K&��hn�"DE���^�s�p�t��a���k�� �;��v@//�����^����a�����*:�y�`���Or�O�\v��Z�AwQ��Wl��j�z��95��|Ƞ�գR^dEP��W?yPM��W�mL'x�r#r�n%���f��s6�	s�eo�Ǜ��Y��3�#=��Z1᠝��_��P��(��,�'�,�,\�_Dc�\M{��Uˈ�-GIs�iF�����]������K�[:��&o��f���Y��8xqCZ۠�`�SU�s��^ji�BhoU;�f����-T�AB�LJ�_�\���i=�K�wIё��d���?�Q��O"���\�Q�
kލ,8r�t�~�V����Z�}��CK�R/
~w; ��SK�E�
X���Ē������� �<KK"�_�����l��ݨ�&����m��U!u��8�&3e�'���v8%�,(�YW7��H%6s���a�"7s�����: 4��N�׉����s�;�L�K�%��E�N��z\^���	��ܴ�q��t)%����'�5
VIw���	R�(uIb����mo��[��%Ş��	K'}k��$-{�J3�#�y������ف�l��q�^v�_��%����'���օw�Lc˹�`����Pw�ۅGY+#GE�/�������~���Ќ���Q����_�a?�Vې ��1�7���̺�3�?t�<����u���Fa:QI��G#`��@eT=P�fA}5`c����)N�0r*3Ej���݋oz�v+rqnQΊ���e��Ӄ:f���D��Ag	���f����b�d�������7'�6�U�W�yvO`���e���ÁD�g���H#�n�:r,FO��f�!����u��R����&It����#_�M#.k�&b\Ϸ�Sx'h�U%�M�:��r��_a��iX��o��{�٪�)���7����sW�;9��`-֬	y0J8G�\#>Ƴh�"q�[��
��x�R�9�|M
b�ǭNߦ��ۙ�_�G��D4t!����)����U���9��=��۪xx)\R����0)Ll�w7�H@���!+�4Ids̑������-��
E�,�Aq�Z�3�\���qu;'�#�4�3���K�;��0���$�)j��M��&~5 I]�
[�P�ܖ��׾D��&��3�
�u�d��L2�m(Va��ȍ��P(:�/���}b�RH[��h�]�,���h}��NE�=�lD�������BT`s�C�
M�q��N�m�a'���pL�{ᝒzf�g�R�ɫX�=�B�zNNF���n	n�� �?�;�&6����ŀp�}���g*��L�B���@����e.B��A��Mxl���1_�F6��CycǂT
��l,Y�U��a+�J�[�-���ys���A$���T�ur���zf4�����o��-�Ù���fo�pY�;O{��`�����<���Ą�A�gf�W������C������bqeZw�/ʊ���Er5~��q�����f��?��f�(����7�5,-��"Q��*=n^_z�Ft���Jsﰃ��wXVY|�y��Kg��9��?�FF�U�0#~@���,�f���゚���yL��F:3�V��$[	��T$��!˷�4셷#+C�����?SO��}~O���u�RtM'����i��]G������#��S��o�I�ൾ}N���Lk@�e8�>�Sp�%\�aL��
+F���؃�o@�
���`[��Z���J��p�����Jǜ�S��[��b��9�-�i�}����NBT����د1Jn���c(]���nk�E'y�w�CPԆ�l��ţ>C���X�7��m���-s�Q����D����d���?��Oa��+:�Z�x�}g�x`�7��4��-i�� Y��/"��hT�Y����������z�^���by-�`t+P+�/��:�ԗ��$��Bp
�Ɵ�]W���񂪦:���s�O+�^<��Fa��������Y��\f%�2��`�K��11��Q�/}y�,�d3�TW���ׅ!���s�
�l'W�(�ohC���*}��H	h�D�[�������?R^��1~^@©��H�/uѴ5����M��ڗ�e��Zۣ�w��b��R������� t���$m�����"��u6��Pp���'��z�+9�_�D|�Ȕ����/Bp���x�i�U�/q��7Tސ2T܍0C1��S����S��X?��KEk���#R��=a�i�'\2�O�i��`������!ER%��E�G8̖DuI�/Qѭ2��g^���+��M!���ԧ'�I��r\�M�qc`�HJK��-��:\���ʣ�0a�ð�kk�Ƴ@2�Faq�#U��A��&;�$�4�׀����4ס0Y#.�s%�l��y���i%b^�m��0��Y�vWdk�~&H��O� ��bu��y:�ﲗ�ZbT�?\r�u�+!�J��9�4�f�g&i�y����%�&�$�;�\�;�;b�6�-l��2xh�n�˫���y�9#�&�1,�O�$+��c�ek�a߰�&e�qVt4EO?���ke�x�SJG���Ȁ*l$D\q7�>��q 	>������l
ol{{��-���/����=K����qS�L���n}��gn,F!�6�>puq�_dj	!�������{��ō�at&v��6�Yw��,�<��'�N�g;��K{�X\QQ���|f	`��td_����Q?)��Y5~���pF�kAk7��k%Z��,�,���{�U��8rT����tp��/tΩ�70h�,�� i9nY����(���$��� ?��ފ�����i(������!HE�:(7���b?b.���v�J�g���aJ�t�-;|DtKH�)�%����jo��H��Aa���#��&��>6n��c3��~S>��~͏*� �i3���B��o�?1��@B��M=�h�B��u�
�q,��*�����n p���2�P�}m�#&�o}�UFiT_x����#��zB�(���5��Ҏ�]�[�)��e�C��̰bz��u����x�� �>���{��јX#ZO-��;�B�݇�q�|Ps?��}G����D�8�})�1��g���\�h���(~�n��/��nI�]�c�R��TZ�*�8bGI#�B�]�Ey�f�<˧IT�#���g�@/���vAW��F>�dw,�?��R������6�G9Z
){��A�G �t�/����l��,)��Z)����E��-Ә�G�s�?��aܽK� s����cf!��)�k}eZ�5�S�,'�o��h^�^j%��y��_�i�����\�&c��*���7:m>NYȋc�tN	����%�)'�v�6�����<.������Hێ�����-��ώ^G��ݳ��s��n;R<�0�	����5���{�C{��c���v7;|:z�l�s��gA��u%�:�cA�)Ӆ���2�a��ɺF����	SjT@�^��(O��Df����`@'��\[�������s����B�IR�<�=�G�g���ȱd�6ɩ.ˬ9J@�'/u��b���Õ;��[��?<�p����9	�"FI�����e)PVQj!(	6�pHL�AaT�0ox	�%|so��m(S~ĶX�b����nӓ�ߢ�xv�(�k��U�.��P*�[��'��oGL���4<��'�NdE�C�A�CY�Zv�vv�f�{VL�W�1"�1�bxr-��eW�����U����qM�m�T2TU���LVI����%E�$�܃������Sp�	�5�m�V8U���2VE�
$<R����쁷������s�����s({�x�d�SB��m!ɭ'�
�pP�����<c��R���JJ�`�Y�T�Ol$�U��/Py�wUǗ�~ �{q�V�����g^Dh�B�G*���~�gҜ��n�L|m���|�q����a!ǳ�^t#�gĵp}�m%��8��>�̓�l����-��|^�z�5�6|]��6Y��"�/��Xb&6Q�"RҮ�������M|e�d:J��O$�b�����,}T�z~�=�o:�yd�ӑ���BG\ȕ汇�W�L�b�AC�,{т�}��P�`�q0b���jX�M���ci����V=+>^�w��Xe$��'SDB�5�"���z�~3�$�����1,A�&�z��mG�	����i����۸C�����t ٫��$���ݶ��C{X��h� òd�6���to4 0C@��7�r�y�*��./g�{��2��!Fk男�^���}�Ò���?���D�wF���j�MٿD���HC��K�fe%/mEtv��u˿��L�wc��D�t��7����1��O��B��Y{%W2^�`���T1�@�p[f���#����2�� �4�T#�|��a�ݩPV֒�z9�r�I�×3�5V�T�� ��{�����Jn�h��j�o�#��!MK�nH�l�e�?NWC��G�i��oi�2{�u�fH�W>�҈�n w��$r�"f���Nj�T}���3R,�mHV�^����G��H��J���J0M�L�����͌ZVN"�tN�#g�_
m:��]� ���s�
z����g%JR,C��I�f�|��5]��x��n���h,�G����>Z�*��	�Y��ɘ,��J� �ߢ̺�nӐ9zm��7�Aё�|����g��D�t[�D�6�l�pZr��9����+�Vݮ�Ga|d��=��r��?��ޕ%�I%8�����7�����W��Bw�$��pF3�l��n	�u%,�0ϳ���V��}ǩ
�Id��CC
�Ѐ�U��"H_la�.ԑ3���%���G�Y�nS�K[a�Ʃ��Z�o)�S4e���C%�k�x�����{� ��64n8���׵j8�raP-$q�77��\蒦�ML��k�כ%4�,"؇�A�x��@�%���Ft��ݩ��$9C��gJ)]�ۮ�}p��=`�9Ɩ��KNT3����r��e��@�B��À�Sx���f�)77w����i��
QqMͼ��mF $>s�i�Tg뮄��A0eG믄�6 N�3ل�3���A'W�-�R���x�-/�tq�wx�}q� �'��M���S	�Ҿ�bKw@q����
��<�2��ޓ}ʫ(���5���n�5a�`��v)<b�1�v�YR�H��/)�&�,�<����g������od)��-_�TwЮ�Ub�\���o����t��hr�T�J 3��M0��m�p��쭒1S�F>�5(�7Zv��D�hm� \�~h끩#%o��H�fvfȯ���K|NӉ	KS�)����������}_0lT�\��rOgB��t�����B����7�\�Ѡw��*�`�R���^*��A��3��~)����&k55���?���.x�kL�t����;�^�Ů��F,�R��M � c��Ƿ�ca�����R]���su1����qI��7f���4�yYcpz��]Ӷ?���B�����.NQ�:�o��Z��ω��]Ǖ(0\�~N�F(1Z��Bap��оKǵ�h@=�l�U�H�@���E
��V����s?5�pxG�|ʪ���%},�`,u"��E��l~,�o��i���l�`�v�#?���K{�r+�S��m�K��LNؖ����O/��xuGg�=�?�XV�g�d��9�d�T�N�/]P�d9�H����ޖW�`�X0���f㙄���CZ �zY9�e�8���>��]dR�b�����IN:���+�b�`X��E#ӕzA�X�"55��ꚒR�$�l�Db(���e��d&��\��" >A�