��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�I�;�b��v;-j�f��-1G)zC�!SRa��<���9��11�)�)�4�.�U��|t��-@3tt�s����}�C��)%^n�素�r]	��Ξ�����-'.Q�R$��
y,���DJ��S[�<Q��ŵ�Y(P������Xz��I�����m7�E�ED�2A<~��f��	<h/m��a���otd.Z�Bj�<��x]�
K4y�'��J,&�&�W���샃�L��I0�5Ɋ�B�o���[ƍ��>�Ԗe������\����ի�7�x�(�F�� ���Y}c��z�y�W<4U����,ao g� � <��ڰ�K]�K�~�!j�K{�k��'��K��oX��Jˬs*]Y���6�^�:d�� B��FKIv���/�������&���{P�[���mǾ= ����ch~�G�~c�ZQ�<{���8l�wM��!�Ά��y�N���8�'֮J���\���/R+^(r; o��AW�u�]����,~}�]�˫V|w'x��H,}V�8���	�����=&��Oru�,v��P��N�~��� �kC��wB�ՆTA2~����sr6q�t}��}No�����ݾ�~�^�c3�:�hŢ�T "��Tu�[F�zZ�K��@��|L�N6�:ֻ�~��>Җ���-�S7��$vx��+����
�ջ3�����|��k�'#.�w�c|�E���8G�im��(����}�%��-m7�� ����E�>�=CL��z���B�������s
�Ɣ?L*��J���C.���C|�k�ˬO P��C�:C�*#p?�G�V�E����%λ��{]Yogn)��/Y��/��1������}��e����O���S=�a�����	��ԏ�?N�ލ���F�rn�֗�q[QL��dz�ל���c�v��B&N(߶Is��3���!o��|��!��=ͼ���Bs}�$��p:�✮μφ$Q�$�/+'I�`A��е�:�ű�7�\�����
cz�+m &����/5'��⦖s�s$�?܅�V��9��kC�G{<�����SG��2���TlY0<E4����,Y����iU�Ԁ�e����V�-	L��/sl #��	��p��ԉ��fZ���p�υ��{C����@+F�W��p72�� ݅�aAYo:�_E8H�<�G	eZBё�-�ۨ�qߞIS�cu�z
vdP^��kh��Y~�/a8�N��;b����).�����ߡ�<�ՠrڒ��v72n�����A���6u|�_�w��@fVn���A3f#�p�ߪV]^	fT�G>w��29g�%���B�7���G_j_����Ϫ�,�Ti�x���7`����<���6���Eպ�miM~�!J��Æ���( ��W�U���:���MC����$�n�Ȧ;��b��d?��9�]�L�f:n%�K�7��+溝]��{
���r�^��U�]�v�!��^���9�tۤ����.2	�W�����$�z�$,k���z$G]zO@Upv�u~�5QŬ��*�Q��>ҏ�An ��#I	�/��D�������ME��ݒM��:�)lh��h�M�ƛ~"~�.�»�=�0\Is ��	n����^mtE���=����4rs�}�`UV�$f�,�fQx?��e�3�Ԗ�r��J���W��j��sy��7���v�Fw��	q5�+:~.W�~�Ć�zy���IFOQ������*����:ꇮ��M�*��$�%t^��=�F��	'p��V�%���P��d2ㄨ�aܫ&�{X<��؋�Ċ�S�u�+�=.�yo�xG(�m��9iz�����<u�8��8�C0����/��8y�l�̭+�ۃ�C�<'���XR��w�'���+�������x ݷ��m��>���ۥ��Ht໿����f�h�����%��-o�S��qY��U d޾Å�\���h�ʬ�i�=Am65
DRu�l��7��Mh��cF�q3��a(�v��~�/�qKEE��!6���upSs�7:q����YW�)�z$R!f������=��{а�.W�1����|vwm.2�L�T�j���U&.��X�5�;]�F ���j} {�� �&�9�"��`���|Bc�*J
�����.��G�֋�h?�T�0�0)��}0���a�7S=L�� `ݽpX��@HL�c��Jh=e??X�;���t%�!9c��{mD"���äL�7AU|�j��_HP)��w���K0�bi���6�&k��b����\#��J$�� �0X�?�tY	�%`ڷ!�0�h�}�wĊd��42zI���Hd'�o�G4���Uj��8���ݎ)Uu���q�`��*��7�U%�rk�J1V��ʽ�*�V���0If�\�� ��ЃS��ܱ[Y�G�`Q�a�"�Ѫ�A��5n���O�րq���ud��m�p�MYB��vuS��K�y�E��q�?҉�� oY�'�!oh��G;6�L��L��z���w���f�K2sÝJ6Z<pu��T�pC�siz���mU��u,��M O�4�*��϶�l��c�����yU#^wh�GDg����!Y�|(����d{rK*i@�����04i���T㖔�D��F��ZÆ�u�T�|�iܩs� ���Ml�^@d\������K4ӊ�z����ttLR��݃ ��`���_�sS��bV�a�ܡ��}q�&שnhne��K��h��"��}e��ҀZK� n��E��
���J\��y��m=^�LT#�`�H�_�	u��s��:~}ȣK��7HC�y��?��c���9�W >1�C0d����ռ�zM�=B�|
����0��b�j,�v��`!�����N�����
e/^ffH����!sj���� x�J��f����Q�,3��Q�,4WA�g��ˍd/"�:XH�ct��}�ۖ ���?��C�P0�a�NrMRhA-{�p��u4^u��Ijq�6�n�I3���E�]ε���>�=� >*�m,FdE˙ٸ�?��q���b��gA�!�8mkA��8d^��;�-|65×�*�r���_�M���`[�ߖk~��R��Y�_09�>��'[�q^0�5��)�.T^hV����7�p�{����9�Z$S����@���D�罀�Q_d�|��������.�4�,ϯ	�YEk8s��������X�q���3eCzw-g���cF>��(~�`�}�\X����l'fVX��Iݡo��چ!>O-�����1�Q>����޲8c��k��8����Zk�wZ3�H���q��[�]���N�׏C�_E˗ԟ�`�{��攢��ut\zM��ncq�e� y\P�_5y	ˣ�Jz()�|�����+z�(�r+P�,�,��W�V;��0��d=��=��l�K�r�#H���5pd|����������Q��y@L&Tt71T�]u�-[��~-�F�����C�͚�'��/O���'��\�|�ֽ�_���5���4�~e�Z�ã�`�9��}N��9��f��ͪ�~�]t6�Z�-y����4�un�Ul���_���	�[p�S����s�^�7pƲ|���[�p�+����E��x��F^g��N�W��w���L�X��gK��Vc>�+_B�[��@��؋�A�DK�;���!����||g�p���r_?�P��ħ�_ڡH��;� ���U�!�b3xչ���mE��\Qf�$B3Ԫ�������s���=;-w3X�'�B��l�b���X<dS1N��tJ2��[��v7�B��������|�VP��n"(���݄�s������NV����Ck��\�+�����o�QipA
�X!�y��Fn�.��p�9tO���(�x�D���cG�Y�蕰��˪��]�6�~Gѣ=ը�0h��q�P��5�m��<#�c��1�M!c���g�Fԝ���\���ě�̨&����ǎ�V��I�x�6m��E�:T��:_d����)�I�}Xw+6?항wF`����FJ���׫X��E�)�jz��w�E z��Bk�x��`����H��Fk�I`pM*���P��Aזּ_l;�L#`��e�ʹz�\�_N�x$@t>�ӷ&S5GLR4���s�	��q�x��+����E��fK��"봙��l��n��k��j��|~8����@�37��6Q�j}�ƅ�9!�%=�#���Y2 G�ct���\`'��:y΅
� *	/�m�����\�>��O���0�+Ӗf�Q�	Q�|�����Хֿ�u�>��]
�Ey�>�{�F��&���c�7�� ��*��#Ŷ�A����t�<f��ŪD����m�v���Y�,|��Uŀ�F!ŐШ)Ζn�#f�C)����A��sҢ��X�%��*��i�)����N^:���[������L} O_��>����h���;ي������M[��N�¡��T��I)/")�Ӝx���T��15�=pj2��t��[����3b���������`��	sY���$La�����Q��&K� :
¬*:D
�]+ŏ�N@����E Vc+-�dq�5z��ʹ����w�9
m���B�����z���^':�L�����n8�FJV�z<��1�W�K�/8㮓>����c/[���)�I�9����y��g
TX�cMU���D���3Ũp��C-5虡�qs}��{�( �3.���Hq����=T�ԗ��HTK|ˠ�y#@��=V��q��?�anf��5q��..p�T���r|��-�~��$Q��0@�����D���xÒ�`���~:J�����pދ�-	Z�EV�rҪ����#��y�#����������V�ˣ�D����8%����<���7 ���(�b���
�ޫ��O��!VSA�ޅ|�ۛC�`��}��7G@4������N(� ���*�Ĝ�'��׷=Z��jKY�`��d
��y��ÜO�S�,�^ �"F6e�6�"�����
@��[l*��<��}�!��J�j#i����'۪�tu�nm�
k�4�����+DL�*o�|���`� �vu���YFTy�!*ަL�l�Is���N�x5��F��*C�;�X��~�\��ݮo���.D/Q�O�2�L�]��cC�������SI�jB�.9����U?*�=��T~��H�|�{y��<�����_�������3��<�[��FߋZ��1�@�he�&����g�hv�͍��e+H+��6�$�]_3��*(MY��O�Z�\9�9�d7j�������m�)O�aBP���.4���6�8���?��_��O�,o\����}_a��E�+��5�\;nl���A���D�W��+�(����N�<�"�l����׌�O*Y��2KE+Sk�K���Q\��3��f�-*i���s���b����WW���Z%� �)�� ����pb�$��@�6��uH�]
�v��Y�W5�hӞ�>�B��4
��?�3hIFb�`������jp9�,�����Qw�jo?�����h#�8�:�&\p��]/��a �QI%f�A����_n��$'�
�[9D���~�E=(�����{O)�{���x���Phou2�`�L��9��^�#t<��.��W�t�J��q��0u��źr�T�`J�'SG��?��ߩ��������WW�t����i��k+�?�mB�@�w5��CZ���{�YU�,!��-'$es�ks�g!���Ӳ4��Jﳭ��9��_$�u^�p$v�	��9{��ji%�4'Fo���(4�;)_���8��+7;�p� �� @�/����L�1���F�X�e�3#�
A�S���b�5	�n����u��'��>�"������o貯v��Q�����m�jG�$�D�â��\�A"S�ޚ����7>GT�U�����c���$� l��L��M(xH���V�˞���Y�;�j�/��<���P����ϯ0n��ȥ"�%Yn�P�a�k��%a}�G���/H��a|o�V$���ք7D�h��~"�>gmOΡ�D�F� L6��eA5�[�fx���狞f����	��N�P�1C�!���$�ͯ�2��A��q�'����c��Cv�&�Bz�?���G�(�\pR6R1"��#ǔ�hu�=#�u ������fo4 ڣBg��$�2+1�%� ��5�Q�`w�L��>��/��ǼG i��}� ��_�ɲ��[,7��W�)�:���f.��Oy*���ŝ�l�J�ȩ�B�:;&Z���)~���x�8u3ʓ/3�@Hb�|x?���-o����I
L$���l��	2)E|#�G_<��~q�j�Ѕ�hD�h�$|����ъ�g+�nɗD�c��mR���;y�ݔ����3'���"Y�|J��s��~����*��S�4c�]���8K��C+:�ݚ`<0�Xv�ZF�bsXb�3�>6n �.i�͍�;�v2�#Tx���@I��K���6S����2j����U�ў�4�a�
�-]a��L�qbq��I˗����z^ ���$f�בv�%
��AX�n��f�UaTr����i�;�j)��r(s��ȠfL+�ՖƑ7�wJY���qJusz�|n�Éh8&�%`�dw����-wŴ���:��$w��
�Y��y�K
T�W�_��/A�Rz�A�,�#��im�����C��iE��Y��E����߆��-4Z}��E�N`W,���9��!�\@It-��ڌ.�G�8
�L���E�ƣ\��.Ef�>_A����� Eދ/��%�S���D	xf:��[��t,�~�9|�Q%Zۼr���7\�iPI�`�lŸ��I�qލ�g�	R�$�gX
�3��~�λ'S&5���Ǣ|A��G��kʪ���p�h�.3�k�#)f�E�����8p�D�M�r����M�$C{$m��x^�v+,��kk�Z|��Ɔ}S��� �Ɯ�)��ws�g���6�3:�s��I��H����q���2Ý2<[K�lb�����,1H�LCuV����"6��#)�!�d�|]����[fx�M�S�V�v�Z�d�G����j�j:����.����m�.(J�78�&��~��=�C���oN*E���Fg�;��H'��܋��iq�H�ZX$γ���5�3R(�n��tɋz��	�f���ޢ^���΅���J����V�(�c����9�-�lK8[��k��˞W�8=�
;l�d;����d��NR���'�Q��G�O�"����
,x���F��Ĕ�1�+����	�NA� 	�.�@�)���[!I��=9�~ �Y�Zb����sՂ8����Ƽ��U�~kd����FNC.�?G�|�{ =�'���ys�����}3��9�Ӝ������\uW��-~�EA�7����5T���et�KJ�Db
�т������*s�V��������ԣѮ}'�n�` ���ס�:������.̀�ǈ��c!&^���ݡ�3M�݇�`��z��3�f�F�}8/������??��ED38�����9°����I��)�:m���d�e��5Z��];�s0_S�<,L��ϩ�!)����x�|��E���g���f��a�� h�3�f�!v��dK[�齰<�l�L�=���트i���\���mSqo�j��
��*?!y��&#�C��:�%��':fSA�y��#%,�w�
"�>a�����NM��#��&�����` ��!	�WEM2�=��د��Y���hB�yxl�s8zS���)���91�cx�!oS��)�Of� �S���ʎԽ�)�*�)E���g2PL�d�zrT�1B����_�c�P
�(���/-]����)!@j��pf=�!d)>{J�}�N��8��Z�uL��NmM\�>MA����V���ӷ�s$�5�_�KЬ?��.,w"-o���>9u.��(���#%7ǔ�v�?v�ċ����޵g���Rr��t{�.xYs�1�6;@�SX��(Y�X�4mh0�u�c����w#��ӏ��&��8������i���3+�z���f�i��V`w*�v���'�\�%U7�!��F���5�k���.��߄��YD����WC�n*�BR�\��yx܂�������BAG�.ν�Ui����g�;H����HE���2�Z��y�~$�d(��X�!(Ӈ�2�E�Z��F+�g�ԿZ������kH��&�ww�d���e(1\�k��k�E�5_�r��
Ԅ�Oj������Y��=��Q`��lֆ�"3���Xs���iI`Vre�g�B_�ɂ�N��\�1Ś����;F~f�MOB���]�ht���C+�wa���%7ߍ��"� ��������b�	���m�Ē��PZ�T�r�c�vZ&��@	��%�i�K<T3FJv�b�ӠmJ8Yrq�l��� #�hLk.WF٨���1�����������B����W��bǋ�z7G�#@�M�?���Y��XH�Qʺ�hs*5�W�=�w���Y�ܾl���,�I����M8&/����[g���1���ܔZ�7��	�� \\/�m�%�>a��ޑzV�w.DL���<C��:u,7�q�=������T�����?�s[k�x!�P0~'��|�W�$H�d�"���Ј]�_��-���U4e�
$7�+֏^O(o!O�N-0¸�7&��ه���[����gN�TP�#@gG͍��6xm��+t��c��~�kZҹ*��MS��nV��,y�wn�}x)s?����j�cb� �v��3qu��9���^$�4���`g�U�ϡI��a�/i<�����U/j��=�OV����[ԧ��v�|�<W�ٍ���	I(�4�FT�/�۹�����V	Z`��_7����/w�w��+�&D8��2m�w^��=�V�����8`]<��� ��C`+�CY2�_�j.� j�r�R��Cg���w�O����/S��#�Obn��-at�1IӸ���Y7,.N�z�6}y��ĺi-Yb��,p��l�Ç�����Ze��m�+9����Ǻ@�@G"�v��D�
��#bK�;y��;�$J��|�Ay��y�����G^c��\,<y�A]����G�
�	�NĞ�w���N�z���s1
�U��T��j���� O��BU=����T{�>Ͳ�&e?�D������3��9��R�᪊�ĕ�$w�$Y0�_�{���'i�.�s`׌��:�i����i߻8Eh[�[Z���3c�(vkky�.-0�ė�چHI8�����f_��CvU�G��)��8a���nR#������2)pjOiHe�7�=�w��c�};�`̽�;��ʦ�DH�m��60Q�Muj��G;�H0���cZ\W�M��p���D�0�Q'��$�g�鿨./,��}�!
�(-�rQ�+Xn�>�*�^��3++MH'��-?U�����x]�88��5���&Gk`����H�k�t?�j��m���!�T�C�hk�3��W���-�f�`��)�X��z�%�����S����H�T0�(aq2���r'�/���
����>c�@��$Њ@Ύa��ūR΋z�~��S�^���MV��glöM)'�Б;-.H��X|4I�N\p�jL2�4�l���M�2T�i���Y�c�2�~.���?wn�5˛�&��
�	�|zh���Ϳ0�m�j�[��{2�l��1/f�����y��|j�w!����S���.| �$M��&���|�%9c�/�H��6K��Yw!�'���� ���&2�D�S�,�4���崀���:�i\���(Yt�O��P8'��M3���k%𰑩sm�$��g�//��4/h���s#	7��Kg�0�>:Z/'��q�S��/xm�$ȝï�G���+!6�������Q�f`"y�vg�Rj��R^��Tbd+�
)�s�c1�^��΢$U�����{�I���`UI`�<�'D��@�,!�F���9-~�m����APH���_Qq�'�S�fC��O-�,ݽ6��������<alyJj�Tf��^��q�f�f@k7�|�@"U�+�`$��	v0N��\bΠ�[�۶���G6���l�\��~J25��0��3����$�[��d��QC��=��?;6Ѫ��{����GKA��Y��=j�����+��O�BgWB�C��Z���q2��e���f�.�� �!����e���o����[-�#�������歩<܇�� �������Ғ�c�В>��Q"Ĵ�Fg2(�SI���A�������p+T{��1Ǹ����,�%e��Z#Vx³���&�G�����\w�i��-�ٰ�-��[J|���*�����
kә髯,et6J�c�3�FA:j�Ƕ&������y>�ڹ8~L`��gd*^�������B;�c�
棳fQ��vo閒-����	����Z��J[�$��L������a)�H����d����	�R��H�h�u_~�P�2�4����Xn�)��e���0�b��(�ھI�	�~�͵7<��;�[42�O�D�/�������`�\�sÞȬF�8��΁�ަf���S}����p��	�Q�4#�����k���_ҡ��%P5x/��c���ê����U|ZF�XX�}�il�:�TK�{.n�c��B�
Ĺ���X������j�%%�3r�%�/�[�~T�^:�%%Ma��[��e�0iY }����'��%v��8<�|.+�{�����������Һrf�.=���F�',�/#Ѡw�G*��I���_�����qI���8��
?�oRUGh��A#���*�Kȑ,��h?=�Q���V�g�ׁ!�ٵ����B��OW9:�'���_�X|;��<���M�~��:	!���*�?4׆u�b"�����s5V4a��i��d��7������U82wSjh'2��}�wӻ��
pZ��ڜ��#�M�(ޱtؐq�'lA�� '���Ul+o�@�sJ����L��`.>}����@���Xk��y��9mp��f��T��
7�Y�Eb�����i�l�