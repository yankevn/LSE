��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��|��b�*=��{������[Vt!��L:�RȘ����!�T���	���m��I��oYC7��pz�3���?���~�xPC֜!�%��fVf�kH\��A0%���9�qSZ����:'�ض�VIǵ`3��E%�,�-Ǖ���3�D�����+?��I�$Eɴ��$p��DtqC� \��i�H��PN�����҉~8�Y|�TM��kˢM�q�2�$-�h��2��I��!�-��I�5��[5�]�����#��*�o�{��[��b���#���I��"�tk3��ƨ\�)��F�Ң��@�vc�/�;���4��dӦt#l�Ŕ_̓��g����mHm)�#�-*W.d~�e{;HL��̶U�	�u�Be��E> ��{�\}��2Z�M����_ߺ'�4��f�`L�Xt����c½SpjWx`�Ȱ,�����d ��\΁C���dΟ�)���Q5v)?�ff�w���	{ʷiM=ejҝ�
�b����5�)E>�m�A,|���o9����+�Lf�N�9D��-����w���ri��Ru�����A�<��\l/`���:� e���FJ�i^K/Z���*,f�� N���31�����[Vƨ���$Q�+�ߡ����]*�0�G۲���NQ�����j�_^�Via�X?ü�/݆_i��e(�v��5�wm|ÜQ�����}�"�+�a�_�cv����4_�,�+ڞ����p�1%��b�XtSc�^���H�#������x�*n�FN�����)��ɧZ�_�y�����&�]s����MiD���j���&t�[�hK�>�=�}��o�a�5"h����[����q~O��F��X�@��В6e0V����[y���qܡ�C4��B���`�X\ D��������QVe�3:6��O�A:a�?�n�ԛ�D�x���!T�,�ᘇ2өz?���_����piA~�I�ر9 r%�B��ej������*�e��D������e��n]N��{�e�R���Z�,�V����o\Ŋ�CO�'�PI'\0S�9��w�a����{�{o6�*�`��Ms)�kaϕz�K�����=���W�i�3��wظ���_���噍L����{�=�q�WS@P�#g�Y:�1\���C,�kPV�4c��k��D���F_x#�Mڨ��_i=��P��`�3�g�ޟ>���-+���Y�J��g?V�7#��euW�ruRa�<9�Z�s�n�4{Zjd"�xʽb�����)���"��yI�s��I��5�h��M��1�����&������4�����ՔH8>8Rh�� ����o�XX��
E\��p��V��6���27��O`d�T�s�E�m����֘dŭ�j8�B��]uXT����Ta�ЕB��Ɉߢ'�]"�6�Fm�����y;�!�7����2uf��D��Z�����
�K�S�0d����WwJ�0z�^B�!��Y��*$��j�w	���1xb�!�?��?�棱y^ӧ��XB�,N�'��v�|�iH�u�#�Bw�?�zv�2�ٓ�n����*�8�f��]�w}��}����Mo�js�M���/!�|⿦�V>���غp��i2�X�Q`,��d��#�1��F����1���fjO���5���i�&@��/U/�t�y�|�|�j1
S'�:�~��n�����E�<��� � b��
��<?����4�����C��t4��u}��qK���ɼ�q�Q��m�wI�.�S��Dd����9��u꘶�%$@jW�����8)�s��M*�ɒΎ
�TrĀ��~AH�8��k*�˱F�Ly�y5��5����<�q���F6�C�����-��/���Ǐ<�$��j��W�t��=hh$/�6��x��J�����t��~�a� �����&�81�z�l� %��GG��s�;b*�J����wb�$���*&�UR��2&Ff���w��0Vc�"C�φ�����$�k�,�k8E��$��%�׆����v��v�Y�o�;�+��ю����R����n�	[
��G�b;"_N���������a�_l���߽�;�m�\h��È��f�A���(d�!���� ����[9�9���!*�ǒ�p�R���G�*�{�-�!��X]V݂G��JTW��$Y�#�{5�O��o�����.F"#���3����-dK
��kO��G]x�e���y�ݍ6�1!ӧ>U+��G��'�Iy/w�a�)����C�׬�HΘj�X����fd�i�B;�
�'�t�F����X��
���E� ����������Eq�ol����5��;����h5�j��o�l=��{(X�y/�ȳ��U'�K\M;3@R�܄�����B��������3]݉��_T�m�t�.�`�;��m+i>zyz�_�D�z�[��V%�+'��.���L��}������"͂b�w[�j!��=�]Wj�_R�_��V�>��C�eDQ%Ձ��p�⍡�,�it�����D��=�K�������Δ�����:j4�
��K���b�V�g��D7~�ze8�U,�"0�ߦ=܏�����t��]u6ت� ۻ	5�$#S�ߋ������>A��YN��F:�7_��]8����NH��}�z�H�Φ�ڐ�hUT�=�Wƨ�s,
.���KJ��ig��'T�A� ��2�ޛ�I?&a�$��󧱏�G"�NOC����>��l����3�vw�b�&��XAa"����^���?+���A��y�Z�~<h��,(����i���:҇�<:�ڵ�6)��$�UU	�M&3ww�{Z\,��w��x�'�	�5����fP�+�K�`Տ����2���Ĭ��5�u�fR�JM�}A�?OwR?��/�p�����17F@�#���&��ɂhE�1����b�s���^�q9����$7}��^� #���'ЕQ����m2�/֚��l ���ǐZ����Ւ�Wx+�uhnʹfN��|҇Uby?R�u�ä��?�1��v���`����y�mf;�¤h�|���ظ�YW=���ЍZ�h7G���H︺Π��w��<�ŀk�oG+�*�?�ˈFzF;�i"����i��Ȝ��v����C��o���w]�q$���$��r�&��f�G�	�ɳ���+[hZ�:�C�����Kx���e���$i�D;Q�=X�������ZB8��t�Ԩ������" p���6�����+��*�K������1OQ?�N�L�l��h������_S��t�쩶���-Cړ(WNp+~�����������!�o���7>�y���z1{��qQ�Zax_��!Ґ��%�X��I {��{fl��]+��΍�T�L�<�J��Y�<�����\InI���9�����+欸p�g�n�4pb�)�`1������Y�$M�]1����
\���� �5>��O���D%0���o���!_�gfD�ˤU�?�#y^�x9۫,��{�,1w�%�#��׵7��z�^d�@���`����\@��Q`�IzT���k=���O�~��z�@�^;��ó��q�W���	����@���SdM�p�ڔo�b���6o԰��|��˃x�6���x���߼��e��@�ꐵb}qq�(2u����MH/�U{?H�L?hmHv��ĺ�߽���F�:#�[��^��8��E��x�J�8�EO�
�	q1�7���v�AG��9���6G��X���`�E�y��-�	��}��w���$�7����WEԵ��v����{�$ܫ�ŧ�C¢�H�i�|��y2|�0����9ʽ��X����ւ�J̢����fj��*���n�k�=��JPv�w�A¯�Vb'a���B���6�Wl��Zl�J��=�܋�c̅.d�E��/�#���� �D!g�Q
���9���E�����u�ƿ�����D�.%E�LPq�Y8�Å�f�u��J������-�����Əa{�R���A��ڲ���I��l3��z�lI�DdWlT�I�	��?�ɜT�Nr��F����7~[la���9��a��콻�і���P�Z:k9��yq�8��׍�.�Rr��v�rl�fz;~���<|�#�Q�����B��9ғ�FV���U