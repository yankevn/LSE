��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~��j�w�9f63�cbGr\�.��A�o���M^7��(� ����&���z��p?��
�j~�#�j�˝�k7L�0����T����{3��́�;vj#\��ݬJ�a�~?�M�s�m%c��OD�����c��V��G5�m����E\�Ĳ��K��tAL!�{8�h^�őT4M�zS(Vm=N����|Q��QŦ��el'���Μ��� Y��A�^�Rz��0����������E�G�Ƀ^�-}ǲFx��XU�U��lpA�D�k�������mNZA��sNu��^|Y� g��zD!U�bxO�\���ѝ�6�>��#ľ�Mc��˭��٧Ƽ̄�ylg4�����X�tu��H��T�F;n���d�֑K��e.�-�6b>|�r���KcZ��{i��tfp?L����j�W]&i�Ynl*���j�5/������t�P��X�O�x�����^���̬C�^+��GΖ0�5����mƲ�Y���/�d�0@`�hn���˻����O�J�m�/i|�n(ḓ6xg�<S٦ZT0oD�@��y�^	%���?V� �k�o�V�����*]`(p�P)Y��C�Mm��1��ve
ʭ�Jʄ�^Gg����^���]�_*�G͍w�w^˩eX7B�e��4�>�Ng Ƿ.>H��͍WJ���g:r#s",ϲ0��	�P��%XK���6��&Ǉ*1Έ�$�\&R!�N勠s�]7~`���fs<J��Q
X#$c:�2.hKYx��L�^�o�_Z=e븲p��������(2��kH�'<��FA�0��s��B�����ζ����>5�X�ez���$����H����QtH��ߟ �E����,��LB��M�������@����^\��"= 1^���H�B9�}w[*�Z/�hׇ��à�L�|s�xj<UV'Tҝ$�F��1gE��yWR�G����3�qN�y�ĸq�����e<����.�4y�i٤������U S��1��p3`�F��o��Ql��4���I�p���]J�O��~{R��:�!G��l��;||B�T����cJ|�ykɁ%(0��S#[��v�X����'ӵ��H�/���O�V�]@��C)�sP�:Y�?�g����yS�^��S�tr��!��SU��9x/��������*:�Jr�����n6m��˝}�*���+"+�,����F٦1���!*�`kbb~�X�������%F�T��p�}-�X�`}Z���/������T<�&�U�����'��0�VΉ=�$�i���i�_Ma!B,��cD
Oz<�Ѱ\��/L�e���!�^���(sNo��`+���"��8�����٧��D�ݡm?j!$%�%���D55]Du �ޜ��kR<�?�*W�/��&�Br�7�0�o�͟��+ASk�d����"/��sLK*E9kCR������J���.k(��^qs�}������n�" ��4��&cjF����ZQ�x���1T�&�{�Jw�z���VҤ���T�v�8Js�K�9�O&%��Dk&�/(�)P��.��ù�S��&����Si��Ƥ
�
5.������:ӗ�Hh��,��֥�vHWG��?4X�h�X��N%���9��5�y�Y���7����H�I��V\iloo�8���}-kO&�8.���0�z,(��G�H�&��;j8Ѷī���T�	��g���T���dzAK�.�&=��������j^�_��7��[�Wt;�*P��j��<6��x�J!����ݧnB��#�t��#�?�{�m�Ի>A�����>�ሂ펆*0�0�ȷ����pc���n�j��j/6]�F�à����a��'/��L�d'Nރ���1)�Z�s˨q�d�_z\V*^!NY'�?傃�Ù<�,�VM,U�(K|�E��(�	"t�~^�@Pc�'�'��۷�&p�Z�J�Mu#�S+�r����Ҿ�<\J�����y@�eT��t4�_���*��A���v�<�����������\��@x���W����jj��6��[tv�71x��}J�w�����4u�1^���~�t���J��B��]M4`Zs��ә�)�nWГ'��&O>��
�Σ_��\��)9N�tE\�Ϙ����{�w�N/ʯ�k��=���=��K�ӈ������	R9�`��yOKX�h}Ȁ�U��kY_>T������.j�+��h3��ej��t���~V$E��8u!r��rV��.�MBG�yC�H��*<��M�r�c�W���3ma�S�^	�no�W���h,�����YN�(�i�4J ln��g�
���m�#����hL������EG��[h�<B緘�X�e�3�����?5�E1����R,n�J���[z]�-�b�{�uU�(���Z�yk?�"j�����F�Ϝ�Wp���������6�m̆uK������]y���k�����O��M"�{T<�O��m��?gڛ~u��9�.C$���eW1��H	�<`��o����J�8��T�5�fo��a#'�W_�����dPha���sR�@k��<���ȡi`ҵI[,�!���{�@LL*�"/*6�����aE��Yi+L�X*�d��&��;��hV-|���)G=�kGt�k��[W��ˤ��9X��)�R�Q�\1Z�x��#M��,K�R�be�3�4οb&u���������6?T.�F	����uAx|�趜�Ǩ�Ō{���i�'��[I��1ԝo`S�г%A�
�~�Z�4+�b�N�Fs��� �������v���hmȝ+��P�O�^��%�<Z�qopއy���R�z�˥���.�c���XR�w9��E��b\`|��r����V��e��E���x�Ϊ�g���;%}T�_����s��&ߋe��A�j�FEK��[�-�Є�AuPA�E��%1�&O�������[|�:`/��P��c|��6u�p#Z�v~N�B����o-'Qk&�H����1��ߴ9wY�~��`4���)�����u������j���<R���v��5��3pf�uY�
�\w����a;���ʤ��y��e�K�D*�.Z���ywAu�BS뤜�7��`��[!�H�62��t�s�P7?�x�~F�:@*,j���� ���}O��O�Αʅ�+�� �k����J��
�':H?���e$Mg2�i;V���]!@oިo�s >��Б}��L|.��L�4=�
IV��ǚp�%���Nec%��c��[U�̡����V�--D�nb�C����C4�Y���|٣��2�����Cp��e�Cj�w�6C�̻��]���װ[J���9@FVǴ��Xvv���q�#�I0�P���h���cy%�7�KF1L��Mª���)�J
!�jz���Ys�m�cK�)���)��\yh�Z,�7�3J��[N`;�΅�j��=$�V3��P0�f������W����<���19��\�6E���k�XF!���x�4�m�i�MM��
�s���!_װ�j����� ��䮅yU6t;���Λf�ϣ4��,�Q2�j @(L8�y�n���h���� *�m�.��1��J�sco���R�_ǌ\x��~#=�Q�t�8�b��K,.��wB��uk�o�zՙ��3��|J/q!l�꓂�E�������1u�PI@��Ā٨.WmUe�3&�R�&ID�u��t*�ŏ�9©#��2�:�Ĉ��/k���̧��sKI�){b ���, Fܖ#ܤ�b�����ʂ;�؟Kf�`Z�{Ɵ=�[�a�?�v�+&�j�ғ/�zk�"��EP��TL�7�[�Ac#zQ���Zļ�����H����wPq��#�A�q�Dw��rȆ���%S�Q�7X�&���a{�6����L���pIt�yB�!K��A�CQ�yc�G$�S�^m7�ZG���O���S�����������d�����k(�yS~$�>�1_��������3h��itH�^�I�9�k,���!1Ų�=�c��4u�f��S��87�����E�'��
��MW�d?����B���t��#3{*�	�TA��K�~ =jR�e!��}A� �߈{��X����3�&-�I��!��Hԃ�"��D��A�?�Ⱥ:�	��o�m�ȯ�A�B�yݨܸ,�x������$l�SR�����kc�]@�k���h�(�8Ff��k����[�Zv�V2lee�+>,j�}C������g�8u�	��ۦLd9Z�M�C���%�R�v��]��t�M��u�`����:#�!�5;�堸�O�/Ur�&� �A}��6���3D������L����}L�Dĺ�A�몲t+��Z!'�������KR �]k��}"讂md���9Ih�%��=�(������j�o�y>�����e ��۩n�poH[��?��?C$��Mh�u) ��^���j%�/��E��Ziy�$a%IJ�c�ֺ���Ǻ7������%��D�9���1k6��-��Uį&��'Y�b�"�;H.��c�	��r<��^���Б��	c�Ֆ<S:`��nJ~�Z�:�P�UOK&��ӣv��0�md�5�����������C���H}�i-�]�&Hg�u߼D�&�i_ˉ����,/�_�MA�X��\�g"�mH��mP�=��ã��R�����E�^%�N��1j���I�X�ͦb��&Oq*ȩ��O{�@U�������,��q;8;fū�=��Ђ�@�R�a��iZ/��%k"`Χ'�[��L�q~��21&�YG5a���u�O�@E�K��G,}��g������;!0�u��12ߣ�ل6�����#�wJ�w�_�:Zc�Aq=����>R�L=�n�����q�qY(U�컎�e�
cg��F�i˾ގŤ�35YU��ס�XB���$X,wS�Zzs�M���ȳj�.;yZ�]�|Ӫ�M�ńi�H���8r��Wj��L"s�K�+�!8��@��_�?&�"� ��j��T�R��	���A�(Lr����p8xl$���d ��	�Y\�9���B�Z���"
�����G`��~�Bw2�O� +p�_u�� 1v<�gY��7��K�Ȟl�F����Kw��݈X��`
�ѩ EH�vX���Sʀ@�I��#2�e+����R�%���{����%?4�~n���(cX2�0�k�!lG�	��iac�n6~���7����cv؁`>+Y�4~���;��	gl�e�d{c堆|�03�0^2O��JO���!|(X�ŰE 0�U�G=����{��-��a>�����ि�[f5���K�r^ǖ��4�0�;�$�G�tǮ ^30�_�6|L�BnW���!}t�C��G6-,���9����y[)ّ�w������J��8Av�j�Фh�;�>'�Cѿ����)���D�؃��z>�!� �]����H�����?Q���Ȣ��4|�����	$Q�9Ш@Q�c�t9bwP�"���̶�se-܅&�� z`��$J�$	��Sb���_6�y���W�,4��c@k�����` |��㶰<a��<��@�'��ПX���d�A/r9�tYtV�E������3� ��"��l��'D���y
&���?���L��v'�L���T���WkĔhas�L��x4=�{J�3^?�n���	�݌�t�1k��f����Ef������4-s�/S��ϖ�6B-�c �l��0^}z�j����l���^/��?ا��qx��'#ұ�</����(k��b&L�p����G$h�I��B�QE���ϚF�S&W�λ�����ml���I��� m�ɻ!��1�N���y���!�e�0�\4f�,'	~2KT�ǁĻ��f�����?��r�r����9K禽��۵1z�{E`�j@�9����E��S.A��;�e������'�����)&xR�$�*a�2i��&��3���/�E��-�K�~X�u�)����䰀��'�mi� *Y�R7?��/W3�^�����WH�t'Gx��f��ѯ��� �O����J��SX�2��#8k�Uz�c��+��m������[х�]�t+�_G�Vf��V����wN�Ka�~����&�:h�H����?�楾�9��R��L�������X�ӡ F�Tj�.CM��C�c{`���H��#}���q����1Jb���|{���+������^�g�S1�]��G#Z��3mLl^i�ö��=1�?����K�CYQ����cYZ��m����Tz�U6�B�"A�.���=�iG�J��S0c��H�E�t���J�!i�_�#�Oݠ���ڥ�ʊ>'u;�iG�t�T��Ti�T^|���F}_���e�� k�By��l���=�,��	���
9�$�G��A�w�8�g��X�[0�Ǿ�|+&P�r�}$O�vˉ������u�y��e�P��0�<K�j ��'p�m!�,FgloSG%�	��rd�@e�w�	�p��HL�kݙ:"�̞�.Ә���}��~���O����W@t�Ob7���W���Z m/Z0�o,]G>-�� <iun��x�N�Bc�̉���C2��VAz?]�P�A��M(�J�e|i�Gan�<*�J��)v$-�J%qԙ���Q�J�a|;s7�lqs�Q�Q���ˀ�U������?��V���\�ܲm�L�ȡ+H�G���
売yV�|0�_:���i}���:fҡZ��yݕ�p�Y 1�S��O��X.�*�����MYW�?��	��k$ �ӱ�T��㘟s�`���R����nE��W�(=f�2�O��Yҥ���D�rs���)tc�c(�k�>�'I"v[� "k�	�/&l�o��zs�Hq����cx�H)_���3�����¾&?�}�V��dG���@Y��Nq����\5��d|z��SL�q��+\�Ѣ�Pt}�ĩ6.]<|ac2�������I�T��j��p/�4$G9�mu�2hՕ�2)Dw9�u`���;@B��@�o���>��Sg8%�� Bq��'�8e)b8���h�C��%}9�;ö��ܘ�V>�)Uw�d�O`��s)���7�FC&B�c�8�x[��#��o-ʹ7��i������r`l����g��/���cj.Vr� ��Ϳ�M�$=7u?�w"�#��5�-�%�UY����:9�T�x�?�����_�Wj���N$
�f���<:�8 ����jG���fs�-��,���� 5"�a�Ve�и���bZI3��(���n�]?�h�\�.}�F����Έ~K��?�ܤ۵�]��4#<�+��3��^1Zod�dB:�mY*��� �1���uE6�6Ϩ��g�Q觇R�p�JH��&��T�v{�Uj��tC��^�(�Z�}k��j>�I���JY�[2i�^��^�����[T�UZ�^W���	LZ�br �>v�
S�ᘍ��e񮹝�n��Rn6%��B$\��_��i2<7�a�6e��*���w�"5Y �&+K��0�CZf$E�����}��v(��jS�kN�"��
̘G�7Oa�>oV�3�DQ$��Q�-c���ca�lk�����d�L#*�4ֻ�4ӧ���y@{(��O{E�z�$-��H� �����6At����B���:� ���<�K�x%�S%tW3�g'u���`�����~1��U�M݆r�<�.���H9�Ƹxr��29Ǎ�n�z��6q�R������LSzkԲ{+k��Q:h�XڧVK���9��Ӊ�,�Ћ�%]������C^xC��]H�r!����\��>y���B}~C�����$e����f7��ӟ��-���i3����@g`�Jl�P��m�q�Jvs3���׭1��x��Gw��Œ�&$	%��rN��� GN)O�i�����;.8-Mjh���k�LY�:' �>�vR���d(���Ƿ��jugdA�ecr��0Ίx�\���MU�<��Mzb�A�Za$�W��X+�*��#ҾI)�X�&�@MD	��*o:מ��w�$-?ډ��U���.��e&U���ws�1����<����u����j
yB'y��Fe�J3w�M�/�@璆4���n1����ys��v�} Y��ޕO��R<���5\p)/����V��G��"KKҤ[$��`��b,�a�];�(�qఏX�A����ef��u}��ǚ�d�%�Ct�o�cl���������0#��Z2��@eB<AeS��6NK;yW��l��i��@�#�ݺ�TdD�M�����E�R�`�׭9�i`��WU�R>�����I�ڱ�O�b��Y���u�P(E�T�@d���`|�0�X�ݟ`��w�������5��K��k4l���ٔ�>o�����������ӽ��:	�,��xZ�2������9��y���$��6>���	�5B�H���5�W�Lӛ�)�)� )	!�ϱ`��햋8�T'�Q�[
�h*5�"Bu�}���ם���K]��f�9�l_�u?����Ē�	� �R{��
�{�{Q`ոZk� ��=`G��3���� ���@�h��F<�,�QX�'k�����9�!���YrZ�N�5��b?��l��'P+!����R��0��97F'�VN\&��`$+��.�z�Wf-e'!�B�{X-���6d7�!
�!G�\��ǐ)"-�o�l�5؂z��I���>�xc;H2G� �nX>et����GL�1��9���w�����C3�VQn�����Az �𤓱R��p�"5ܳ�%ۥ�e�hF¦���C�0����p��t��q�)܊Y�t _�X��zK��p�0����k=�0�Y�Nu�x���p�|�,���_]��p��F;�~����\�~�9}C6+�ݣ�Ԭ�m�oS`$�/�e�%�=N����^D魅����$�g#P4�)��ዹ��Y_������E��R�4O�F;g�/[���d���'d��3S�O����L#�Y~�3�y"9���Yqb��cbj�6��%;��|I��$�L������n,|6���Dw�1��ItJ^�֕���e��?�w���
��hٖ�e�*�GTR�*gʹM�[�W�����/J��M�19`��v�+��MK��nC6$>��$n�<j��'�O�e�f3��� o��I�*�n�����z��:h�2?��~�Iw�p-/k�ˢ.��:�p���/;�!o&�?���=&�<�.wi�5��(#�)��YiB}I����$�F1�������T���*���S�%L1�x-٥��=���}KEv��}iڽ)l���%{��9MG�N��+�G��� �������[ZZx2
������,�
Q���ɦG!2eGP*�[T�cj�R�6Ĥ��kx�g��ϋP��=��9c���I��d��'��j2�X1I����rCO|J2^R4��08�l$�w�,���;�8T�v0��s�xB����/�l���e��ˢ�R�_��^/��h�acE�g��
(����G�l�"��']�[$,$=�+Ϋ��e@/�j�\z';#}c9u򌋆M���U���Z�Sڄc��_�nj�؜�$���#��͂�H 65J�V;���3.ވ���@Q��Y(�dx�O�"��f��~�b��'PAd��RB��J��L|�&'��N���vy�*��S�[�|�߽��Tl�����Gp�xQ&�6J# �9��\�ŧ>�!�v�����ܻ�v�z������H�*��;�T�X�P��Y�~Ԇ/4���%>�������"�d�;�E,�
�g���-�4�����W��mf��5g!6\��%���@��eRʯ޺_D�ˮ˲<�p�`���]'��H��^+KC����s��ɳV3�ng4����-S�yJ �-4$.���E���­�qOM��M7�L�	�Vh�i�@b�G��(���Q��}�����%�
���Ca0Y�T��T�+h�Y+���:�4���_i#����bI��0�F�D�C
[�w�#a��$\��%�C%�����MYLӷY�$�g}C�i�݊�݊�+�fS�F�D��O�`�G/�8���J���R��uj��_V	��VeB�a��Ŕ���b�I9߳��'��G굅���X���9 r�}L���7�YY8W8E��R�z�<���FӔ����~�W��w��[_+h�3*Q�F��E:&����G]W|N�~�o�ٝ���f��Y�"ic92���ߨ
B{K7�ǻ4�\>��/��nZ���l�W(trsc5U��LY�����U��`����"<��J�2@�A��)F�6���J����T%7.���ĳ�*_��唳�f��SNtk��/�"�xWz���K�/�ܿ2շ��1�r�׀���i��ի�5��7cQ_I��a�[EyJ����&��dm*°?�?�M���t=~�M���rS������:�:/�ٔN��ɸV��%�� ��Ys�faء�Y�X�d���`*o�O3�뵱B��c�C����aPU6�A^h�����4K�"k��X���Kr.��~t�nbs8E��Yt��U,��q�ކ�/s5=���V	����pxG�~vC��U&�_I�2�k�	��gq���Z�w����XV�-��j��pD���� h��dl��qa@*�������Y��A�΁2��򨷘�ʻr�1��︴�W�	GX}B�6�i�A�rL�x�j
i�����3�a-O�	���@��(R�� S�՚�ibU��`��r �����	�y��(js1bN��X�d�F����c]�Υ�D������DE��7E��Z>�-��l���x���f�'�d��=����ե20TpN�x���I�n�[���"��I��r�s�G�44J�ʂ�<�b\���&�5��76@���V���ȪZ�4j����\�p[h1PP�oj
�Z.|�bx��/�Xq�� ��`Kz������yj�I@�-Y���W�uց�=��	e~�T��̹'�O��%�"vT��� ��Ay�nM�	7��.��h�6���Ʃd�����:M��}�j	�ψ�5pj��C�Se^��	@^�k��=�z�k�q0��4��f���ɢBr�-@�x�P�X��z{�۞SZ"�<�`+IQ�;糰����*�T9�����B	ED9F�L�Ť~�|������-��[�6���V�[�8���@���-�k�������Hb4�3)�O�Ho��	�.���K��E���?)���!�!g~��ˬ㭏=#��G������]G�;����'o��8#'l��:�>_��u���}8l`��SC�x���EM˟�{���_�BD12$n�1# ��|����e�<��-��6(�j������N�iď9
5�����#�'������������b��W�@u�)�[��4�����1b�h2�w�y
����9ǘ���n��A?��P��v���`�p/l��0�*���&������!�^2c�5�&�$*x�� B��L�dzB���A(�
�fVMX9�+� }tS_l��N(bCP�=蹁�Tm���c��ɬE_L���trv�r��~j�2�eAنı�!�EȠ(��=�u�g���FQ
���G�SW�DM�f����)w��,�vɝb�@D��x:`����oA���f�f��}'6����4ȸs
�8������k
�uWQ�1�����S�2�&J�����ەA���qa3s��8�`%�i8��t�̖�ȿr�����t�`$��^;�i�Y%�z�*]$o���l�S������_ֳy����|NY��dk�ʳ/ML��uA�I��Q�b*�Ӏч_�O��Ա�G�0�um�����GƏL·v��g����	Q���D<�F)��GV��}��Pl�s���|�����if�������e.�� �jx���ǿ��$`��m�`J͇溝����[�$-���+�1�`o�k~-�:7�w�����4���6����K+���z1��W"m֝\#����C��~��5�(�W�x��>�bt�I���Z��v�P�}m@O0^ � ��3Y��-�ڊuԥ<(WC�I��_�
���̯�=�ZB��G{�c�y��<��e��X��Ӭ��1�%�Ũ��.OZ�6��`/г��$����S��$y;*�gD�p��i͵(���<�GӁ�Ȏ:�"�i�n�ԥ���e�� ��xΉB�s�B�[PG�)�>L�㧓�e""�k�؈�޾��5d'+�i~Բ!��4��)�@1���T���@&Z�@H���06/�A���S�HU(���QtA�Yb{�8$-���Wiz��WF�2���6)Y���=F�4����ٜU܆�&.�nU��3��Tu}��tm�*�H�fC �"Tl�@t��i3G�y�{�D�5ŏ:�ί�� �W�873{M,ǟ������wP�`P��oFd��s���d��
�P8�� !����
��U��ƺ�������M�;]���&����'?q;�1�Ƈ��W�z���x���]�EFj��Lj�Y��\�~�)��<�MT^��Da��E
PT�E�⫨#q��g��NBf���pa��,���I"�R2ٕZiX���� �v���������dI?�gvS��*(G�DP,�zt�>���U��YbW�,���c��'q�3B4�V��C�\�+�{��㌮Pyor|�R�	.��o�`Hc���Z�2�}��մ��ډ8
9��<]Z�v����+���P7�b���@����)�LtN?P0��b|xb�'6�����5�G�,2�SZbV����M�K�I�Pǅ�O����ò��Ք�5�$�� ��DCP���I���ļ��XK�<c���]�kl��~fu�|W+��jx㚻!�sA�/*9.�M���M�@8Q���̎��d	�g�b0��IyM����Aa9����rOEG��߈Z�"��E����?��e�)�1��j��#ds��ePYY�8سY�݁������OI�p���HDh]����Ad_4�c�i#��%�-d[8��c&����p��Zz@�dH��\��Fa�JW�r��	ũ�J�p	�K���UP�*/��f�E��$��'�>n�o�h��O�'��* ��m�ލ(��F�dlW8
�����E_�G�|	K���/�-�rPG��.��˦=\>���������TU����n�����?�WPa���E������]������r�a�R��U^�mLy)=��\S)��(O��gd箍�Ҹ�!.�w�sUY/�䏱	�"���T�Ъ�d��k:��s���!f�w�o����i����;^z�ʃ�MK�%Rׄ�!�/\�?^Q�F�9u��#<��6���u�ߎX�Ç,����_�qD��k�IcMAl�2d<�-3�����Q	��a_Hr8*;���'#����������Y�}�:MÞ9ϱ��+w�-P�\��+�E@x���WT�BU��1��D��2��M��!9����P�>�����S���x$�4����2�H��V�7Y`5�1IG���x��F蟬F��Us�Y���p�b:Z:��f(y�|��Lw�������ŋ�S9���t;Ƶ�Z
����iE�iL�5.����|�B^zXvM�g�N[�(���l�=i��j��Z�97W
�#1���=���H(��x$��&�P�4��ĕCծ�?P���W2�/;ᩳK0�ڥ`���`��T����yKU`�0Eb�7�W-CE��ܔ�AH�����'uk9�ppR[.o9Y]���(%���pAp�M�ݣ����� J6�n���D5� �d�9��5&������:]X?߱��cB�g�UwSW��K���zB3�ŠYY�K�}�0�$^2�1
��h�����"������<�P5��}h7������bw�>{T��ҳ����ꩰ�^�<>�{Mp�e���x�ϮpY��p�j��ԍ���#��]���Ǜ1h#��gO�LQl��i�e��#��ẰנI?���8�
m�C2a����Tޱ_�y�w�����ӷ0��!$��rNŊ�4�۲P@E;LC���XR����ˎ��},W���,��I_FT=rW����N�=n5þ��%��v�K<bT�Q�ª97�NB��@�����<����'Y��ӠiY�Б�&�( T�OIjp��V}�R��a�fw-'�9��c�:�vo�r��GyPZ�^��}١#�Y�6��$�	���/��(�w��c$�,U��ڰg۔�.+/S�h}P��ĲW ��I���e�YaBS(:�N��D#%3�����$�u���c�(��e��t�ڪ��B��v�(L⺅�Ӫ�@�۵C I�lFZH"I��\�"����W��JZ�N��JP�No�C6�}
ƞ9���9��H��g̗��w�
�t4���c�/:i��Kǈ�Vs]�M/�bEԩ� Z�2� ��(L�G�_i�#���-q��A6�aJNr��r�FR�B����b��?��m���,���<`���u{S����qElb�*q�r��
(�\`͖�c�ąGMy�!0lv��{��]��V'� �~[iY� �ҜP+L� ����� �-�z҄Y�T�xJ%���E�*lE�Bl���Z#�H,m�Ôɇ��>��|F�q(ڨU_�|Z��EU{%�T��͜&d"�̚=�*
8�u=8W��V�G~�EZEW��M�s4������R��9-�r'7�(+nL��֕��vz��6��j��G�4�&?�������l�;o�M7��:�l��#P<O�{7E�yݳe��<��oU`�C4Й=yŜ��v�8)����>����4��)6�դ�ޏ
��8̚��ߌ��eY�Z�
�}F�G;=���R�(�FF.$��>Pn�2�+m(���R­���X���?��m�Q�r[��+�3�EN�K�R���S�7~]�����~�:���@�7�= ���QA�Z�g�#֣܅Ao��~��������#��OI��k���;�C�w�)RC�1ʎ��5��L)�T�1L$p���6��*�s�ZMH��Z�~�E��7�M��ykB����rnﳳT�L��/}R)�(����v��V��4�\g�ܐY��1Ar��h�x3�������Ёh�� G8�T��t�@*`�:Y[�g<�q����S��e�#���#�_� ��,>RP�ZG�n�CTA�� k�{r�I����~)�AT|�4�� 3-N��JѺp�3D���0�Y�U������I�}�+��B�ߙu��N6������RTa�&�#�&#��Xk���� MQ!�'}y�(�Y��_'�d�Sh�p�'Z� �N�Bf�2�D��ȵ��S�\���"�ؕB�O#%p���Vߊ�tV��4KZ��]L�0N0I������P��Sb�+ȫ*%sR�����E�N�u�.^	Z,!�F6��$k}{(΁|�Ќs)p��D�h��\�H9�0�͹d��x��S�\��lӧߙǂn�CD��}]v���i�ۂ��b(G!�Af,�v�,�����W{Dޥ$�t�{�(���g�k�h>��(��������֎=mM1��qtcRYQh��Y���ݘ ?�wR�%�I2��AD0'���oЭ�}��2^��$���5Nf�8>�.�QҒS�}ŘE�r�NN䕩�ٙ$�֎����a��ݬ+t�#X��w�T�J#;�S��� vɩ��غ"�_�&�rn�A�J�я�KȈ��J�w��\rcLl�i�vu-�$U�PN�:`\���d�L�����=�D�F������,��'��!�mG*�f<Djb�D<�'��;����u�r!�;'1��� -ы>��s2��A�ab^ϝiR�,v���NϿlB��3ٷ!��z:Q4-~�cp,�;�Y��x�� h/��ӹ%s�b�p
%ft���;s���@2&�f��,�A������U�������R؁�܎���^o:��w�3���+2Ґ�ڪo�ҳ��9�(kB����g/��}�
%A�Q�ɲiV��½����_�K�[�P�N66\�^�p5��#����{�,n��F:����Y�[�^n�M��s8�A��ܽx���CԦ"�M��+��Y��.���κ�Ly�%d%���@��zx��O怸����v����mj�̲'��ԩEӏ-�X�6��pC�w����I��<|,CI�h׉,��"UEU�OF"�H�#�·�������������|yG&]�H������B�zA|�Z`%8@����q���V�]VqQ1��h�gU�γ\S}��$bw�Qr�����p!�@����F��8� ��u��+�������~bT�����UX�Yd��w����r����"d}H��J���)�ȏ��T��� ��ћZ$ϣ��^�3�J^�y/f��i&��9)�jz���N$5�p��`Y 3"�an,�ڼ[�����u�D��?=���������O@�yE���#K�> ��=$�$�q��b[��W��N�Ӿ��Ȗ��;`�Fpy�n�d`�OW���
(�1����/��#�~R�;��&Z�M`d�v��ǈ	yj��	����UB��zz�q:��x���J�᾿!8��� ^� r#��0��=R��ࣴf���Od�$�}�����X��O(�A���@o{[w �XP�@SayJJ�3v١��f���ɂB��	�s��]B%�ā�
r4�a�ܨ�y��L&���jNY&�n|5�жi������#s��o���t0ُ ��s���l�#Z߮�d�)�޳c*���i�$2='��bB�LK��7ңi�N�E�<:��s���o[
SK�P8����S�I���8�I�%�B��K|�Em3&PqT�h���yש�y�g�E}b(���=�U��G�fF#��P�qf`�|�����׽2�%9�٧Ap�#�H1�������)\=%�@T���)7�X_� ?�_�+g��+/���C��=�m�0�yDJn�e=�>.����A��B7��26�!�]p��TFFy��+���iv_{���9��76�ILċ��������f��X|Q)U��U�]�km��F	݉Kb����W#�.^ƨ�s:��O���<�R���U:8(~�+�m���;͑��gr�V�Ȗ��,�>U���ƍd��1#S��죃�.�!@�X��Q#W��쬑tOD�[�t��z��$�@�{�R,@�u��ΥD�k��QI4>���W��ߥ��`xY�i�LʵZ�Tc̭��P��5�g�!4$Àp�Kb�6��$��R�pp��p�T�_ �'<{ӄUg��|��(r٧'_s�s�A*ƚ��S�U�}|�;�PƂ0�G��9O��c��@K��/�h-%8t�e�O ׃��t�5��0G,Z�0I��d=~��\ݍ���d�,l��͒��������DǕ/��A�)L�g7A����L^r��U�*�X�"wB咾���z�S!n��&��)��g�8:q,{�)�,�K��J�7��qW�m2�CV�.��ޘ<6�=�l*�Ϊ�7+��p���*�FK�~�-�O�/��ؽbr��n�g�&#�<pWi�����kV	b���]Np��!J��Bhw�ty�
���X��`ݖk����ݫ�&l*Z�z��������p ���Џ)�D��~�g�]f���={�B�{r"���=8ybfڠS#��/ݣ��U�`��j6���Br�}3R���@.�1�ee��,��wfG������q�El�(��!ꦊ�,+�y3�C�_��X*�Ţ�D8�g�6��2��t\ ��ɩ:���a�2ao�n%4����a���J�Ƹ�NJ��d���#��ʩ@8�F�\d�; ��}em*ϋ�e'#u�r�p��܌q����@���x���!���c��Z�-�v��8ːz���;����gά�P����Ŏ���T<\?�Y'�ٔU�L�S�p�r�lG��f������7@F6>"�d*���f[�}�k�4|́G�^�)x'�l,���v(�jB~�ڴծ���s�N�ʶȶb�(���ձ�A<i��t6Tk����[e�HP��jp�a��^1��S3�zmE�~lK��3�w/�_147]��8��֯���ғ�̔c�zV?����ݷQ���	R�ę�z����.�7J�{9�K���e�3w�m�bLU�|�1ĭ�IKؓU�2���J�M��*8lh���9�AMY]V�ܽ��0�I|`��aް9*<�Ԯ r�Hi��|�9�6MD~T��e�f��pMW�w��\akE Y_F��כ2�A����gt +��>�^p%ѫ�!�W
ǚ���ֈ��c3$j�E�9��ͷ��/(�� 9���nųQʙ���|L ���f�8sVQ[�}#�[X��q#���H�2�D��L�ѣ���� ��Ƴ~�\^�+���~�H�^�'��j�ϟ��r�`TF!Q�	�ˇ�`��&���rl�>����|	_�Q䵐��&��_\�}ӌX0K]��2��e�+������*��h��3l�i�r�S`��֫�N�y�^��|/�q�,�������z��(��ӓ�V[���>
?�\{�N�0q��Aa�"J�:��.����RV��qț�Ħ�^�܌B߭����d8��θ�Se�>��Y�߈��4D[�u��y� nE,�a�Aմ�ɵ����;UB���*�Y��� �Z��#|s���%��&�ߢ�L��!:;J�`u��*v��G�):/�E~l-��-h�0�F�P]8$Q+���o���/�K��t���Z߃��������$��6��R�3�j�����a�@E^ ��)�`qEW}��}2���ʂ���$wi��0Nt ����5;:$�UGj�lz��b(���*���@�`'!�臮�G�����@6��F&�O���3���^lH-_��g��^_J� {�UϐM����D�ƅ�6�a�Y=.��-gK���p�b'�&[)u�֡nϯ��<r�Y��tVv��l��x�G|l<��r�^�S�h�J���>v�r��Ǭ�����N9�H����Ue���h�k<��р{�M����%�x]H s�~�۵4�]&I��<X_YI�w�� ��s�����.H>-e��v�-�����P��k����n�W?�e���(�fT˸4�f���c9��`���x2ވv�׷��} 3�c"Vh�T�{���$J �e-��H�n�,�b�����=���~r ��%݋���~�w�n���X?�P+x��K�	I�.��ծ9��l݇ަ��u�nx-�����#�x@Rrz{'�|Jv]��-�Wg��`o��'�Z8�k3(��_�/�x��娢�&��cjG��}����a��<�8Z�2��
��p�eç��=�M��q6���c�V��QV�z���n�y�@�������6�$%��s�+ɾnS�����W&�G6�_�^5W��>�Z����<�x��p�K��oc� �n��ޏ���g'�Dd8#��b�`(���Si,}CW�$^M��
A�Q�6!�P�km������5�ۻ��n-����	�e݌�Е+oPM�����(X/�q� T�u)�%�^�� X�ިU����T���0\���!<}��40���|z�� E*�n��K!�~{j��[�O��G%ؐ�K��������]��������wZ�P��L����7{�V��E���d��m��P��f'��6I�;��D��m�|��H��h��ԴP]|tR6���Z��,"����e��QtYOSx{��ɠꉚq[�֧p�jW�e����VmM�B����Z����C&8��;�ي����;�zFa�Nԑr���L�TB����	�`��&,Y{��G�r?�r���>�au�@S���� b}IW���2�E�9eT7Y\GK�aJ|1���2S"ʣ�$l.1���^����l`s�"o�|�\�E��d�+ ,��od5z�{�
?����.�S�:|�>^Z�Z�k�2�@(�YI%
�Y7�@)�Ej�d:�*[��&����S�y�������[0�Rv�N����寡`�UE���]oд/f���l�Ƨ2$*�n��~��sIsq�RB��,'�z`g�J�Oi���o�lA����gff/m������e����3`{P���uO!�X�Eeb���+�C�ǱBG��1�tW⸪I�r�_M������Q���6��$<A������KxaKV�����D_�T��@�� mS��JIwG*,���j�b��XK�o_�< w�y0����������x�:gI�%��M��n�`�q,�is*���+���f��d�*A�IG������j��AE�|��t�j�䞘zi�247輘C/�Q:�]L�rd�c{���ھ\`��<�O���fX���ث�R��=�K���뭝�a���ƹ���U�[D8�i�߄�v4�*�Q�l3ZôD�R�(�K�/\�{y������'��m��f�Xe�����4�f�k�x�6��(i$D^P�Ո����|G*K޿�s���M�#)�~��Z�ر���	
P�#���f55ҐV�T+C��m�WM�Rc����g�i�<r�c&� $�}o��xců�pë/W���0�Q���8�R�?�ԏs��o�x�5B��6\���ϴ>�,>Y�T�.�)C
�j��`Z�Ϲ��� ��d�'�CNkk�j�A���G��ɂ׆�B����;A�1�nj�a�5���l$n,�Ϟ�K��`w6���ՙG��`=����$�47��2�c�]~�1�� no/�$O�7��T�}��S\�J�J��{5������r��9Z���t���3k��+����	�ү��Zj1����E���t6�`����U:��)��;XW{N�BT`9���Ipɹ?�"�9��۩�I+[��f�
�_��U�S����ђ̂l�3p"/�O ��q��w����=��ޮ���C���d����Thz��5���N@i2j ��s"�m��AA���>�D��p�Ş�)1!�x:�H�hr��E�:�H�U:ߏk�H~�RX�V�n_�	�4�%�:���k���R����^��?@ZaJc�;aem���3b.9�
P$������5��V��R��]���6�l��js���ܑ&���2\ʞc}S>w�����[VO��k�D���6�Nw�hR�/���Z��g6x�rS͢�d�>Ep�@�0�I�0yo���o�@�2�*����N�d+�ř]�b�w1���d�/�F�Sog������/]��/���g�9������B�n�m�gq7��p)���8�η$Y?�߰��U:O���n�&^�ɗ�gaG�L�O�rE~�|�m)�Y��Xj�e�A�u{7��1��f�֣�"CU(�ߘ���@�$hyWj)i<���L���e�q��-��}pLY��vӈ3 N.�
��֚r(��h�B��K�+�$�>�|�٨��I�܏��p�lY.4K�4alȩ�It�C)��r7��#{�Bb�ڷދ����u��Ϡ}47����*Z��ښ������ ��o��������E���tZ� ��R8
N�7a��'�	�0�~b��«c_V_���3B
*ImH�CC"��s�ߛ���%Fl��N�^l xH�x���ޟ���x��IhH��
֤�D�}o7��
�7��\ K(����}ՇO��n�ց� �O
ur6V����S8Ԭ8o�Qq�⠥��rT�G�{/��wT����MpO0����C�����5�Je�-7J����h�w��fZ{a�9�^��Ds�/���Fr���6�,7l0���3���̹J�2'�z�u�]�sv���@��,F��k=��prȵ�ۖ�T��8�E��nA�p�V�NVt���������9��q�Q��0v3i:J�K��6�zS�tO��t��Z��:��c��qī���b��fF�%�@lxq�n�Q�"3q�O;������z����%�o�bImL��3�8�Փ�x�W����/��I�no�����/��gI�����mo6
�:U�L��P�B�5��*ٹ�}w����e{��(�v+a�z;��	n�#�|�iQtc�j�6���
��o���(�w�dgs�qP.���&w�4z��b�9�7�z���{}.N���r)+;T�T{������7����y>�[�ux����,9�G��m�ͅ㑯��F
Cy�Hfs�T�	��	o���k�������݁-&���~7�X��5���QywQ��^3���͹�K�:����a�p�S�̃�M�Q��Q��:��;�!���O�C���3k�&4n�Vkh��y^��ʞ�"Ki"�t@Yˮ(�MpN�fbHϸɝ�1��jFt,���Ż��0��	E�5)�)X�~..y�}�n��)��N[f/���V&�V��>^�~��D���B�[)
�D����K��T�Iޞ��ƕ�]Q(�,B��x���(4H�#�+lޘ�n�v�����EX'<��睗�n�|����9�A{��]I�����t2G>�s+4ݠ�= -�׳x�o8�o�ɭ#J7���Hv��#f����k*���Px@t�?�����Z�;�?�m�����2���Ǻ���*�T��$X�L���"ɩ��[�ܔ���2r����|��ȌG�ti��2޲Нaz��X����c��ʛ27M�ʕg{g.�g��a�6��@����p8hX~�/�|�U��_��� �.�͐b>�:�Nt@k�<=��
{��@�se��4�����;���B~c^��n4�ɐf2�˩�0�T��w����Q����O�̇���J7Ci&[�p(Z���s�%�Z�����F5D�|B�p}1^n=�k?݁}����Ƹ�J���x<m�,y~�C:�Zp����~~�^D!XP���d�9.?�+3ey*F'U����jQr<6�^X��Πi� ��h_G��8�=[��o}7�	�j^=��%c�k����e}�}e�
���/X�i�� �$���Γ.�J�uFni����3�%8�&��5Wzu䦽�uq�ޣ�ʰk�΅�>��O}��8�j��	�*s�l�2R(L\���;��-���
|��e�$���qT��BK>�i.o�wl�)�����.#+�7w�A����Ҿ1DE����&����v�͡�����[R�{͹��zo��S�g^��+�z8L���64	��fY���W�=�D�}�����t�|>��t���v�n��਄�.���?0�G+�3Xr$����9f�
��CLV���$"��ķ����w�O����6�e�d�L�Uo��|#���������pE��+_Ʃ�l�|T���?:�7�F����M����+xlIV�[�#���W�
©�G�c}��WC����M�
��.~ �p�j�#�B�چX���_�wg�4� �����b� ��s����*zz�<�H���-QU�?_��E��+|��C걖WT�4u�����i	�n�)���\�w�tE���;�4�2�xW�V�Ձ�)�y�C9��J��0�Øt��+2�9�S����p���m���S�8'�H8�F��뵵�����]D��
؝��a7EEJ�zk�9b�Edf�%ҷ��J�;$f�hZ���_���x���"+u>�O�QR�)<"�� 6����/J	_p�(�1��F&����bǛ	����'KK HFO:nԟ�oq;0|"���W��	-T�팄�je������o�� �o��za~�!��gvw�*���c�)��qj@,�W��`��|�G ����]��S1a�b��UJ/��'�0z�sx��U'���}�K6�;�lw�R!z��>X;D �_<N$em7+|��6:m;x
lMSB[�&mhTa�lGX�."Z-��*�e|x�E��t�6_�EX��k�R�/�Ł��ZZ�Kv�a���� �� �Ui��o��}GA��I%~�V���q&6�b�=Ypߏs������Ej�-uS�qa�#�8�W{F8\�եG-�.#�<��lЄ�����7u�}���n�ʧ3'���-_��)��ޠ'rp�ij��6����.�W?��_~����%��˱��Ih�v��k�ȼc�_?�c��O7v�A�����Xx��Z���ވgi�&SĿG�/u3������f�~szjd���Q3�О.�5�1ǬW��L����z�M��歚���ބ5j��v��F����p,(��<�G�$���;����~�O�n�@G%�iRJ&X�xj�D��DٳB�������b��ȵ?�]��*F��%ۮ~��l.�)e@�#Kq�$�$8f0�u"��!�U�
w��0h�0σ�ͱ�y�P��2�|X����Z�x��yēVG�C»f됊�LQL�#�ҢkX*a頶�Յgк,|��A��X�}�m\Q7�ۚ �T�z��Å㌮�l2�
j��U�i��ѣ���|~���L͛?�^+���D�Q%�@��{��HX�PD��z��.OA��V�0���A��맃������g��<E�j���Wu�^u��Sp�6��8H$23��F��N8RƸ�yt�?&�jׄ�q3�E����q��/G|�>� ��3�ԯ�����#��p��(�x.@a�P�`-�FFO��a�̖i�$3��D� _���k�3I]HX�Y>�V����2��?�ߝ+��l��9�<�hL?��[�֓�A�c�
n���~j;�aѼ)k�V��3r�Xj��I�6ơ�r�s[~l�Vg��7�!�������S���1��
S��Rj��H�@���Z;�ҙ �R��Д�`EQݝSLr���S�F�a���E��x���?���?�M�Bh����s5�N|_���Y�s��˝�ł%c�ڜG���?�jb��k�BI֢׺9��#E�J��d�����؜m��簜���	}��B߁t2"��i;���9֠��M��@�(^��~��|�OŨʌ �K�o���W��.w<��!�ZH\皬j�(�^�y�K���ED���
G�:�2��M�N__��S�"�9�����B�41F��H�h�!�-�*�|�p�����{Wo�,��b~�G .��]�r�N�jp#L��aPp��A�9�'�>9�7ŀ�8�J& �X��w�[�iA�׼RO7ŭ�2�4"q,}�c�םͅ)���K��U(1�5d��l�:�x�"��Lvbn�BU���܌_L�����9���J�v9�4�=FF��(��zd�Մ�ʰ�Vd����p�Ӓ�B �O9o�ƵϭV{������KP����j|nid]��U�_�d8�~��1m8�/m�ʀ<W恦}.XM~�����l"��dIP�U���>H�Xc�7{� I/XN��E�S� h�3�
N����dA����s�_I�l��Jq��U\�jv�W�Eg��y���I���B P���׫��g�D�6�&�T�n��b�����O�?��>�/7��Ǟ"S<�Mˀ>�4M�jRȎ����L�]Ki�Ә�P�(�c�)8G���n��\��ʤ8"��N�g����"����B{ң̩�Z����w?TyB>	��-�?qZ\SI�A�**�[6�͘�ˬ��ܑ�2��/�&�\`<�Ҩ7��q���,t�(��hs��؎���gΦ�[�&�K��1��7!D~��@�M��t+1?��=�=�,� �FX��\I*��l���
4$�d+u*�R�^8;��SQ�|%B�Z�;lb|#_�|���J\����N�C�S��(�v���2_�h$�:��� ?��U�`�Z�ᕈ�E=�G���鹫W��2|�bn�=2o���OT�<]���7�~�z�3�_���������E9��~*�oZmi��u��A@�,�������4�
�|J�o�^҈4�mp����'���0!�A�UI!�Le�&��ýAEg-à^p=�ꦜguU�T�E��ӈ�C��AuT�����p�]d���V�:N4�:s�?̤7�4w��e�O��-������n�4�K^������#71�t˗����������f��7  E��mMII�X��n��á1�7�N]�BYY��y��3�M�<�+��}��O=��;e��n�;��o5����~�5ml!I�w�OI-C�i�>��5��\z�#����^1K���
��T�_!���~�@�k`IWp#������v�P�+wb0jqRO�e"J.�ҵ�rh[!���L�4`��[W�� ��w��:�	Q�qK����B#]��7�Q�\"����.єM5�R��l�J`���	~3ij��f`�i69U���#��).%�"B3c�XXB��u�zq�]9�s���to�Bũ�'fHd��I#��F��k�ez���"�Iª��=�����w�`;	KI�l̑@瞕w*"6��Z�����R�>Z14�ui�_;-�����f�2�L�eK+��"~?�Zx�iv�sZ�s�"�H�)ƣ�b&ͧ���K[.h����%;���;�.&�M�[�	�Uo�mά��1Č���G$�J�B,�h�L+���3S��Z<��S���Y�C�5��$~��b��i���[>�k/�-�T�w$����^uR�sR�x��>]�E�y<f��������d�@3�~��t �-�5�L��׭:��_���e��+,l/��*���q�vv��,��C՟���p�s-@m!J�-vklי�S��g��1���u��@����x@��r������z���/o�V�As��
8o���R�n��Dt�=��a�U�����yi�N��{ğ��6��.�j��xg��	��ieRnwy̌����4Gq�:%L��9�QEPVzs��
������H���"lwǿ�Ä��Ԇ21�����C��;=��Щ���k�~�@I xsi�KXM��ʎ�[9�z�_��k��:q�>���� eG���Ip��Ͷf�,���ս�^hk̞�A d֤!�)]�T��%�c�:U�sk�&d\�yO�Ku3z9�/:�ꣵj�6}�B�1���H���Jc�� QU�#!΀����D�;���]�k25�/eU�*~e�\H���}����@���7a��f�,����+�H�uP��j��z�	���J㖝p#�%V�&�_'� 3+�m��B�Qg~R�BA��kjaС�� �"C4i3�V��{B��w���U���V�靖�G��,i\x/76�Y'$�N�'D2�>��B�A�ѭW,5,��)Q�4;q�VZ�Α<$G q� Zb����?J�׾��X�X�*>���w_e�	Q��r�<���Az�:ڜ���3/4�(�qcbs!{OX��U�����c,�&@K2���mԥu� �A}���E���fˉǻ�����C�A��������d2�!��m��j�`���=��<�1C�^/��`���7#�K>fp��[���F�Km4��ɵ�wI�B�8�?QrZ�����L��"���ot�E�l��?�5��j�r���R?mvŏ���.:�o-���p5a�2�mS���q��1m5�]���;�}�5�K��\�嚋�`X2�A�G����l��_�?����`�R��+*v�uT���,1I���=�����O���[\�Qs���h XOO�sP2yZ(�G�C`|P�g�������1�%,�w����6m�$�V�*M~�Wׅ��[�2:��O��D��C?�E���<2��U�{P�B��S�X�oT; K; 4x7��x�
�~gd=��nk['�^��P���.��4��<i��ؕ�6��4h�c!����'�GQ�n���Q}�僋}�ƌ8}X	Q�N�f�j��Xs���0�ؒe3�}禐�Ȃ�c�:�ߖ�Sn�-�	=�B}����/��v��]�M��u��)K���z/�_�E�n�n2V��|Ą��a�̟Y�w/���l�ݚI}( p����&�8�|}7���=74��*�)�#���'{z�G<\e펏�*^2O:�����.�!ZI��4�Or���ʼl�]���2�T%f���{�F� N���6��w���3�4�?�n������K��Jb7�s�ٮ����V?I���l�r\*kKv����
�о�ɟ��$�%�[ 6O
��7���lɤ�{h��� !��2aoĚ�U�$	1�}uZ��e����7zk��dE���:G���l�W����y�ө�w��[#��r+9}�)�;C��!�x�S�m��f6`C�Z�߹r����UK^
q�ʨU*;�q�Й)Y���(p�x�!8u��P;�������'�|Z˛���2�D�r�1pA<�#2wT���~bܷ�����1����Eǅ�����^sO�3��D��6Jd�*�n�� q�� R�>Ah}&��C��4�E��VQK���Du����B7�I��4xM�^�w���1p���Y#�Ê�������=Z2І֛gd,� ���
�y�ZUU��N[�XD�vN}�A�)�$��5:I����ǌ�n���V��Ԭس�I>�M�EgBH��F)����>�~�u^��\A� l�M�]_#3&9���R&J��j1rc��[(~�t�m�[��y�b�$�hǶ$v�؞:��I�����/�vB��ڝu`��f4��6�D�睟$�Z���D�a7F&��4	\���.�̵dq8�h�;|a��=%iQߞ����~M�a�d6�UY_U(��������(3�ٷ�-�C�8�������!��%�0�1��^0nQ0� ������ׄy�35��l��&������ۭ�Yߦ?'}<����L����>ùa:d ��%�9�������?v`�` �����
u��d�;aX;ь(�_��Q�U�v�ǧ��%���D.�Yל����+UYa}���������N��É�K�ʧdϡ��t������1�U�al��]�ѕ�u����&�&'.e�O��Q�
�{��u/���U��X2y|�|�|�	b[*�O��" ���Mq��¹���&H� ���QIoi��>�����	xd09^��"D��������n.81�>�y+��u��(���B�gZ����[�bX$oS�_r��޺ͅ&�|?,^�8+v��Ga��G<y��Imf 2��2uHV�'�_�cn����.	��.��x<���v�\ >�CB���{E�j�@���;����-� ((�@��ƀ��7�����s�t1��3��.��ۋ��;g}v����`2\�H/����Z��,�lh~����I���滿�b�;�#\�%i�D����G���
/����"��n�04هl/k�X��r�rK�����G��1e
����k�ش��$��2�^�T��j�t�H��|��}��OdS�z �A}WfL�[wtwf����Yr�FKq�b�L K�A-�*]� �H�F��E�;��UǗM'���sbr�\����=�wƘN��Q�\8zI��RP%ܔ�K��� ���QzU��jNO�b��r����7��YX�y��Љ��xw�jA@N��ZY������t+��U13A��Ύ>
I����j���_<��N����^H���r�]ԉ������\.;��A�d�gq�q����1t���� ��Rx�j%f;U�ۏ6��t���l�m�GF�i'�/���6M��h��s�T�X�@od.�M�=S\�����V6�O�]�ϛv�X�i���g֛5�<�ٺ�dh��t~K,��?���["M�ZnB�$��v*��$�v��I�qj�i_V�l��|ND�L����+��-r���x`f���%n���&�;�7�i�̆�� '׺s��%�'Yp��&l�]�Rh�&��lY��w��#y���F=8��,���}��P���J�ղʫ_5���^a�Ԡ1M�8��.�nE���X��,���`z��VI�����)�H�AK���vF�j���*fy��Z�R���)1��{:B�aP��ӬB�����W̕�N(%�J��.�O����gEH0Y��{-1���Yq.�?���6���d��0,��^����?��S����nn�!jDj���
	,��fE��'b�Y�5ڃ�7�I]Xo��my�����������)yiFkc��w3����"�s��4d�.I���<�J���L�s^�{�KC|&Y)�65�4�:R�L_�u"a ��C.G�@#h�򽀽B�I�����^�;�F���9,ĉ�Lb�R�y��&�3υ㫛O���=
,�i�Do��Y�0%�ڏH7��6�`,���w��3pǼ�4� $����^��w�rk0�� [�K��y��#E"w��}���pb���"iS^�0�BY�ĘtF��c�I�C�^r�u<}���]��3w"��#��̾f����Ð��`װJ���]�(�Ɠ��pb���a0
���������Y3����YJq)��F��)8X�_���6�Zq�~On�6��ŭn�L�>�[+�up"��/n��s4a2j�ܓ�9I�S�E�4-�"��}���ͥ}�U �Z�z�XuJ���c �����Y[s7$eY�4�S"�f#S�] v�P,�H�g���́aoz��	�����]���B�<�5@6 ٗ�6������s\@���y��0�X�?m�=���T���]I2'P(�9 n}!�>��B����FzA(`�f�j��ʎ�F�`�Le��?�<L�D;>�=�zW��to�Q�X�󶵢\/�����F��(�N$wnh>�+�.��_G:�D�r���L!ș��Wi���6G�Q˱��ٚ_n��Ȓ���~T=�]������0�砿v�e ���4:�Ǌ+	��y���#"�$E��@rk��FN3����}a����Ǉ��iK��,қ�D�ڏ��Q��까�}Ct�O3�j���p��j�̬��)1�l�����$=x�vXq����'D�����v$؜Wpxl���Q�7i�}� R�O��?<����&@g�.'1��O�� YwY�Pd�gC9�P`���=	ω��s	����~��� �.5Ɨ�|a��餶y0��5�n|�K_���O�20!���	���U��FA��A�O����kZ��YK��I��䢾�4���G�f�l�I��Ç8�=�Z����!T?x��$<� �Y���=)�>�ݓ�xR����pˀ���������x�mrS��Z�t8x�*����-v(��4������j��F�@oS��-7
d =��:1�ޞ˅J�G�ܥ�^=��{SĮLc�"X�%�yͪ����U�;9����?�:��C��x��+L�ܠ�\ �?��GK4e�a���������2e��6�rf�7K���ˠ��o�Z��%d�~�0%4�H1���@��=5��<�ح����V�c�S�y�A�&1���D1��]���R�����K(ߥ?b��R_1�2��}�����<󮥋��\T��LI��Lz7��f�'Z���#7f��}gC.�v8��lm����$ ����6tE׌D6ص�|��y)�Ӟ ���cX��v:	��s�ͫMP��� �8Q�
�_�2�C���N��E�veQ���ٶ���+A	�p�O`�Dڕ>m�mOy�@��#��U�`��B�� ;������J��Oz�wh��J�xa���?�P�Y�l��4)����-^1�Q�Z{I{���p�d��.ɿ���T���Vۀ�����`{�p�q&U��F�����<>��=�>j,�����&p�a+懠�� �>ѫ�����l������A:�e��\Z=�B`���4���A
��Vܕ���G� ]>"�V���{|-xo	/����'�K'��N���P�4��'4?h	�n�o�ي�x8T�ZY�b��ܤvS�b Ղe`�X���,@x�}3�]5��Uu���u�g����U�Q���[�#�m����S^�2�%1�{&v�c������	�ue����MصT�{�(��)�	�t$��1`�) ���W�ֹD������g��\�Hy��9>5�C7� 
��q&k4ƿ'J�^-�PVe|�动�ȟ�x ��huC.}�[�5pU��3�&�*��p%��,�Z����$�6)�r� ��cz[睴Rʝ�`A�&�G�)��g��^��o�b�W`�y��@"�0W��]��ZA����h$~LT�qt딉r�#��� d[������[��z:?�K`z��ֻ=�"7c����l�FZ#9��WK��]���W~�o�2k(���ˇ}��"L�5<���MF�$6z��e���:� �T'<�c0���,q(����8�j��[?���a]q]]�$�[A4�u9�' g=l�Gk�Ń"%����T ������T�������,$-̬x���t�����w2aP��<޽�\䐔�fp�O�t�*�;�h�����ڐ�~l�j��m#l c���@�PTn#��{�|��w�V�ۂ��&��o�����G��Q�7sם��'�Ԛ�oT�Z0�me��}��E�_���$x"*��R��_�XV�c&��ȳ�m�a�H�H�P���C<����ׂ�ؐ�ۿ`f	���tF���c��En�׎�@���%�{��%�o)�/&Pט�A�h���wh�g���tk5�[��C�u�gw�ѿ/�[��-����#:�֡�2D�<�ҋ�c����p�$-E�#Ea���I��L���k�}ڄa� K��H��[��Z9�9��Ѭ���Af�u�iîb��o�,7�\P� �_S�����,1����*�dM��)�����:�d9�9��/\5-UU��� �=e��,뢵���<r����z()����ɐ�y|����Ӌ�h��Ue����O�K�{Y�Un��_�d��,#�*�6�T|AI�p�\a���Z��y�hu���b^G�M-n渌G�ޤ�Ð���"x��arkY�%��$����?ϒ-E����F�B�9���i��?.�w(�#�ua�KÜ2��)`���m@�"^�2��A���L�8�?�_.���/��X�Zg#GW�tV��)���	9�N�5�-bl6|X[�$��g�+�wk�?c&�*e@.���5�jW-��C�%_��5�izE��Њx���<={p[��M�� EjV@r���lԑYv �I��e|�/t�Ead�`z@�# `���a|�-8]�>Xy.|7n��� }��R����~�i1��	�Fn���1���^1���_�}��2�=�d��^{���>�E}�$�#[����nRl�N��j:Q�}���'���|[�j@ޚ���q�Y$��4ފ���0+�pZB����$9�><ǃ���2(o�,��l'��p�5ͥ��ŋs�2��Ti^��1�kbYi��򊈷r������a;�Mn{^G��O�Y4C���Tf�Nl���ҷ D)П'��i|їp�����E��$I���fmFn�Rs�`�o�^BY*	,��_]+�u¼E��F�M=O�5)�[�����(��G-'�a���sXEߏ�5�1G�fy��l�?�@�0;��n6��6+��.�{��V>���'O��꽊[l�s�J.$\D鸖J�@����f�Q���-��9'�hñ�lA!j���J2xu
����Kxc���I�ԑ�]J����x�Z1��7Y��I{��f��F�xt�!�6�9��=���"A�^����k3AO&�X�WQj�Y7�~5��Sm	��=�>��v`K0��qF٫y�t�%���R����f�b9C�	�f���bW���xP^��H\�=uw���C�W�v�	f6&���5���#�� �������Bg��m���e�+����f��0<ĵ>����N���
��Eo@��&Oփ�࿾�Q�3�O�m-*g����<��ꋩ��:ЎX4�W<M����~�sjO�S�ԇ�<���ʥ�я{U٧�T�eO=��^m�`�.f��х̩8:�����Dm%����%�Iy����8�� ���\�����B	s����4��JӔ��fZ��c��v��|Q���i��Sܒ'�kW荂�%��X�6����&����'�����/��%`DN� �W,�M����Rai�z���sE�E'w�W��ʋ��5��=�o3}�kAZ:��N��B{���{9̺���(����!��jS���Q��^���Q��|�Cb�F� ����?�j����ElMI,�
�ш<�-؋?<�(<M��E�������_eXd$�V�؞��]�P�� K�\,��n+�:���W7�)�x��D��ĩ��)Y��/x�D^M�����"hy[\��SZG���V�V���)��뙭����e��KW� c胅���>��Wa�Id��J�\e,�!]��H0K_?��� �J��4}ކ�&V2L�)��E-<���|�(��æ�\��7*�'/w�����.����>�*��ey5���pr��~^���;�`��Ʌ	����?�i"�ѝW��s{�����Z��yLQ�gTOTYt���Y0~��@ٯ
	p3��d�Aἰ��t���(���:~�Ý[��eگ�>��=�	g�/B����j��Hީ����õ�^�����pJ�J'zz���Ʋ	�촱\*�[��m�;��س�e���-����J�)�z;�(Ǽv) hA� q06���Q����V�al�W����P>��^���~�=�Ӊh��!��.]���~lm����c�9�K�.):CH� �`<й��w3Uk%qw�AS={�t`����4�e֛�$������y�?������O�/�������z�	�kY~8+���ù�l|���O4'�Hs���N)1>[�����j�r;��b8O4O����9Y���p,�x��ٻyZ���7����~�Z�K�3:C��s]��"}2v����M�T�0ѿN�\��W��,S'���3�#���Sn����y�#�͡"�{l�V��c� ��q����0�P�6�?�=��I����yTU[5o��8n�Yo�a������l̓g~�L:!!���\*M�Qw[�g(�c���V�#Z+pܱ�	K�{�oM~��a�U�.��n;��uÄ�ј��W������1����(�wZy�k�:�E!�9ޱ0"�A(��HfwC�t8v_-�΢-Z�o\'�Q�I{�y9x��Qd[0+e�<����x�>%3*��U��(k׬uW���F��g}KQ�l���Z	)��J���LlL?J���{ߙ��J�۽-r���<�a]s���xC�NU���R�g �u ���R�*ʦ����2���W�pp�$�՝;6���/��o�'3��%!ԙ`�o�~�ݪ�hb����@)"F�ŉ4M��b�j]�rB���?)x%8?x�:	��gj����`�jK5�	څ�JP56�IS*��!���|��j�9��ݵ�h6g_셊qh9w/�o��B������ӓ2�y�zV�4{O���Cb�HJ�s%$D���!"��oP�>3��7d��0��Zv���xK��U8��=�1�8RwMWN�A�G��l�T��$Bf���. �4�ѽ�7f��o]HZ*�nM��{Ey���?1ǯ��V�N9/93�����?���P��~b�o
�I����ή����r��oNDF�k-���H����&�B�a�q�ڢ7ZE(� 0ۓ�PJ������mo�ն��9k��=�x���=H�}.��0�G��%?�9'
q�*��dreIY���$^s��Ty��j�߯bk�u�6eF�ƜL�ag��y����j�5 ����6e����=mH�{��>��8M|�=IPe�d�Gc��a� m諄=I��A�:�d_�nS�p\���j^+-HO��tR�o!5�".hm@װ�+g�M�V����Y�wv�~�O
��-������"��$;���qy\Q�'4�(e��M��+Y��j��-��r�!�@�P��w�	s�h."��ߜ����w��MuA�6�ʁ#���(���˴.��9�~��:6�j��o�І���+j}����'�Փɯb��7��*j��Ʀ;ZG�wf���O䍮:-��#;T����`~q�5�{�x����R���c͘Oh�Tz��{�ѝ��?ܼ[X~D�t���á�d`�q7��'��)�?���2����H����˕ �©j����|MԉHOY�uj|1H~~�����G���� �!S�m�w��e�!g�*/��a�b��(k��vC�h�㫈Fl���������ƶ�*賓�z���{Ս_vqR$�Vx[H�~��b��wS����1Y�S�)UH����gl75(�=)���~M(�KK:|�h#����qWf!�P;k����b 0��h��\���΂#�J�2󈩽q�1	����҄B����u�G/�����I�n��4���LY��P)\kZ��+�Γ@�TdW��$y�%���G}��\n
T�S����M5ᥥ� HZޑ�F����~�	c����+�F�;;'���d��W�Cs,�쐢r�O������e���<��!E-ܑ��s.��9��z��ep.\y�.3�2�-vV]4cp��	Z��pz~��Lf{Q�j ק�LD�J/d����_�����S���r�\z�*&,�=vQ �d#�C9*7)�M*kd�߆�uHAd����c�f��*��1��>Q�<kGƷ�����Z��tQ�����ӎ�v�P�q�Hk���|�s�aI�O�y��՟��q����������%XZ�RS%�B��������*Ck�++�ؐ�b k0f�Fq��4*C�=h�t�o�c
��{��3�)��ghj�J�
�IxZ�B�_��HlD���A�S�Jο��c=x�8���f7�-����7#*»��~���Qh���KP@���?�C1)J�Up�y��/��kx9Yǰp�J�~���R�k,�:�v��!�d���?Tf��2\a�C,+3ۢ'ܟ�?z�3@��b��er�]NQi�s�4�}����M+;>��v�զ7�_3�#�@I�I���h�[������&��&l���[�H3���i�Q;̯���1�w��=%��(���NE�_� r0��ψ2�ait��������������~V�����S��j9x���,��Bq<W�i,�]q��d�[K̶����8��.�O�=���1��27I��Cvn��k��_q��I6`;'��_�
q7�KES��<�t�c��Q�A1�o8�!yS@a�6WSD�6�^=
C���#pZ�uB���8+]
�N�6��FY�Wb?{"׀�w���]�u��������,���$oI�{��`F�t�/h.+�L=d�'i�� ��R>�2�+����E�@��p���}p��M�y��M��7r肸��>�WA$P��鸴��9"��x
&}�|f9E:�K�D݁�#oXg�+�')9��T�K���ׁ�)L��
ǃXX���TD��Όfɤ�$��.c�{���M+�@#�zN��Z>|}���L��⇤�t�gč��Gw�o9���%=/�E7m���h�����7�'�stv�Tjk�.8��Gd�J��q��p���If>���\��-Cv�n���.��u�ɡH��J�2�tKan���d����*:i�[T�I�L&�t�ի%K�����ʂF�3�0��>���>���T������?��n�lq\�eI����
���?$BeoZ5�Z�t�z��픺�y��O��@ݦx�Şvܼ�
U@����j���e�2��I�U��*u�%���Ol�E��v}�3�T�"��tb�/�l��v³X�*�l=U M���IkY�h!�z����E!{\��B� ��J6�we GQ����3x��󎖊����~@Q�q$�[?���Mp�D�:xi֊�Xsm@(� �lq��lx-7�7��&�"�*���X^s+�}��n��O���,�Z'�es�"�j�ؕ�R�LB������3��1�^��Vv�G_�]�g�v�$�M�],Łrb�����ׯ҂K5+�ن�C�##��0���-AIi�$�o_�ϙ|���Jw�������Ձ�\զX?��G�f����g���������[J��;;�Y��F9b��"��	����N��%u���AV�0�Mwp3�5;"�| 2���%���n��}�Y�	n�R����2�Zի��;��~���9��6 ?��@��U��ږ��v�ok��\kᜊv�{西*�^q�ý%�hj�{��Bg�2  �9�?g<R���[�71�c.���I�eT����}É��:��Q��,����J�ah���x-P��t��	�#�����-�mTG����)G�����Iy}�˄%�8�Ul��M��3�� ��D~ �?uA�V�-���'��M���
���B^�|J ��0�����e$�:ʹ�����)�⡤,{��7�0I����.�.\!��A�aj���)_�#)<&�:���`�wc7{ᯗ��v�xV����;)B<�@I����uk_�Pw`b�St����Ѐ�M_�\	��JWb/���$L2@^I�s���0�m:��n~�ꨩ�yNW.q��~v���i�?a|:�#�to���Gʭ?z�iuN�8^p�PV�4਱w<���#h�(�r�̥z�)�u�ĭ�D~��do΀�B�ջ�s�g�V�d�f񣎀:y�7�S�+`K�ȧ���8�-�Dڷ��#�������y�v݆�,q�c������N��6T¨'�ǧ^e*n�U�h̗֩�]�A�h�S���]�J���. %(b�_AUWI1m����n���L!�-E���2����2���ܨӪ�H�!�Ӄ�:~�)'�ؒCٛ{��F�.�U�^�*���7�GW�
�/���L��o��dlnd8�q�>9S��/i(\T��y�+���MD���$�^oRW�f�7�^Of���T[�5;��x���"^v�b����^��5Y�x+��r��"2�"�сp��rVG��>�Ħ����c��b���%��
��jn���c��|����U\�<GycԱ�  Q0�'���FFp>�ZY��G/Ɨ�ӃR�T���ҭ>�P��)�w]M�K'o~�s��S#V;�����_A��hћM�t ��Y��h�f"�~���yCp�e����]
���^ݒ�䃶�7��P�B��ۊi T	��=�,mvb}���ր��0ʸ�b{b)����̍�g�go{�V�1�L�)^v;DP���[�a�3�ؼ` Z���+ic"9jl��ܴ�EB��l�aN7�V`�:�GY4as�y�#��V���'s���p�o��I�34D�S���2+���uڅ�Wi����;�1YD���+��T�X��+�4yKގ8ٛ**��3�o)"`��td��68�@��/Mc�38e{i�yT� <2DZ��F�"��?�[��ֻ�~T�䏩��!-1���?*��"9�:�������T`hBz���駗]1�{�=�l�to��Q�i�0���z0ڍ;��"�[��O,����86��ѿ���S��*�x9�3RDSy�_'?�6>c��Eyř֖o񴛒>��}7�����1_�+9����6��t��0t6\L%���"��v?����hH�p�v�˛������9�Q�A���Y����Y�'ۉ0*�z�����V���Dް�h����c4��ZW5�ǰ��Kή�B��ʫ����<�n��Z_,���_�r⣖�c�ӏ	Y��@���M�j�4Q;*�D�b���D2�b`;�W�KX��_#�t�G=��4���G��컬[;�P7��q�ɭ���
�.}
3:7:8A��ܩF>]@��K(�oCJ{�����< '�(�5!@�'�<�g����>[��MN������ͨ�~Hx'��z�5�l�Vu�{'Y}��q�G0R��������A��߁�%<�}�1	����<�D�ZD�/���;}pα��s��pu�����qtVѫ�M$e���r&�?�ّ>L��
�gjj�	�c����Փ�?��3���V?U�>E\ۮX�&F\��f	�x>��L9�Y%���*��%llޯ8�$�$���"xB���f�q�sQ��ԗ�O�Ä!����<�{	x塹L�Wux�,��N�
ܕs����]�] �������Z��@�nA�1����l�m5*�i�M�9� �6�=q����}/ ����^����CKB���[����*�B"qA��'�2dc�:��@�gv�f��X'����3��JE�&��~���S��t�t�{`]�B�ݶ8�IN6�#���k�L`hQ�"IhXy�j�d(��h ix�J	�)��|x�=���3�*�i��@Z��m�G2�zkga1���A�����>Aŷ�n�\
�؋b���yɃ�(��
��"�U�\���R� H�l�j��ceu�0
�����4[�no=��`m���E����qO�^��*|rp[��f�(^�Z ٭�::��J ޚ����F�T�L踉���(?���G�Fdr}E����*%�AA����QD��5
W�H�}OqE+>gQ���̅93�KXu`c
ͺ�M�T-�����T|�����Ŋ+D
��L����}�~dD�N�����>�+	��#�wف[x:���Nh?ldOWƶ��7�G��fc��r M1����4f�2q�a��]�f �����%�o����uY3q�2��f�2_i,�k��NAy@��䥬��%�n�*��܇��x)0x�mӤ�����:QBL@;%��"�4�RܑK�h�V�OÝ����1X��T��Lj�����v��/6�q�oά�l�b۔ݰ���&���|I�Kd�}��MC�#$p�4��� ��C�'^ja!����
�!�x(��Tmظ�'V3���$�RO��t�TH���M.n�voQ���3?�e�=3w�[��ϲ����ﵴS�'I��.�T��y�d�/ �}oɯ�p9��o�Z�n��s@,d�"�@Т2e���G$(��)rŔ@�8�(H���e���9HuHZ�:�"���eD���3���	2ض�؀��4�y���͡���_��R��qռ>����|��˙�-�")Wf[b���[�_Q".�$y8l����W.8�_%�i�T����K��g��?{����R(=�Q�e�J�F0h��������k��L&8�2��=�W�R��nQ�Zp��4�Z���)��y N��; ��o�|����J�}��+��^�"���U��Ve��6��=���5�U���Yn�~2W3�O���� <Q�g)uEL[����K�B��|Ю+��|�FP�~��l��?�<��t(-熮�ˀL�F �c�� ��
TG���e�Mi�|΢��ZЦ��`�B�N[XaRDc��c�&,{���S��P�q�i�s� G�"���N����We��i���7�*t������Xз���m��#��u�W� V�&GҲ4�޻��!��?Z[{@`Ϲ�k���Q�
��Y?��9$?6�~���_�<7s��6����:�ϸ.W��1�cʜ���)���x��mJ��W�����+/����NKā�Kt�q*��SP�d������զ]�ؽ�g���=Ѐ��`ZG�=	I2ݷ�H~a���c������<��>�*�ix4�S��0Z�/H��'q��s��m�bb�wP�	a�,��ۻ�����_ʚoX-��m�Uj��_�kM���`t�CS�nl{�ߠ�j$�I_�v[�4�E�E�q�h/e�S}0i}r�
���<�s9z%�B��L�E��%��{h��+
� CpxxAA��|Qp'�x<��o�އZ$����z��c���l�u%r6E���gyz�W� |S�����/����׊=\��N}g� ��mb��jQT�>��6��bX�<ժ��e���?[�4o��n@:��a2m9��)�a�)XR f�b�+.��2��Q�� �������5@��.	
�q��+��M��_��٦,&�5tĨr�p�0�Q[�y�u2$���_�;��j�M� ��t"��ږҚj5�a�tɋ޹D!��Z	?��x�~�*`�O�gkb�6�L49wT�.�����M)��'��l]�a'�����Ɗ[��k&΂0����)�,�pN�Ty���)��U����Wꭘ���ي�\ax��Yl�wu�Iv����!!#��Ś�wC�����p����ڙ�kRP�*����t�4&�G@���k���4;p$�Nzv�J����5oZ����{t��oՊ�����N>@q8�Gw)���$�y���͒�J�D��1�?%Q�Uag�i��Q���~v�D����'�ȭnê�%bl�,�k�S���b��V��}�ߛp��6�������m��K*,�L~̟ ����4��N���S�.v�외��VF��3�~����:| �:���Sx����
ie��/~t槷^4�+"��)�����EW��_4
2�-L`��l�k0D#0	$Q�r�eq0�r+��XL��FY�)�jB�: `Sk���G+�P�E�#���+	�����v�T��['G��W.2�U�^o���S(a�"�� ����׋:�T5�n�E���_BM��4��{	�E�F;(����:��z��ncwNU����#��ľt��k�?غ���Q�P;�o2�c5�+tl$����j������Dc��~T�@"�5���*�ť>[m��-���{�V� 1�iX3���B�N�dPr�AJt��/�]���M� ���ʫm]SX.b �[k�-�=�VҟH�,��q��RG�'��}��xiA3I�7��oLC�K%�χd�~%�$NuR+�ŕ��@�,V\M��V��S�P�����b��*�W�L���W�{y�Hw�T�0CY~d��V�͏;U0�˷�">T��{�E�t�%������V? ı�0�I��*1D��s�$��1��ל�\�#M��^'E��-�?r�M�+��U'����ɰ��7��&e#'�p����U�F���TB/�1h�M�4 {�Dw�̂ϺD: 5/_��I�;�"�K��Q����1��:�X�E��r�Z�t�b^����g�;H�f�������`�r�&%B�mZb?d�|X�Ѵ�?1s�Ns�z>jJ��k��/��7�N���r��S�"���3a�q�����2��iI�8����Y��>.���;&����3?�ݬ%޶�GI?p[E�i:�I��|����[e���3�u`4�Ȏ��
��;x�Wy�����h�Z�BP��T�#�&�k
��/R�e%6Su�9.��S.#D�U4�:s"�xt�>���S�}S�i;�\J�C�<,y�i]n��A������0Ď��|[,�Ne5%�74�L��U�&wЋi��Zk!{�M�*-y�je	�|�����X��s��| ;�������EV�g� �n�¶�t˖ШKQP��M/Y��[ֶn5�\�ay��Q�LS�sl�=��Zn	(s���Y�r.���m�Z�[|&"����R�;l�����N��a�\=Z����\�	�A���z[�m��ˢ�ۏj8����ʠz�N��He�tEop�88Nr�V��'Jz��v�@�j:�~�~�Η8M<|�'���V��G&���	~}U���������A�N����e�歏�,�VuX
�D�-�W��Z�:^���.��[���w�zh�&e��+2�5_ߺ�L;f��UQ��K�l���k��.���y�������Hk��w܋s�(LG<i�$\�n;����{�Sn�X'Bj�OF(���j�a2��s�v��J��x�`6��
lqQ�j�v���FR��KpQ�q�#t��'����Lt��`4>��N�|�C���ʎ��`,�>"�Є�v�V�,�Y��+��Ք��<sZ"�+{'�O6щM���ބj��2Z,q�+�C�SN˺���o��d���((y�[�5-���*j�Al3p�^�=�ǓM�\�K��d����'����d=�Q�>���q��[�(+ə7V�����G���*� 1lxH)p���""�sE��\��n��� u��?��L��Q�-@��s��͜�hN= �DI-�}�(�}ƒ�b���T���6@��� �RW�*�Z�WE��X	�"�;v��x�-�H{�Y�K
��Xc��E��;
B��P��9"�C~&�Ѓ������m ǧ�.��J��g'�G�//�/�%ޥ��0�Gݡ�����88;/�^&kg	�iʦy��m���S��2���@�9��%m�YЅ�Z��_��#�j�����a�ɴj�>Et�_\�DJ��~�X+a_���y<T���'��4���kO��,.�o���
��t�)�Rܖ�l�.B'/S��A��������������O��w3�/�T�����_����q����Kb�j��!#�b�d�{����!1�y��@�%���mI�g�KtcՉmۙ޶gր�	��O�S	a4T#�j��_����YϷ�*��Bi�a���K�b �g��M�:k��>���� ����/<���!U������Y�8m�,Q�������C̸0W��lCE��j[ƚCCw�|�����0�It ��1q2:��݅dZ���5tS�'��7H�>�ߌ�P� ��b?R٠��E1Fꘖ����w��*�֬�Ƥc
ǌt��W��K���i�<.�Xͱ����8}qu| `� `(���s�i�s�%�F��$y�fb�*�(�|����;Ӛ-��`ŕ���L82l����'�1�����͐,��?L���L(5�X�GL�f�P�S���W�:��9!v������*�֙�T3U�6����-Y4��_1J� ��,��hdÄ����9ޙ�:�����N��0]�T�B��+�2���q6��bcPml&����綃q�'S�~��
y��t��Pc�fC��l�4�@�sV�7�B����a"�v�'0a�"��9�сqE���f��άa����"ra��8�l����#����S�mgz|���u�u([���$�oG�~���r^�����d�U"�+L�"n,D�n����_l�`�(7m�I*�z-�u?Ԁ��t!�ү��T�h�qVTA~���f	d/p_"�L��Ol �P$�6O��0�B���i@0Kp_ę��'j�>�t)n�Zz�Ci$��_ZDXJL�SXЕG�һt����)��)ly���9�M�b��Y˹�3(
x�F*�����|{�d3�����p�K�$Еe+*�cF�b��G$���sw�<�I���y�:�K�����74���%贶2��Y���2:�^�J�1��"���c����JQ�)BI�^��g2�a��Ll_�]#pk1S�
tF�d$P@�%�i�;i�#�'D5�I����2��.��������s!�����K��64����a�F2B��뫌�x���;�*�;0:�(9�e�V8%�xi�I�9�w�u�{�&Pň��|�_w.~�H�F޷��R5��7
I����|bp��/�V�IΎ���z�nM��������}��`���x��kv����y��
�?{V,�I��E*`�l�/ʅ"(��@���A�YxTQ�l����N���H;��wR�vj������ e����&bu�b;��<�Z悿.�(	7x�dEEe�?Q��"�wį��{�R��K'��">��{j�V�*%�&�3����xھ���M��=���j_���0/n��ւX,҆��h�^���?��Ւ�tk�p3SK,��n�~����7zEн���w�|r)�?�7��jA6�ap ��(�WW���i�"���E��TXh����_���ζG��_�U�H�63�6���Gk�]x�|O�f�qM���^X��Oj�q�:��&Ү���Yc���$"�I>�%J+FW;��ӏ�yY{�=Y�a1dUQi� ���Bq���؀o*z�o���]^Z�������׺P�-�^���M��2�A�e��*6ȶ����g���hvcP��͹w�7Q�
f,Ө0"��v=���^��(|l��ZoW�r�W��ff'�����:^�F��jK>e9�fFi@9x��>70g惝�J�"�<�'X�m�F6@9E룬�����X�������e�� ������#~e��c&3��1��l$��\�M��)i�G����>��B �Rw\|�����?�z7�����SzѴ�(y���ѳ��i	t��64��&�6H��B(����Ч`�� {�*e��|С�Dy~�R�E��X����3z-��Y�
S&�/��4��[�nv��[�Q�C@��c=�T�PKBEH%U6*O1rĥ	��7��!2u�[8�=�9����1RT%q:P{e���;���Y�� �;x����d�m�;3B-j�[��C����f�M=�la��!cٓ��s��1Xm"�F��(#�%�%���4Gb NW5����i�?3C�5}�`8�S��ȋ)��]L�7�?��z6�7'�ߋ+��=�6����� ��������dX��4�t�},o{v�$E�0\qݕ�����-ً�&(�N�����j��q�;8��V����j�jF(�rW=O������`����c��|�����H�����I�ulW։������`5���I�G�(����N=�&9C������Z!����Lo�X� �,�r��,���!pJ�.����xOOIO�7$*'����+��e����22B�W7��	6J������lf)�	Y�N�BM�dQ�̖'��HN�ntJ�U���Ru� ႓�����0=�#�r�Z_F"��Ck~�n��e�It���jU8�l���ar�F�52�If(��h�ѱ�f������.
��Z*O�JG�&�����Y�i2މ��@\B�z�2V��o��X�'�,3^a��{@�6�Mcز2�b��<�W�2Kg��������l(ƧFX����>�u{d�7֞�5%ڲI�7��@��p
i�/.����
.��u��\�����	k�\p;s��y/�O���?����?��K�1��GY��b8�z�>/��ګ:_G�T���F� /��{�j��L���`pW�閛!�_����M��-�X�S�� C"'��5m؁l�u\�li���'u{$��.�|Ǔ�v����J#?\����$�����4F�	村%�h���j@[�8З�E�o�`�Ҳ��"��"?s�]���?�t��ē#{+�_�=Cp>t�_w*�.����:�d�+�q�x�iP �uK�M�E!k�037ab[��E����i�w�	�{˱f��w�BZ�i�M��ӕ�s~u�;HUw�F�~���;ޓ?	ި�wD�9����>�a�RU����:1'$�����h�����Y֨� ���!�i�҈h��:�mÊΨ�`
�L�r�����iD���	@(�x�
��5��� �]��8:A "�$�'�s ��i䰶��ӏ;_�B���Iθ%�o�G�c�>�"���l��\Ӽ�ZVgmV���\Y	3\������yO��q>��,FS�]��
w�+�}*�]ޫ"��,(�ec��N,C䈲m
�O9b.��JS�\�	�Tp���!y��<:���V='�L�Դ1|��
<�$洬��e�#ɼJ�K�4��vƋ3�����$�yn.�q���FH,`:`���+�n���M����t�ނ����í�Eժ�I��CY���$44�<0ۉos�>kS֢��f>hD��0ܥ�`i���	BD#�o�&Dt�Q�S���y�Z���$�Jr(��x���i��
R� �3e��`O"�b�AkB��[����	��E-kQ�o�.�#u���+�~ڟ���"��v�<�n7$\b��?����]��R�W�H���Rc���
y�]a$ӹD:s5�����0�R��Uk�I;��!հ4�~�S~�;/�u����H��E�rsa_p�����,Iq��fE�B��?"��I8Ƶ�3��v�� �A-�m:�V�R��p�!쨷��Lt��`P) j���O������"_ ��P����!2>�O����ӈ��A*��c<d�~D }rU4��N{��̉�:^�Y�^tW�>I
��-w�X@��N�SVQ�M�g�t�;S�>�6JR�2R� Q:� =bn8�5��2]��D�SN���ʱ���.M{�-W�~�ȋ��B0c)w"��t7�M�=P�`�4�7��%SH̯�w�"!��� `�mk��	�p7���̴�@-dUן��gDg�,����Lynë>�! ��c3Ǵ�����#u���:�(�Ĭ.2���~Q�}�w-�,ɓ@���S�KgeP9tM�(�D�u��2XF��
|�k�I����4�ˌ�dΛH�	�1>8}"�]�I��I�̮z���P6���KU��-e�`;�{O�r��28�j���ޟp�4k�U�2$��
.�>��&'�@Օ��?)e��_��5�-A':fNV�"���<w��=m�w��Յh������� �GՇ}?�oK5�����-�N��l��!�	2œ�"T���p��.d�V
6�.S}+��=kH�	~��Ж����� ���fr�fN�K�蕸��ȢIX�4��.v�L�M�E��ʌ�ۃ����,�����&-9Z.q1@d�P��aq�qbΞ��RψSV� D n��<7��*e�\#��<������$�!S�'��b2�_�>t]/��S���ٟc4^c�����dm['%����,�g+fO]"��x� o�ˠ����5����0RⲶ��	��͠_ �D#� T��y3G""��g1f*d�}f���jf<�����
�˯��$ʠ���jw�W�N�$�ׯ
~���څI�9A��3�_Gٟ�7��'�����/�y�bs*[6�ApB�0�1"�.5&�����@/��s1��]�U�[9VM)�i�K���Al�vt���"2L���t摗����Dʯv�O�E����1[z곳����8`ڡ�0Lu3<�����>��2�~��T�����R�k*7��բT� [ׅh����l���4^�%�Ec��
�{�uY<9���u�;�;bJ[>~����=��8n�g�d$��ꑔ�Ca�}�і�#��i���[Tc��+��C�I�R��<����}��%��b�tP0�.����nc-~e�b�)I�t|��p�2�~^s��y�Ȋ��(��0߲������ �jXt��i=Qͧ���S�}�j��0��!dw�A���,��W*�<�x~�t��F<��>Guͼx���v�JQ s��\���g��5�ڟ6�p#ߔ�(�+�ګf�K����@�����\�^}���$H�#�)�e+8w�-X��:.$�w�G��2�Q�y�!�9��D�<�ڙ�X�;(�]/ɯX�?�`�O6��s���7
�%7�V:~2)�u�=�􁽗��T�Xw�cy�!��pH�s�#��h���!b����?�'��J��xw|�e��P7����>�d��47�÷�Jצ0�E�xa�yur\�;�+-�+.�QC�Z7 B��������sP������l��\��Q:�4rW�|�[ �Qo8B�`�r�1',n�&[���
 ѥ�u��6���]I}-ͩ� �2���7��N���=9t��vkT�]h\�������R��߄w�9=��1(g��Ge��,>�q��_SFJK�s���+�p�T�u�jR�WH���x��)��7N�T�C+ �p`���x�����]�:%Z鳸�&$��Bj^��O˶�_iX`�6P&��?ɯ���������
b��$��G�[���A|�!5��6?�8�'lb����Ӥ�gA�����Q�t�#�D>'��bˠO+��2��{犟!@���@μ���|����x�3@t�MKNB�R�˕uT�MS��G�P��rP-��$����Ƴ�^�unV��׽����GM�o7E��ԴPN0a~���#�6T��Ԥ�����}�Ե�zN^�3��G4�O^)gS�AWm`�H���,�g�s1wpE�e7쥪�$�E��m���7��!�*�:�������Y6z$����U�^�x
�u�cn��;�i��5���pn����H-[���|��Y��2m`L#9��V��ڈ�WCu_t<�k<�4�_�!�r���~ߺO���%(GQO�k��ME�f.7�{i5��ccd��qJ���h��̋Ǆq�, ���������9���h����0݌(�.�1��G%]�R�)�T��c6�ƌ��璏s�W~���1��&I�޳uQ��������ufrZgޘ}P}�����>%>�4J�a��O��+��p�tg�D����Ə���^�8x�FA	B���L*qX����GQ�.$����6�����#����ѦsI�+2]Q�/Գ9�G+�������lfy��_�*#���f ��ћ�O8��d/�D�|1�\�FO�p�"��q1 ��N����p�%i�}3	,���F�����4�Ngl{�/KN��7Mݦ��W�F���_>����i��9�����jM���ZD�g=�[���1��:�0ꁤ~�W7���gٺ@��1��S�f��ș� s��Ƞ�9��o\2���z�y��{_�kHR��v��ۖz��}:V�hؐڍ~פY�+_
hR62*g��Q��;+6H��HZ�	�x�ȡ��<�FY�I⠠Nowp�y��_K-D��e�꣨3DF8�5m�p��`	��G! lV�੏�J%|����=ZLs��])�*HIU�<�D�|ZX]X7i�m��	����D볙'��nO3²��	gjw�=S&n���#&ͿD�r��M���f���'����Gˍh�l�
��b>��3�B��v�q"@�[(�.D����RT��Vp����s�k�'�PF֟��,��9�����a��"ܹ'��涜��ݕ��0ƾ�6|T	�"#
W�UB�����,�ב� .�Gc��"�W ��OS�y�X�ټa �I�I˄T �m8;e+�����'ÎiWBg�n�!K�|�V�m�2��̥6U:�_�������~(�:S�x~o}�o�H������AXHF��9W/4���U�Z�c���R։=0Ac��(���CZｊ𕸐g8�ջD�y��7%�U����o����<�R�Ѥ���'O�^P���2���m �N��f�T�E����ňI��n �Ҷ����&mF��d��8�_�-NRZC��aMd~-���
۰�is��橹ֽH�1]G:xS������{�_�*p�{n�nw� 0�h�>J�M�X�ڃ�!Y�.�b�EӀٺ�Cי��vOHZJ��_�-��9��S`�������x-�9[�"��+!���}��j�W�xm�!��?�����Xx��AzB���:���@Vi�¢9ל�l�A
wD
q�4>�~�'�������qP�Om�)IӮ����ʦ�}�"#*Uq�N��J�HP��~�|����Rk�TG�C�W�Tn��RY�0��f�%s��^(������}��\&����a��� �`�6ޱV4W�h�#h�n�+���`� ��� u�El���U~Y����q�����~���f \���3�unUf�K���pxh�=i�5xq/Lp)��;�.Fy�B���H8�L�S���!��@�<�ݖUG̓۟9QJqЕc>��W�^6/��X�|2Ps�ٱЯC'6��� Ē�`�4(����y#�a�2p�~_0��>YNpM��_�N���!@���A�陯�ܿc��I��ri{��.��1p��3��4��5\�7��%91�L�9����C����
���\��r}}�g���vIݞ���I#�*��U���7Y�����Ҙ(�����&7��f�,��?�Mݣ�o����Y*(Eħ�����"�\N���~���ȓ��,��*�yƷ�<�ǛN���1���s����3�d1����*0cߤ��SD�Ov�9-|�]�ȎG�EB�aMY�ÌEV�U �����"�:n0f�)���C.w�\�=�෧��?	�X-����M��fnSx&{���uc}B1��BcN�(T�z�k(>l���+뿳|g��y-枧�W�7�κi5q�+���e� ��/SD1��� �f��cq5`����}��=�]r��QH�a"��Q�6F���3t��VF���p��hL�K+�>��l�Y��%,�`1�-��h���Q�*gRZ���¹��6��
����ɦ��G'	�����Q�|��A]��d��8�C�%�KQmT�����-&@���&ؠ�!ž\ͧo�d~뼉��_�*QL���io�>z�x��L�1B��Kv]��d2~KI����_���!iY��rz)K9����~o���G+�\Eշ�ط��P�$�����S��hp��3�<��G����� zGt�IU���JHE��w�.2�;�5 �>T2�yJbZRQ�0�g^G�$�<�oj�v�QC��֯�?�*��@�6��h��uo�����bf�d�g��3|y�p�$i��P'Ci��'�zk��˅�O?�Aq"~�Tp��[�<ɲ�$����p|������4��A �s�>�R�����Q �7�]��rG�]4Ï{��}�MMz� sM�W]u�y���i���'d�E��qoA&�����=wbN�K��K�%�@���2r�u��u�@��@�;F����K�rW�1����U�x���;{��5M-�Ԛ�쪩��4j���A�WM�-����n$�M,�+N��T���F5ˋ��PՑds�j�K$���G��u�d�+x.O�H��������M��RfJ���{��E}2(ղen���5籀���L`��&=���᱁h6���ü��Ć/[�J֝S]	��qg)17y�7�\���b��Y0r��a�-������l����7*g�e�yO#�Ql槔�"�@`-����A6�[!?C���M��(�S��zx�����Y�y���� 	'l���Kc9�n��*�ưt���-4�����D���RD�h�)׺Z���u4x�h? ��c�db&�3��	��eN�Z�ﬡ�405�5��;��Yb�6�9��\�KD8!n�?;Ϙ���G��(��x~�G�	�DsR��o��k�	$���^`dή|��*2��P�����T(id�"(QI����z��C��YX��5lj�?ַ��e�����=�u(�z��x����P��O�ڨ���Ϛ�fH�N[n!�7�̭2Q(��,A�H��KÌ��Cc����I���E'��A�(��<��7��
#�bH����vA��dʩ���ɯ�5}����zC�II=�!�[��"�u�o~�%�%q`���������;Ӕ����,���-"<�I� A��w��?J��T�w�w�}����-�k;&Mi Փfr�3�9�X�稿��[��\�A�#?�+;��ث|���JO��=S���I=�(#>���lh��E���dY�0��GhBI7t�8=��0�i씣�:����q�d��/Rm�_mN{9^��SD�t���Dņ7�C������J$��\<���2�Z_�況t��fBj=����+��Plk^��/��r�~&��w��(bD�,�`8�)0d�s)��"������؁d��UN�*��0�Y�J)Y�Ì��_��h�[{O�h!(���mږ�pa_?��s�ļ�jR��'%�aN��Bɧ��������p;�9��vx�)��މ)' w��
�=	���n��4O�:ڮ���^x,��Af;&�$��5R�%�1�?�s(i��
˭������7��}^��1'C���E�a�H�R�QK�p�B�Y-^9\it�q?)頠��=Q��7��Jb���x�8��-A�����+��u��$�R��~�mJ�h���z� WRz�H9Рo�Z#5Q)��g��$���Ec�;�꺆�P�L�X�xꗣ���������¶�MJ���C����,�����x���R��B��X��uZP��ei9�2oD?�y�ɸ�}��`�HV�w�	��������}=��tʞ�nde��7+���ܦ���8C��ET�;M�s���-%kI��0�0Sk�*�� w7.Kz�L7��@Bf�qznՄq�ږU�(�~���놲�[�ǅh�f{��I��ƫ�;~���Na�����&$;ŹD�'�5D������i_��.{�[�F�_f����~�Q�G����ً�kú_"6Q���Gk[A����N7�L	�S�pv���P?&���rj�ُ�z��S�6�w�Q�0�Fc+��  V��{w���m@[nT���MKY� cVNK{�{؟ceb�KQj/դ)L��|�"�x�ˍl*� N7͓�]�%��&�F�dM�|���YS��ܑ(�l�Y��������z�1��޴�����$26�F֓��	>;%!{��|��Ɵav(Z�U:^l���<�W�)z�"7�H�����!�h##AL�W��V�M�M����%���@V�3"�F�vt۔_���<X�����	�����+hܮv��p��:�O��<	�)NhG�d��[�@�)[���4X��i$!�;��I��d�My��\�ḭ�\����`=�T}Yu�~	M`ɤk;<M����m�c�a��x�o+Bķ<R���&X&0�Qt��,o�צ�&ث�)4^�v p/����rl�&��lB�3�����S�9.���<!
yZ;��]��-w��L�����<;{Z���(�`���j�;��|��ź���=W�^L�\� #q �7�1\��$-k��R�IسC`;OI7\���N��{;�<�&��W��WL:|�9頎"���S�^��>���}�t�3�y	dZ���dfg�E����V-�t���t�2�E/`�m�1�r䌧�s�8'��D��.J+�-4�b֤*�2F���3�8 �ݟ�~��95��
����:���*T�x�.P�eCd�}}iM�Õ�z�\��AAa�p�:9ӽ�%wx��3q����C9`-#��\��Qv*��+!݊��Wsb�0C��iʧC�줃Xȭ��v��Ϫ�J�窽܂@UlmJiH>�y|�>�?��=�3ņ9;x{k��ߊ{7�;MoN�� c�c��2?��S¬�fԔ`�OB�� �yW�\s�͈�M�=�%2�������pls	�Fݹ�/�m	ڔ�]�w���]� ���ڭ��lTD�����mc�M���*�����l�rf����G0I�1ty�������\��'ǑZ/������^�SE{Q_��M��і�`]4��@Q�
�ő�
͜y(�]�"����m�)
��֊c��R��[@�4=�Y�+�#���Scpq�|��n�?�2���I��(m�D�>O��:a�>��G4J��Qv�hC�ı�M�[vt�d��*n/���7���.d��oj���� RO�QΈ*>��2��`޹"��C����}O�Q�=����9�!bn A��%
ɷ���* ~�р2�ٟ�R���}����:��Q4�\1���)����M�-Y����+��lZչ���"��e�)������'0ֿ�_6����kԶ	Z�m�y�������Q�FD�d�� *��v�b��"����� F����I�o�C�����^�jKc:��#x�� c$k�G�	$fϲ�T����|�BdJ��o���[��h�`�Vmh�
���z�'��g� ���~�C�P㨹���?��a�I����\#���ʽ�8ߜ�Cf���aU�!� ��J;��Ȉ���<��4?�Fyr@���S~_�o>�{?�1!�	�з�Ι2�ٖ�^G[k"�E�IB�7��r��^~6�
�+Ű���'�m�9MY�N��R�b7���F�[2fo��Zj��)C��
��C��2��&�q��U��kZ�(`8�G
A�*0e�P�
�>�JU�Ov�gK�7py��>�[���h�>~��U���r|�ݣj7�e��1M�ⷪ�[�8���TC�f�]{C��a�ԇyۇ��8������⟃�
�c_ϼP�PE���4E0{[]53Ml�'�ϼ�'vű#l\�P���СN�澶<p�%���/�orߜ��?����Eq���Bb�~ԛ��ƻTX2i��
��#�Y3�u�� �.��KM�����[�#i�x��{��rs��;�B����U�ʻ�Qƾ�|\�c������:�* �Cef�}��e�*�'gy�=E.�HM,/��k�K��g���� ��W��F�_�Q��4H�w,�F���BcfI�C�-���J�;z���p��K������bA?]���h���&�����J����?����t�7��yks>!CM}?݄��ȯ�k�5!J���H�Xc�a�T��������7�l���r/���i9s3��#Z��s[#�l�:t��ۻ��mi�XPI�œ/�6�dK����zc�i~gWc�����^��\��t���J�Y���6=�9�M�ѷM�,���Ap2F��^��G岞��Si�kAQW��6�8�ˈSi�I��:9�N"�?��{�U �?V�ܢF���H3K���Ŷ/
�+m�wj���&M��<p�/9�Û:�&��:�(��s�u �L�����=�)�d���
G��c�Xi��ZU���P��zYk��
����Gț��p�G���@��[������s���=��1@$����$N.c;��X1��c�H�{��r�O��<(�Y��u���"�����5�ͳ:;�鳅l�SC��ҩ]_�����Pq�P�J��[�S���n;���G��=�Ą���*�jY�A���������kP�)P�*z���5X�2#����)���/�po21Pз�fx)�������~�����%��ӭY���	m,�����فBڋ{Vnb!=RQ�8�Ľo�=��ny�=a����ʜ�C��*"�3���x�X39�^r2j�+����y��R=3\��;)�l��p����޻p������P���Q�������x�L�3�Ͽ'i{I�'!%��y�-d�%_��T�&�Х�$��+jYsb���RWPS�R���;�wM��y�e˄�^�j���,0��d�q�c�~%�p�Ctg�.9�S$w�x�`
��МX!o�
��g(�\r	A<�zX�4HB��E�h6mE @8�
P+C����'�v00�i<��箿3}�ɨLXK�&����h'�3�bg��.�Ϫݗ'?,f����m�|9���V=��{�0�!]���'����x(1T����6���B�:�C�-o���מƔ�мV��x�����J����S���JC��-f��U�6��Ƥ�s������眻A�l�=3�n�MQ݃�4_Y���U��SC��	��~�8�]�<P&����f�-�]�;=��1���Ѩ�tG�ا!Y%&��P�Q '�{��K(���h�AuЬ��h�����y��%��|I�������V��/�`�9��k^�d��n�IWv���	J�3:��h�N���}HV�I�G,;(�zb�1���G4���.��;��>d��hQ�6M ���gr��~dPn���h�Z�b���i��~*\�EĖ`���r������G�|�0�+ 1�.���,�{b�~-a���ݲ���~Jȇ맲YF	QO�o3�'2a�%ş.��L�)�g��w q/+�Ic;��~KP�!��o#��)�v`7�����@�߾X�v^�j�>(?�.Ǡ� ~q]&�~�v'�yf_:|<ĤW�����%��®҄њ��1���]C}���)�C<�'5���Xޢ�[q��F'v��KC��F��e��|������Qh�)	Ѩk�F��}8�����An%Kr��6]��q0@h�U����n��Җ�-ر�H�F��g�ǵ�eA|�E��F���ވ--��a;=�t^1�P�HF�����#V�W������^��貒;%��\���t��ˍ ��?��՜�/wfS�+��e�
F�� =HH^�:����,��y�C�7zOX������h�J��{@[�;[��.V�cX�1�>���
����I"���J�*w��NW�z,l������+knR���N�ۗ�t��s!��?|��xQ�)1��<E#�+N�ъx�z�,�O��zU0�D~�$��.q�C����ʓ�QG	��§]W�N��5����R�~߶I��"s�+�,o��W���ೆ�#�#B��P��|�&�||�Uo!f�r�;����3�Y�Mr���g��\���f���{Z&� �c��T��<��/���
���%�>j~b�b���Xߛ}f��[\>M�T�QI���:ɓ���ЬR�Y^q����L��]�B�fDJ�)�τd��+�n�7h���>ΦD�y{#ryJ
�*��� ����L��ӆ�V}=�l�x�����.|�|��H<�KQqP{�s�tW��Ir[��3�H#�hp$����h`25=�ٶ眣L��U_ps�
@G\��`�1�HF�P!�aizM�xA��$��N���9"�
	%b k�B��?����� b������;���z�����^�����HՈ�1��Q���Å��J��vK�'�q�O���O�bA��ڝ��9ٽI���o>�?ɑ���uà�?�=�6n1�!q�<BG�o`3NL�M��ؾ@����؈�ԍvHq��%B�^0�-���b�X�Ӗ>O&k��#wU����r[ ��#��T���.V^k�Hi)y{��S�i.<M�l�(���PA�?=�b�����@93w���kV0-'�t��D�ĖT@�����-|)9���0� �M1�:L1h�V�[��I�~J�L*/	���$Km�?lN��5������\1�v�},�g�T������?��G�yë����Ƚ����)w�'¾el��)�ͷ\5�] �z����/��C��?2A�M��f�?�2wm�p����X�qջ����J_"aQ����6�R��W��B�dԈ7Ct�t��:��Z�"���(2sHU��#�����`�u�eT�P�m�dk<��hh343ZO��J����.������'U����Z�o⒦pl�A7
yS��g斦��\O�d �*/�a����LgG"�- ������U�*�`�#�~^����Ba�ė�7y�8B���Th��zIz̻*��Gˏ/[-9מ�pl�@̻�����^}Qf���8����B@Uh��@�>�S�28���i�p$�iF�M�u�m�q����/m��[�ܔ��7��*����
�`u�+��C_��/�a�������&$x���V���� ��G�i�N��� �4$��1�v^��|�����X��jC6�IT�4��\}�)l��[�pkZ�p���̦w(3�ֶ������^��&�}P��ѣ�jp�����q<��hm�[_o�3���E�:�)����v����qs�{H��,�$6JG�_�y46^��&�[��=Po:>��m��}'�v7�S��7�" �Ɲ?���}e��,Ijfk����a���&4k۸r��h���&���P�a��#X�O��>���Iw����K�â&EF~f���00��t�f�="2��@G���ؑ>���&)�@�C�]���mt��8�q���c�������Z��[�a�E�w�R��exl���Aтmv�*�p�d;a��R�jV�V��^���hΘD��7Vfqxɷ:�FW�@zU�d�Xqo�f`�s��$Q?��qp}ba6Z��k�}~CB�Ə�?gĎg��>l�B�l'��(�r�T��CE��
=�4����&��Ka�0��*h+K���@��8����~�\�4��R� �/���!����H6≲��$U+�����/��|Hz�(�U�!K<f�4������*������ĭ��,A�做י|�w)$�Hme�X.��Y$�d�>5���gE��q��������mE�	�TU��|*'����A�p��$�xI�����P�K,Y�=�	��%�m���#��#Wc9&��\�=(�8�c�D\gx��b��əkG�ǧ��U�����]�����[����~d�N�ܿ�j��<�5Dϔ=2[B�� x{��Y�K�\a7 ,NrR���[jۡi0�?`#���N�"HB�ˌG'����"�"PA���?v��<K����ׯV-+}<��B!o|�\p���W�(*�.����0'8�^���Jn?��i�#��#>
W<S]�^t�O?@=[hU�,+��\2��H)��t�!o�_�����Z���%+�?�;�ɤ���9��r&"�z��ل�#?��d�1��Ճ��i�cV�܈w4��@��2��µ8�7(����l�-R����S4
���^��c�zm|}H��ia's�cyo�=W|���V�w��.���EѢ$fޱ$���\!���: J^็�> J2tÝp��^FI5�?�U�%l�e8D��u��_6*j��A�,��)�I79e'�t^+C�>�:��|�~[��j��� 3Piq�
�a=j�&AkE��t0W���LHj4�3�~�Q�Ps:�ȱ�g��#����V�i\;iݙ�g���(��Ц������HI�i��6.Al}$�5(�o�h�B�l'��r�8�h]���q
�W���듥X懲��?č=��l-8�����V�.pe��՟��dѢ��.0|��� ���d�y�`�ǫ��^~�M�:�r�����ě���S {ؠN}�(�@}'�Tc�o"���f�l��	��P�!�U��7�z$]$���76�쑙y��n�$��rl�Ⱦ�[O��LT���t�~3�K��eh��]���  �ֽ���xw�j&����5��h��o�P��<�Y����Dv����0i�Y����2^�	Z۝�k�3y�հ)�?;d6��Q��<}�ޚH%qW��9������������j�r����
��tXU��h��M��a��Pm�6�ή�l_�6&��4�؂�"I7"�\�mWƾ��GZ=�ِ��xè�0�'�l�}K���]�"�m���7�t*��a*�}8a/���J��̡��=l������w�ۤ��vk��"�aa͍U�f5�S�w�D'�F�f�]��������B	9�K�	��-�q�>4�s�ے�Q�-3�t �{z����da��Dv�ͷr���\B�2�AW YԬ����{��j2U~i2�������=�1;�
�f2�%%R�$�lWr��`��n��
�'����x���iZ�#3P|��Os�,]V�h��Gڎ����ެ�R��"�̊�B�޵��h��~�\6� (��/DI�`� ^�.�T{��^F����ts��.9���4W�ג�K�9���Vp�U�1�&�T��)��(�-��BX��=R7����)��H�۞��<zG��x����vzĴ��8��q�q���A%y�/�3�o�jf֭�&��?'����*�<и��5�I	P*���ܻ4�l��$�*O�Q� �K!�0b�=~=h�)zj6�� �A+l($���̖�^2�E�n�������޸��ھ�T���e*�6�
l-W/'4+����� Ȇ3į
�e�R=n7��V#�'!�>�OS�9���\�d��/���3nb>���H�l�k1w	|�/��Y�R ¯��=M�=���T����?��S�R���
�[$XX>f��h�G
%�� fh�ȠT���)�����\��x�soVC|�͆l��ᘿ���Txo%�4������erӿ�-�6<gp���\d#�d.��2�j&ֻұB��>��&'�A�>�!dD&`�i1C���EԸݻ3�b��P�y��ݬܗM��Ai�o|����"�\G�|��bMCC��_�mzl��h�Z)������-��3�{�_���ūqҽ�Ҁ\V�Q��K���TB�� P��*�m�j���*((ZB����zi���
�~�ixd�P4���'�ꖌ %��*B�[/{A�0��,̜ܔ���(��Ba�o����_R`�m@R����S�_�i�ny��d-8�V�TC��ށ	iq�W&����b�kꮶm�]�O|�!��k)�)j�|��BaKKƍl����+]��.k��'2���Lů #L���ѹHR��&����H8�IO����N�|�W�j�]X���_�U��W����Z����3��ȟ�Ė�:=!Ts�TX[�Dt�DtG;3N���oUh'w�>d�E�E��&�q��ܩ5���T:�qq:$�!,��B6Ⱦ�
�m����������>w5t/��Tl����@��ll�XgN@4�^P�@S��M5S.��g:l�L�ID�DE=��N}3���W�}��xZ�mϋ�~F,XA���3 ��粫���?R>��4>�m8$0��W�?`�ܽ�?�"'a�p��+�20]Ca�Jf���^�:!3������S�'Y6R��m�l���)o���+�;�`��C�mbLV/���OVjy���MC���E؄3�c�k���1�}�+���	���
�'�߫�)���eu�y��f�X�˱��qm��l���'	?�5T
f%�
�zd�@����kHX�����2(�gI0����,Б�g���Sc����0Km���<V���Ӟ��c1����{	������i���\f�)6�ic)K�Ng�z��)����̱{�+%:�WWɒ���с��a��ZDYS>�&���Qaęt�iCc`՘��0��ظ1L?/E#��د��C�y��.(��W�a�������נz�t�b�	}���{�-y���~
����Gdj�+���+�xj˃r�aG?���9�L]'Qؤ��v�~�^�e��҃�l���W	�)��&K�7�v
b&�J�(�c9le�Kh���ɔ|�v�w�h�F��mW��$E���߅E]'i�a��R��۲�:��=@0�k|`R�~pp���B�S"+7kc���){2���[���"�z納�}���_�l)
��С�Y�����>�MC��3ܵ{��aW��<�	_����o9Ib�m��]5w�~�y�8ó:آ�#U���!{�4b�
��eB�L9�Z1��<D�%�@GY�|]a�2.�<o@���� ȨK���Tj]���~�^����3Jp�o����SѾ�o��V����/�Sr�TE�5�<ϖV
�
>L��x�� �
�#$��D����#�^om.>����|W�*{���U���0H�G����g������brYy���t��=��0[V �E��^�z�^T[� R��'�U[�u��Pd	?"N�n'l~�P:����>��JZ������'+Fd�Wl[B��8]L2�io� �5o%<��@�.���FK3�(������;����8����v��"TQ�I��5�SӧS|͒f��4�D�@��q���I���a>[��Rq���2�(-��"����
w��4_2�C���IV� �ئYPK��Pgz(K�KR�Znǫ�v4B��d�Xڑ�\D+�7]:'�z �3�`Z�+&���i�^���'�l����_o�h�XG��&��  �Q����ٿ�uJ( k� ���PЮ=����J�>_�[?ڒf�$Fq$�����ě������U��-H��N$�a⮓�>�[�%���eS����6d����:��J!���p;$��"��nR��᠌-8�`��D�����k���E?Ǳ�7��r�l��JӘ��ù���1nF'�-���Gm��M*�8� u�M���h�����y�+�Uǔ=�z�X�|>6���DEY`�+I7�YB�Α�=������ȳQ���g�����kV�DmnE[lM������g�"0Q!!���}|:�*w��
��M�*���3pI�Ӣ�%�j���_�K��?����{�Y��:'Ğܞe�0r�ϵ���x�hQՁ�,��J�xH��k�CS�:�Q�|k�5�c�E�X
}<�`�C�@P���p�2M�lt'
�Ljc�D�bῳLT$�a�u0䘧�����X�!6�j�z�B�y�&��?��[=T���jM^nvg���+�@K&R�[�_ER�{c�H�9��a�2�����v�s�T6�{xѥ�땘�ٚq�8c�i^�s�nn|��	��Su�tv�aDg
�|椆I0" p��$��@�����ũ�����,z[b�b���Ew.���|�y풗NP���z9��2`�ٲu6���h�x�w���ۢ�j!X���>��t�.h��[w�M$m���-��|#S��;lm��X�Ru�E4Kl����<���J�	�y�u�����p��l1b��1��ʺ+��8[kcg��_��bYF�$Nt�$"�Ҏ�p�Î&l�>�7Ё8~��V�F�Juh̦_�e�bfy�5}|�U�t�)�#.^@�"�WŰ&,��[�����]3�yL�X�Ke"���A�L��%E�N5�W��;��Έg�����]U��� �U���H���ƿ�`�xC��Eɛ�<��N� D���
�|޲��(1�kn%ײ-�3��X�\l]@K����^��W��\�u��$�	��n��4�5�|g�￾�"|�7?�AP�#�#5��ɪ�W���+ħ)ÿ�* l��=�!�=����L�����}/�f���th��V
NU܆z;B�-܉�}���#B�yd����Vy2hYz �(���To?�X|1�0���Մ��H ��p3�5k݈�9Q\��k��Q�����N������o�)�_JU�N��7�کz2L�H�4p:�Y\:�̳�AV��K�C��٬��tQ=+I:g
1�0.CwO�94��yPE�lI�/p3ϻ�^�
��<�4��kx��*�%۳~N�+J��K�y�H�Ҋ�>oEq�x��7pV����\w\F,T)O/3Z5��'8�����EtPHf��������M�p�y��P鬲� D�[�����V4!�MX��*�'U��T@0}����Cu?�w�A�i�˯����:қ5@���rM���'��T�M���	�x/�+{Z�"��Y��j7��W�96� �6T�E~�qK�/����&�<�H��/J��օ蚳��h���Ηc�q��P\��瀷�r'"�}�om#얚��+�J���]��Tƕ��9nE�S%Oxw�5��I�n����lt!+��~�4��)d�(��(B���SZ`�8�8�4�y����a5�B�	��I�8|��#�ETW �7�"�"L��j�c������ ʷ�����P�K�}k	�WX&���a=������bU\P�����9�M ��Ы���X���O�F���e(���(5Nb��/�Yإ��{[�v���h���0~�d�:���ԫE����EZ��ĕG���{�*x�����<�o�c�J�r\���WVVi]������������C����_��Ɨcc���yţ�Y̳/����ln'��.��.M�>�lۿެa(m#�X�VR��0�&�rOו�"��kxu��)���q�&tYNK�|i��r�,
��u��]^�h�����NK
����Ӑ��M`s����!�ZX��)F���-��Uiʸ�<A��݄Tk�v�a-�~�ah+��ˠ�4JQ!W�SL;4Oɒu;�6��ݷ`�wʬ��I�-/x^^�~�&,b!���]��Q���C�%mQ+�6M��T,�i1Am_��禬
L)�V��rH?p��j���O�eI�Z���eQ�c�2���+����{M��	��bd�:�-i?۪b�xJ�
`EI�f�ڕ:��]/��ۥ:iˢ!F�ɱ����"$9��N�:7�M�<�	W� _>5f��BB,c�FЬN�-��ot�θ���Ϛ�8IJ�2{���a�J�g+}>�~�- �#���	�d(��n������1`͛V��)��MT�x:Z�����HV��o4�"	R�("������Y��g����9�s���P��~*�B���.����o��O��-��"��HYK���?�:e�%\,P�%�hЉ&�ur�})�JJ? �g���0E��؂�Dv�c��}_.c]ID�H��KG�Q}��#���޶�u��Y!V��An�c�Ķ}w[�*���=�"����$=���y�G�o0��k�܋6����NW!��x���HFo�ɸ"JiT���T�O^��\��yvc�N��أ05+�U�^�(��J����3��ȉ����Sf��.���?�eԬ�|�m�Gb\��fD$�!���َ���N�3b�,;�h��t;���UFûI�ES.��d�L�% ��G���ߢU�:�H�O�@$�1���I�G�T�<!����+j���/C
/x�vf�)~
䯝�ެ�o؅��MK�s���ؖ�+�W�D�,��Y�SI���p�Q���bTt�L�����7_�-e�h�`��h�x��(i����Ny�f��r�پ�w�v/4l�k�O7�e�pz����F�1s������%O���@��v��U8l�{��C������p?4��-a=[H�lO�P�d��E�sp�����rM�ޅ�V�J��P�5��/.�Jd5J<�����YC51F&��B�ʉԒL@e�Qӥ%�����ނ!����H�հ�b�/��rtFf�ʹY�I�u���¡��ZN�r~wl6!"A"��N�b�a�
��ݚ쁁I闉&.Sy�֟O��]�A�t�aҏ��5Ӹ	m����h._-t��;��G��v��Ff���O�/$.T�^�9Ɗ5������Ȋ���S�޿��.WNN�g���)��^s�DY���\S{��5_kXjoL�4�P�v�����_�#y+�`[�q��,ծ] M�A����
��dՋfW�OecZm	%�^�+�F�>�Ca�h]V]9�q��,�ةH7��b%�\�Y\��N�1F%kUOs^ό\��R���OUv�_mqK��E��Z���v����aH�3���S�:�);-ׇR�IV�l-n����9y�VR_�:��X��0���ͮcU�r&qƵO�<9���$�=������������O	ȑ�S\�J	�qa�#?g�ԛ�@ŧ�_5�>�ʆ��#�������W͚>AE�i(��c'���?7X�TH��0�ϟ �3��&�´��|�
�T�c]���(��mz�&��P�R#4��Ό�ϩB�O���h�X��8�:ò%� y��y��(><�ྖ�`����Fa���n2�����A&���<��2��#G���iz�~���s�Tz�	������������C�a�'ǢDmi��U�c�G� ツ�%������q����j�!:���0�_�;�!���6���䑱�7�1f	��X9*���
;H�L�r�m��`v?��=�����i��	O%X�>��)CǗ��M�����k��u�}���x*��΍9ǣ(O�b��
:99�0��OX���DA�=J��fo�uˈ��Jn�;ƿ���:��L�R68�Z�wu�@m֏��?���i��5�>Em�O=i,���u.m�����Ϭg�S����ė+�O��=�>�݈�P� 	�2���X�}I��� o҂����5>�q�v�q���sr�5ZN8{�#�wjn�}���tU	�k�l\pm����3�R-)���Z����?�c�Yz�.�Qִ��)��D�HG�O#qF���&-Mrt"���2)t�P�;#2F�$vp�~1���d�R:g��޲�T�2|���%�w\vu�Ǥ;�p[�L���{<+����uP~�`�P�g���;k�`�n�2���^xd���Y�nԓ�8Ű~��sWu]�����G�܆7��M�ˏ�\Q�7A��,h��]ƈ�t::��:�[p׌K""
^y�	(�M�jr�K���k �], ��֔��{��c��d�Yz(8��W�����z�	 5M9�y������'�m��j/�z��1|���X�r��E�a#i��{��>U�՗~�]u/̠�˱��k�GzYzT7X��Jղ����fBa�Ĭ>��Ꮹ��yu�=#�F�ũ�"G�fZ��uCϲӞ����Ǧ[N��X[)S�D@ˀV�o�B�ğ��ץ��1��Q��'"�CЊ����L%"�ؘ�4�����L��6f�4owd�LwJ^N�ws~�i-+Br��B�"��(�cs_dG��*.�,�lc��ΐ4$���pȀ ��U#)N���4]5oK�v��C�Y���K���p���M������V��������*�F�^x�]�k�������a5�n���y��^c!qzr�b�����X�]l h��Mfx�2oY��S�Ȃ��+�|L��yI�â���9��{�M������ђ���YNt1���1t�wE0�|��	V¯��Q=Y�P&�$���.�b(h(!+{KH�A�"�.O����VڼxVD4��C�h}����<�������[�Ƀ�����¡[���bC<J����¾<���s-��9������I8�AK�s�ג�{���)�B$����2ɗ���3��Q%g�X�������Tn��Ds.�.�OK ����5�LU�Ot��X��#�>N}�;M9q�:G�X�����D��o�q�oA�|e;�Z:��%�N��^x��mk����Ve�odl>��Q��E��?��>�g,Yr����4� 8y_,��3����G�]��%f�C{��uz#��E�)�[=��UH�U��G�~J뛙/��N6���YjhW`*��ܘ�U�ӭ�����i`�).�d:1!���9�0ZIQ�1��u�&�k�K�f|M�H�X+W�u���Ҷ�h��(0��RT{�u+X���Ͽ��m��?�Ym*X���7Θ����|����ph�w����K��i?M� �'�C�Px���Bxh�=
Ȟ ���1���y|��~���u�ݴ��D��a<�<�Y���L�B3�6WkΓ�)�ỿy��?�g��
�ж�
���F!6&j״�d��Š� ?r�r�3Ղ6̯���Ɉv���?�*��JH_��"�������>�?�o G4�����5�}Ŝ�%���g�q��(������iBsX~���0��~��9�6R�\�)6;`�ǆ�#e�*�x(p�g?T(�8�l���q(��ܐ+Kgp���Q#���߶bk�_D�� �i��s(�H��'V�|�����:�
��<���H��qWM���ra�h��~�ы��-7Jw!���&%u�}3#��C��"#�#��+{�WX����x7�{�b���I��QT����L���|�@�����Xn엔����$�z�f_,�{�ӫ��� �)ȽJ�����g��@_�	��,��N����o29���p=Ti(�N�v}���q���z�4�v�㑑[�&���Ǒ�^��(���	:v�(����[��[�X(@�n0i̛�b��V�?\���qO�yػV֥7�|+���GW�f)���)}�I�g�Z��� A&�F�n�����3T��![�{%�e��\U�.�93�A�&�Ӌ.��4Շ��Ը^.;�+�j����_C~Aک�,://Z����a/W)��_A:c׃�⣤0��.K�`�X%��t���2�DI�蔛�"�:�o����e?ۃ��8 5\�������c	��1N��RK�Xb�ve��+��#�/�n҄2�_w�I�����X��3 T-K�pw<��n�:��{R{����FM���;���a��F$��Ոm���к�Bq�a_PW�r������^%����׆r�"�t���vpsZ�Al��+5�S@L�(�A�jC5�?�҈����?�B�"�E(y�2W��%�RsF^b��p��K���|�N/�%9�p��T{Tݏ�1�8���2أW>��m��ӿL��z��� #$<[K���&F��6{�	�3�s�
����;�5��T♈V.�օsq�y�`�ge�~�]>Њ�Z:�~� 됦bP���n�]�$LDWkDr%b��@#�����u�}�^&n*�C�0�k3���~CY��O^$8^)@�FB
5Tx�#���&Ԉil)��ٻ����uA[�r�� ة��cR3�X�*�'N��c�6�|L��'�d�*)�nrU�l|u~nv��	�Q��G��}���luQU|���.�f�[�T
����R��swY(��Q��U������fXM�>�;Hԡ�z3@�2+���+ۿ��4�C�k������4����wʵ�eb���y*�Q���O .�%V]H��������I'�g�T��==�j�QV�)0�g^�7A�.S}�\��(r^-��a]�BNQ�z��%Ir��T���h&z���%y�K�4V�:�ʴ,���K<H�0t�K���ҍ���ӕ����b{Fc�Z��vy[h�0��R4�Oa}N����z��̧V���*䐳�s�4�D!B��A���S�b��?�V�����'~�Ȅ$�m �i�)o/h�a�X��$�V��Rf���Yu�<8kI!�E*��h��}ft�	���yj�������륧|OT?�<��U�!�E����!�vm^��D�r �|���DW:����렕t��[6���Y���i�xhs�Jd��dK@�y%ad��^�t	;������l�U�Q���L�]j�@�/m`�4c	�=��ĺ�,���mU���w�T�Ar]��Ӵ�+fQ,��>*�,]����_.(�"WƂ����-Ng��4�T<��d�ʞA��W8��W�[i�K�h#�Z�����Љ��8{#zw�7�,z��H�D�1�a��̅
�⡁ w����[�Ὓ<�!��@<��+�P�����bf�n��R�P�M:���_��ey��$�%��>��y4�4{+Eg#��3��m��m�H���xk�g���^(46	� 8rr#�+?��CP 7&��P�XT�����G��@{��B���]sA�v������LC��ޗda�f�=	[~/�����n�oU�J�01�m��q��'a����/%�D��s>žt�@�&t�i�Q8��[��;����21�Xó��[�;�����j:馵����ظK%���ހ��tă�k
=�v��"S�O�q�m�|V��Z}[�ug�o�{���ow�y�M��C�"KL,#ޭ�'H�Q�Q0�=o7�x�"'�B�A_�U�'Ҋ�ȐW�Nv�Z���°[�|��?u�vp?��B���mS�q�Ze�!4	(w�*�$?=MWf�p"�X��j���]<a�o��6�ʭ�{��Դ&|�,�y���:T۱�d�I�~�����̘�a�0׫7)�=��"vެ�⁡\nAf�S):{1�[C�Ti
���Vο�c��� Hx����Xw��M��tr�S�
���E�1��f;�p��o�?�Ҏxu�,E�b=�9���7�	Sl�P$���/�\�,ц�y�%j��zF� ����r�-���gw�u��K���Z�%Ͽ�{`�r�z}7~b��̭�#ov��N�>�Չ�
k���ps��#�F9�ʹ���Ct�.Y��{[�^�9vUyF|ti��$wF��'�;,�wH��%�X�G���x��������%��|�DbB�X�r(U�t�־vx.6�������<��$栙��0�t@�o��ɥ�Ɲ3o�2��m�?�*�ߜ ���F����.�Q�q)G��X8ѕ�k���vWF)�{Xʘ���kʢ�ԭq!�Xn.l�!�Wl|�ea�6� nZk��Srr@#�;����ʥ������Ў�娥4&+�� ����U\�)��ʋ=�ڹe�pq�|w�}��X7�{+�� !��7C������qm����"�ɖ�L��%�P��$�x�G�%8�f)��â�:>bQ	�S�Ч9���u.��!h��aW�p	\F����D��3�|��3/%�,Gb��_u�,�G�T/�^�=1��W�����Vsx�P[ЙR�Ȓ:���^��TQO��A4��^g� �d��=~nz�Z�xY��f�m������Rb���(F�-t�y%H��'�W}R���O}���gS\F{�dT�B#l����ɿ�3��ݶ��g��w�%e��P65�Xz���2B�H6�,��-�1V�����
l=7����/�ANjݧ�p.~A�B-l�0���줒%6�T#
\hj�ܥ����YL�[���	e]�R{s�h5�*����hF�H��&@�_[[E����
�Us�P~�Jt,���/�O&9p���.�fg�%�!;�P�f�ėX.:/��;c��F�Ik�<TbyS�3ʹ���z�/���`gtX�~�������<�N �e7�������W翳bm�bp	ڌ><u�x�q��K4�r�[�� څۙ�-��[���k��G �Wl˹����>��,��w�������2&$�|D~Y^���6���@��s���:S� ����%���vj]A�sA�k������+�"�L��,-�3�]Hm&Id�V�����'��(:>�/�2�[���L=��׶�v,��Z�(;�1���2_̍K1�D�ǉ�\(��Vp�)0
g���৯5�K��ԗLU���Y�f,��ɃI��`K�`��7q/[�`%:k�g[��fC_�y�p� q^q�A��z�\���F���I3�06�Tgn��9�*��/a-r�
JƠ �7�C��{Ŵ0#sfEn>��Z��d�5�M�hӕ�	b}�U���mL^+i$z{�S���Y���h�]�=�,/e<|�7)컓$�l����B�u��c8��¶U:S2�<���VJ����֛*n�])[i�_	��$�:q�8������G���C�G�4 S;���K�'�>�z59|{��m�1���	)xֱ�'�,E� R�w�����ij���6�Zz��\�a�G�;T�+90�"���O?1ﮙ�=��������mL0��iI]�	]����y0�h]RZ짠Z���C6�k��_���Cx��կ�Q_�N�d֌";���-�K���&�,��	�,���[+%�`ǫ�{h:g*�_�)����]&��Д�$8�B4w��ֆS���L��|u���w�������q��te�Jýԅ���-	��jQ�_�S��&NS���^Љ�����;����.�)i�u�p*����A[�]f��d�ʹ'�k������ǔ�3��%��.66�Ftz嚰s��[��W�AD�j�}L*,����E�>ȱ��Qu���*��mXa��ܙv\c8뛊��ș�=����/�\v���hs|"J�U�"��o��1���U��Q"/}u��&ex�pT��=��$����3���-c@�n�j����/��A�斢�n��}�nKER��|�
o�෺:D �^�um𔾧j; ���Į�P}�<u��r�L��O>cYo�b<D2?���;0{���S�?H(�r�r}&z�h�����j�C�e�(����ꒄZ�0C�ȋ����������ػ�؝<�h�eMY���^:�t=B�4:"m]h���sbϞ��MJ�{[n���C�K�`��Y҈_G�.�o�lL��-����4�Y��.�)H3H �%#�DQ��x�'�}Id���1���=�)�8�j���[�B�"�8uY3���Ԥ�`a$�����������i8�O�?�s�{�)�(�(��%��uw�u��}�}��<������d��3��6��/�5ųp��be0���E�s#�V���m�%�N��q��4��X��U�[O�!t�����^�w��ǂQʑ��`��4!�U��s�xk�mL�>� ��tʶ�d.�F��d��[�5�#�|���EP�x���@SLዐ� ��_�;�L�j%O��f�0O��ĻSt��r���]T�7Kʾ�H�@ٹ��~s���⁙d[��'�����k���o|�;h�Ծ���<��/��_{�Q���B�Iy�8O[��ڎO_�H�r�,kܡ�R?�s� }�w��k��߾�yB=������|�]CU=���U�0���% IF�\�I�;�Cb�LdM�E�[~�N���A�����2?w5�+���N�/D��%�u4���=s<ϥ�V�_��� :��ǵ�� �NGs��\�����P79���|?�;%��������ߧ'�����UAz������Äu�7��4m_���B��Ik6�%�_� )�ID�v�A+��0�3�z��@@�_�'�T�MX]��"��J�tJ��ˢw]O��Lxt��Q�)gW&?O���r���e�W�|�r*��$4+3��<㱼�Fϗ�t�C`�)�Q�#n��y�l+�Hs�l�rhlQc�-V��M�+��T9��;��(�b��7�&`�5�FdO��<��P��,q@�O��PH�7N�u��ڻ�A��h.���;B����Mt3��	iu
p�g^K�Rn��x�:�r#h�o��7+�70�h&/v�Ô�hg`M"�-}]���y�x��ŉ�P�n�IOؑ����='��lПÉ��#*KU�E<�.�P{*��uȗ���]�]���ʮ*�����*���.�%/����E����
I0���/�]�����Ua�k���=~h9�_tBz9��P��g^��v]tN2�⣆��>�p2�3l��Y1a�ǣ�G6�nFG�����Ż�m�d���N:��s%kv3�o�r �]���XL$���wW^�'�e�]" ���A?�P�#����"�:�Z���4٫@
I\���������'�vC�Eᤆy�c���L�d�_c<i���#j5��ze'zK%
6�����9:����F�(��g3ꞔ���
h�D��.�dl������3yBk�����-���S��s�7D�
�c�Ћ�W��0 �[�E�N��j�^�~�+`�4�����{G�#l�R]�H�� �Ð��mmp�3�(gN��4�u+���$�.�"�6�x.�%�!�y�^gƣCz�����?D���s����ߒ_��<V��SM�>+�$����Y��F��N����2WR�YtlW�9�p��4���RR�=�(�x�BD��c�(u=�V7@�x@6���p1�ʹ3�G��fF
�|��{Ȱ�q��N�׉A����*�¸v��-�OH���f��y�<L�@���&�F�C�M����i}г��(���D���s�Z�1'0|�J���>E��`P|����Q�v��{u���~�7\�L�舦����Y}����*^ubk|�6e>C�̹��<�����$vjW�k���>���GB�λm$�-w|}�5��eO�Տm�9�Q ��b��O�n[��m���JM�==�'��5�}lɎ۸`���L� �]�I��/·��x�Ұ�ćB���τ���]�u�)QE����+��<7nÈ����{�h%���(lr;|���m�l &��ۜ4��*t�������JgO{�'���h3Q]?Rկ#�c�ǎ�̠�]�T��`���6��Ǎ�����n5��!F�梓,@�4���&�\=�1}�/	�=�8�Xo��h�$��N��m8O`�i�zt;�Uw|ņ�l_�gud�>6�x�f��fg�/��u�� ��&�E�k$oUz^��E��b2��tuS�j(\��]13�V�Q)  �y[FБ�#^,"¦x~G���wU�5�Y&�,��s$�!��]��A���c
��aی���l+�H�S(�2���_�L�]��x۲D㷂V^�����K�i#��\��@�Q��;d��@_Lb�L��6�0N@���(tT�f�.����i����U5����F�\�.V���鮥a)�/UY�d�2,=��T5���-1_��N.9*���%�,�Zu�i�2x��qT ��xѱaPX0�F���x���s+?�%�j���3
�x�k�3��e �E�:/��$7�a"ML(ĩ�(Kv�C�b4��$���d�X0S��(")��q��1���j���e+�
cɂ��<7_ߍ�3x�b��g�}�y���[g>f�4]W���hd��d�S��)?Ņ:��p�3��wb� ���bA{���;�����}捕7}��F�o�5h�/�;�IP�G�hN�*�"�����7E+��R��nl��T|���i�.<�(��>�]�+{y����Lh@��\I����v�K\������2��
���
K�z-Q}"�9�Yf��*��}��<|�xM�u���ZA�b5��:uҬpV�PeM<hL���,��],+c㇦ո�06ZI�D��W�P�o�^���'����"53�\�n�7�ߩh�e ��O�
��{M����Z������}c����>$�����^$B�Q�v=5���_p��byUJ�1�J��e����v��.���n`��:a]Ӭ�M�`g����G�ǀ���`��ڨ�'���N��ͅ>y
���"]�[�l���d�#0�i�`}��E	L�0yu�"�W�QF9������ � %����m+䰴�pQ�{d_/��j�	�,�[CF�s�#�z���o(
Iv�9������\�%�$I=��?s�h��?���r���C�L='�N��?�Z����i�K�/�9��؞���A�6��x=�I�[g��D��	�˺ɲbI˙���i�Zz�����_wiэ>�|E���3f�Ď�����h��pK�	
�23I�N�� 29Sjf�Խ�a�[@��c��'��[=xB�h���J
w���hҳ	ָ��[�K�?F2��+B�7Hl�����xJV��g� � �����a��F�	S GIZ���5����9߬��}H�Y��u�?(���FVU���K(VfLe��-��Lĕ,D�08���e�t�/�=۱��K98�D��Hhk=7)���dq6#�ʶj�
$��Pl��6�M�S��(�Qo���qr\+�^P ���_YծW�^	�{���f8]̸��~���a��À�¿�������]G2Α-�&�\�@�.z���=�1G�b�S:�m�D��$c�������G�j͑>�D����+]�,h�QheĦ�#Q(��M��в��jG������j��p  ?�8.��|������].�d1�)�u��3쟬��{A�g�� �=#��ϔ������{8VS�zʯ�\����z�� ��D�؇���+-(�	J�̀R�IV,Y5�xl�$�������Y��IqĿ��UE������ib��|o�פ\�����k�*�����=y�N�]?ђo�Ϫ	�y��'��au�(T@!��_��)���4`&�Y��<����S!eZ�h�B{�W�THn�.;; =��s��o��)�ȍ�4��`�k�6#�̞I���MH,�[��<=t,c�#��\�MG�l����u������w:nlw4w�+i�#Ź�M�ݵdD��@��粷�{R�.�T� ��G��y�d�p��Zw�ۭy�'mv�v����6��cz�d]�g> ���N[ YS��I	Ɏ����9Kӓ�ܻ�$jo�~��uǿp*�A9�C�|��xK�zh�C���E:~�h���^��ɕ*�����e(��k�ݤ�)�(>k*o�� ��&`*�5��a�1�=.!&au�,��y��5�imK�&?���LV�V�x^�}��z�`���sM$�~�V��j�=���=ї� l��a�$�Ig̥��#;V~��k^Xߧ
�Ȳ��R�Ĉ� �:̅��u�a"��{N]�%�X��a��P��^ɂ�E}$sֺ��=0CB��;P	���r���&lj
��BdO�ߤ��=6 zD���$l�[�`d���}PE/�����V�䙔Z=&��SG&S9r�G�.Ɉ����x�@���dK#ZW���,�_3���m6$�nU�Q�|C�J?�<��"mp�`�j��P��]��n���|H���K����I?�Ǧ�O_DPW�������/���;ȫ���t���4�7C*���a������z�)���h�Y������E��"�JVhX��o�pA:C/Sϳ�� p ��[ׇ�#��Dv^q��u���^��Vz�!<!�-�)������j�͕��J��;ͨ��~7Ɗ�S܈��D������"���n����d�U{��A�0��.$B�=Sޙ�D�aD�W����E�"9ظMIb�C�_���3
Lw3D�Y6�S�r�B�c�Gj�ڶtg05H'1�0���u�~]5n0�
�.(��*��Cs�����I�5%�O�i|F� !�4���l�x�_yX���H�_s_}�����q�eOm(�����B�RH}W�}5�.)�L�G��y2R]�"1G=S�ؔi���G���a A�K����K˞7�Lf�=O"�H�S�G����T�R]���5ۅ��K�`P�M�2��7.�-!��Z�P�H����?e��(����thۊ�Y��@��Y=����L��)<b'fW=Z�\&��|�3���H�C��r Ǣ΅9���\��:�T�M*d}������1�dA��4�"t���W�BŌw��j$q�è�[ݩjo;��ۉd,ub{d�u��a��H|�U3�u��L�f<h����^��z�"����%u��}��5h_��k�Y�5��@x��m�پ"SȳJ�q�`GQ�@��?�@�� Wn�)|I�+ö��>YxC�	�}KWP�99U��s���?�J�iS�MX=��D$���Z\�dQ���7��s���б�SK�ݭ��x�TZ=�q�B�7o�P�`�:%��Q�@D���'���4������A�&���k�H�k����7(���:�12����7Ϊ�x�Si����9Mt�e=����=-&�=K'KEvۋA^�9��-qA'R��ҮO�I��~�2�����=����RfZێ�O����[R��@"IqY%@�@�+�O,���� ���9����#�Jٲ��G^�Ѩ��~�[-�����.=Ĉ�Q��o��'?��'1�b�38~u�Sk���cu�c.��i�1~�bƁd,���&�f��Mͯ6����N5���FŲ��hʟ�}s�ŗ�!`��2�h�SSov�b�*�Un
$��X#�[B�q54�󎮑��-������f����ŀi2�{�*(��$�ń�OS�M���K��C�H��	]���~�Տ��i��Ďn�Xn+���[��8D�-�;�?��a]�Wl5P�� :B?,ԋ��a��ꂷ8�UL��M{��v���Nd�?<���1���l��tkb����%����fYd;`+kri��q;O
��>�s�J���̸�蝜`�
�	�j���n���,+2��������}A=J#�EՙO������O�K׉{�z �ʨo�8-ꯪ�Rh��1��l�;��!|���amۊ�����Hqo����*���?�{����9�
�ILXze��h�+��L�Y�
&�.()�j���F�Z��ީ]�O��S���o�N�����S3Lh�!Fj�W|�o��A�l�?�.����s�Z� �'�sR�L��)�BI��s�݅w��69�y���	Z���]�^���LT�
��ӿ�����bNT志*� mR�����7�촐��n�nd�ޫc�^^�,F��B�՛P��V��#���H��U�wT9�~�Ù�!r,d�
yV�\0�K�ղ~d��2�n���Tg�b-���@E�q��d�����N˹���d46��c˞��G�xʌ�Q�^������:̃A��E���t�1�8��\}��Lod��mzJ��j�F��>�'f�BU�k��D�`�q�=>6���#��(��/������ ���r[�b#�,}Sv���>g0��Cu�Q��Ч���V�pO�j5?J�3V��1��bl������2��a�X� �{mg�`#Ц�}��c!]�|>�w�����EUǼx1��@� �UԓO�
B]���ᐥF�����"���r+�lR��l�m���p��
��\����9�-��q�R>[
'��� f�U8l�o"��uڡ]�q����{�sͲ�b����F�gVa�~_v/���߫ڨ�]��9��k����J�Y��Id��m�ɺ ��bҋ�ϙչ��t~�!�Ŝz79C7L)i�F����cl̙��/��͏��8��4�#�р�j�9��'_B�x�Cx�.k�f��_�{6�%����AtI���_��i��� /A *��b�x=��1��_n��DсP�A��6X�w�᤮|A{/���:b�,<�:8�B5�Nc}� ���f�}Xc��Rd�%j�S��{���΋�_CM�H�|�PY�o;mT=�Cצ<3h@��)Iq�_A��'BD�u�9�+15?��X�C�(k���<q��#PA~dr��%��)�.�p����p��������ח񞦢J��P�'�'dy��� 4�;��'���x�98�����qO��hJ���BM���w��L���H��X����]r|���C^�o�Y멷	�y�)��"܆G�:�%X���Of��̦]��>�����}t�ǌ@7��d0d��䗹9s\O��y����J��X}B�o2+�tiO9ٕ �'������[��n+��`��OY��� YD���\{�Ê��=hv`��讣�F;C:��&���Φ��U�>*D�� �� �	�t��z��p����P������=� w�����;x�����u��N���,���#W9�f��G���>5��uCc��e��]b�(ՙ���5�Aӻ1��IP|��r"!Z��!�	���[:=��5����P�֕��v����7��GD�ܚɬ�+�-ÿ|�C[�����Pcv)�����Ú}8*w��E���T�|�ί	Avɀ�9z�݉!�$�5���