��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��� ���/M��ٻ�x��h�{�縊��D��5No5��L�p6�,�e��{Ƃw�Vλ�66[�^8�E}~,a�V���ApӼ	�l�y�r��cb����b%˂���w@N��~d^���4D�E$Cגߚ���kt`���.��C�3J#���)5DM�ߦۊ&V���� 3l�F�,/N�E�_��	��%��.~��{��'��/�n������Y�H,��w��0E^<5Y�=��j٫�y��w68R���5�Qʍ5����~D�	0f�j%�c��3���.W��S�Nl�n����a�������)(���ڂAC� �M�oC2���U��	�:5�u��gr�������5�su�L}��S�e�v��x�٬l
n�G�w|8;Rj�7A@�@���v.�a�.䡁lt���������m7�ȋ���rL�qVk��NMX�r��(�Y+��h�����FTj��ŻBy,M�p뷴�"���*vI������S�L��]K("Mk|��3&�@`1C>֥vfa�3��w����H��s����b�?�$q_�H�$�L�o�A�����q�i،�H{��|���mHW��A����N}
�� ��i�R������';g�:46���Iz�:�����
༃�E��`ԩ��=����\�D.OKu�|n�Y���PQ�qJ�ڠ����,�����Q����Z�;T��	d�`�Cf9յy���ԵK��'C��,��W�=�%�J3J��;X�@
�lN�B��=��]v�ɘ���B��pP�θQ����A��G��Omz\�u���"~{�r.��PQ��sz.T_���$��i��>^�����Ň9�6:�'��F��a���T��l����P)�F�&ۺ��a@@D s�4�ql�J+�>.B��M��7�b|,ݚٿô�	����y��/�^3�Ռ�)4*��F�XVI�� �8�����<�z�J�8��g�&tA��, x����S�BD[g��ˊ����ȋ��>���HQ��T�7f{��'�E�k^
m=8�i4u�������t����B��l0��\v�u�P����B�ל�B��E1 "�gD��<���F�����Q��3����䚤����,�N[�NQ����>��QY���fN�o&/7}�H;ݢT�����O�!kz��w/��k_}C:�Vd�̩1�\`�1[�o3�D�u�����i���km:�H�w�{Fx��w�ۉ���{��Gόy�_����a������".�1�\)��"�VK�RN�^��v�`�[^z-�i[\���~g嗌6�vl!��5b)2��:rYw��ᎋ�4�XR��!ybL�Lj���j�2�w�Q6_K��E�s�xCd��$�N]�ُ�6�� ���X�<��d����z��k� &6UH�,�ڵ����wҔ�(�s.^�U��"�?Cai�S��4��O�C�W$�W��{�7�##�p�>4����[_���ȘW|��$��<��H��ڼϬN��}�RXw��T�Z"�WB���@u���"{{;kt���(uxʁ7�Jh�}G�b뿅���r�[vշ��zI�k�=�K_u4L~�<�i!0��6����>�]rGk�^l+OW6�S�ʸ�ۉ��
dbޜ���ջ��3�?TbIc�M����|h{��P�� ~;jp����K˖Q*�\/f�$I��f}߈zV��Il�b޺�/��&���!yW|*3�<��&&H��ط�j��ҁqe�KS"�Wd������9�!k�.OJ
��/�!J@"����	����o��X/��Ğ?%��!Q�Y�.q�nZzX�<�,��K�fB�%�jh�Ё��)L��q�7C��O{TT��@]X62�U,�B%K-�d��S�}�&G"�O��ז��4Dj��Amb����x^Y��YTt�`�f0C����\���X��Ɋ�%=���(;��`W�0d���~��@�QGO�6����Q�ὼ@��ڕ��xCݘ�#���#8����3��N�ݐ���Q Ͼ�kw�k�����f�7����Z�d+�QmMP6�>UK��ȔN<4��t=}�1\�Ee���,�숱+�R.���v�'
��!�c�D�_��GrU�ig�2p�����D-�Qa���X崷}1J�U��E<�H����x��$�J)
5eפ*�\���1l+
b��.ŉH���'٦����?I���[��
�F����}͹ ,h�y0�Di��`ܯ��	��@	�hB��H���t�W��G����ͨ)vb�L�g�{X����
s����� Z7+��l�����"Y[
���q��U��v��9t$WU�VQW����}�ٯY�/V��J�NNe�oY��,�jC��u�P������
�q�gk���'�����/x 黾k�]pt�L�ʂ㏨)+�e�$LDc2�X�������)W>&^�����?�y����?L���7k�Ƶg�۝�����/�����0b9��j[�J{�J��yMz��m|t@�z��G�˞T���>�����҂�ܢ���k{W�`d�QF�2���S{�>B�o�?��=�{����g�ˇ~�����-�81����9*��Qeչ��/,=�*�Y�\��F$���0�o
�ܸ8�ޅDm��6�=rX�X�@h�Gb?W�aҕ�,UU.��
��
�V��j	���zh���w��+��#�b��Nѧ�Ѓ�E�^X��싿�Uzz�W2vN��E�������}��*�� P�qx�DUdD�xѰ��H���cI��{GA�j7!P�e(~��[� ��qI�R��v�1�?:
�D���ϣ�**ȼ��zi�fB$ӝ���>,@�)f@��:D}��hk��'.��}��w��^C~���;��� ��}T�!���a�'1�w,4�{_ɫ?��p.Yu�(*X�Ex��Qx�X��tP)�j�V"ͼ�|8-�iIĲE��^C�<�a����`�U��9	�g�>^[�	�ҫ�i�!`Lӥ �#Kg���W�%�y��؅7&D"8VC�}Hρ�Q��uͧ�A�v�V�7�8�u�]O�k�΃zXu%%���qԛlhᣘ;�>'|<t<b&<#�¹��5w�df�ىl6?/�P��_eؗ[
�[�K�������Q;��. zM��U�^\D�l��ᵽQ���$����;L���^c�:>�&���y{�a4%0`
����g��.�,���9&�S��M���佴8�h�}�\P�~�R�~>���GoRaY�{�5��K2�J�)\4 �m�hdS�D�бޤG������������$w�cV�4o�`�g��g~5��K����������{2KQ�y�&�U΂�p(Z������~��#�{�l�n
�.�Wt�C����{������%��~ j]�-��&Ɂ{�	Z��j8��lI�>k��+��J�(�.bN�������݊�8#-�[Uv��3v&���\	"P*S%r��vE(�D�����u|��*�~�%��yɂ*)b��To���G1��C/��0"Aـ���/�%>�ML<lC4�[���$��k���kqR,J/��}>-�t �7:�:����ĺP
��6b8o��X��W 9���͛u�}�G�`�'����{1�a\�����n&�Y�D��AKl�m*�Wx�k�d��p�,��9�x=��%��
3�<���D���r�j"2{��㘎�`�����5�aJ�FS��DjD��[p������P�;�j$m�Ր�,���~�M���-Z�s����@��(�bp�8X�7$v%W/x�=47�H�����5�"��v�$W�0�p�u"�K�S:�<K䳸�v�D��̅U��iذ�7�vr�z\fl$k�EK��� ����@'R�U������vTd32��҄�������U
�Ի���5�b
�'"�/|и��Y�8������H�o�����0n*K����@Ԯ�,��|\hEY�y]DE��E`�2����;TXb�� �(���4�����ԅ��B����u��_M[�a����`�BG��˕
ʴ�	.wI��m��⬸*��]tU$�G�t��玫K�]�W��'^�~8=�&�u"t����)}?k�����bto6x��Μ�
���W8v*Cz�SIqS��}��~l�Е�_����]�@�&����k�p� ��t�v:������|�,!
6�X1rɋ��D�y"��$O󵯭i&�S���>j-d�Wt��sj���$�II�/Ѕ�!�A�-���t�5��(XPPؽ��T㬲���Mi7��A{�� 5(Fl i���DP�CiH�!��D���lސ��/����� �0��5�A�纗��2�=��I>����.����۷�|`��H��e����nj�ť�pA���n�
�z!�7�L�U�+�~sz{�Mט�?�켪�T���{� ���#OL��TZc�Y����p�U��p�����v�Y�xx@���g�@�Wd�"�D�,��6�F<#fJo< N�������sP�q�	SY�c����iI����C��� ڷd�Y��g�-�٠���,&��^�*𧔁�mu��Td��k��<fmBˑM���#��(2�����{���n�*Z��Y|8��+�#LH�UX��9�[�[�%��m�R�c�v�S��G���\�I��K���6 M�������%���F�z���jC�w��T�MN��=���u�����[*�;�6�{��\R�����3ۼ�4[�Jp�#E۳څں�#���
!љ�zƘߔ�����b��#�कY��ռ���m�	�Ӧ��ix&#����P���>��2��x�[U��XzэPl�H�+��{b����)�8��Y�����%C��|�p+޾,�7Y�S�|�ƺ,�uE��
W�nOS����6���%�Z����Z�̪�w�_u)�~?L;��K�
�#�k����T��e�z�|^,I]��cS#�J�7k�{�zlָʽ�k?Wѩ�� �~m���W�ì��5>�9n��'.
�ZV�)2�p%"�"��c�9��҈XT>̒w=��k�������¡Ռ&�&nnX��z�/�{>Y֢k�w��l��5�G�s<ے�(9굂	�K�����ʂ�/��r�1C�~ ���%�89��&*n.q*n;���sPF rU,�ڢ��2{"��Wg��[���d
�Kx���Pթ1��o�����ֿw�Kn�_CdF.�K��d���&��pb����,.\����4�g��M��q�ڝ�p�e�$��S_C$����3��ȥ���Gg��9�� �7M ����>�,$s��V�Z+?V�|!�n�E��]�q��5K�� XFh�s�x,9P�����?�:���ˀo�M{,��%�$�;2��ɶ$�v�7J[�/gG�`�~ҪuQ�7KS����7O��d�$��jE��5l�R0+�r%x��b9�D1[$d�1X��Y�
����/Z'm��z2�  �s��ݧdx���'��>
ҲU�Eq`ۙf�
n�wL��r��_dzSP27�/�} �k�6	��������W��9������6*?��e�S�J�D����y����٥7~���n߲|(�!ΆjSyVg�P��X�M֛��q��X�p�ݗ�u��y�C���%GKپt��X8��p���.e����0b�g���n���u'�"��%.��5�zk�փ�w����rM!�Z�ڄ\V�����)�����?��� *�ο4q���m��l8�ۋ��('��s��oH���.Q�k8��g���+mg+:��,?�ԧ~�՝��W[���$�^Y���!~0��{m�C� �~D��b�D���6�|�zġ�O7����hN�8��^& Vu,��e�c�l[>`���r^v��VWܣdKf��k����.[�wac��6��Jl�L�g�5�����s��>��n4Ҕy�m�t��i��9}�i�!���Ј�KJi(���РN��!�X}D��^�*�De�?C-���yjX.mEA(F���؜���_���O[ɳ/-��Hצ�����Z�T�]����4R6,���!����>u���slH +8�o��_�x�TR~���\�[I�{oQwf쬅����CL��C�u6^Ф���v0�dܣ���-�R2�4]����3b	�����F��=���fl�P����� �WoS�o�k��̰��ɔ��DG����B*y�_�%{n]Y��M������ �n��=���)ܘ�q��LP9�XǢ�3:�L|�;Ax��#�W��!�n�rH�̈K���C�n�RP[�����b\y�Abi���t7��a�0V{���迌��Γsp�k<=%�B����G8h�X������o���g묪�N�<d^�_ǑO��~�����@��	 F/w
X�X�Y�����Hx�	�A���1jE���ɐ/��pL�;/��js�Og�g�3�����`���*[���֤� i6 H�h���k?< juHr{�U�8&���$FwL��hh
d�Z*�ꏦĪ��`�eG߀�������UNBpҤlk�@aRw���-����H����R�7ۥ��$�4��>��i�������j��C7�(?������>죾 �I�^(۠t� �dESH�to:�R��@�?5p��;/���F\�VV��|a�a���v���t��b	�S�[�]q�kg�����E����W��F�{��b4�L�{|���W�5��2=m�͙6� ���x���\N�T�6�A���y9��.��D��m����
)���=���`6�"á`��@�lޥ�B�)�Xӈ�*�H��r�_YZja�L���t-�e-���-�QHtO(�w'��[�Ś6%nY���e�QE��ܺB��ΐ+��J���G�#�:�5����H��>`I_�SԳ)C8ͣ��Q�]wQ0C#.����{��|ӹQ\�?�GP��UZ����ݴ���5�d��7����ey�y�5�R$�4c��]�0�m߇���������]���
�X�%r���`	$��nB�C��r��K�M��u+�"�/���/��Ղx�rs�tl��/�Q�e�0u�M#n��Wb7�>�����f�dl5�-�.��w�n*��(��sM����z PY�ö�?_ h���o��іB8pa)djL�o$�!
�t�"���5��F���z��z�x"�r�;3��?GV<"�.���ml��=�o�ҝY�wR�j����W�C����4� J�5~��z��8��G��)2��Mu��J�7�-RV�@�d���*�f�ʚL!Vi�G���f*̪���e\�}�B84��[�/�|@�h]�vG���V�(ɽO�-s�����g��~ƙ;�,��eKqxVS���)��9�<Æ�rĥ��29����or?t�7*RSZd�t/O��[l�~�ޣ�2�?t�9�h���;7�e�)i�Y���(��.8�S�o����կW�� �ѥ6*�0Ǵ����aIp�l ��E]Y�K7���q��Whr�����2ȗ�^�<�v�w���^��O��R�-�Fo�?h�޿��vK�[˟j���#�S��K[����m�a�
�H�:� �*K��w��OtHbl�B3[���B'F�'�X��v����IK���tYb��`H��.��L��2ۙ��N�1n'/���49�h&/~�v: � �����e���Y�C ����8��~�Y�|�E$�� �7��Oƒ�?�1x�*kνW�̅�b����[���^�Rm�;���^hWv�$�^����bqwe��y�<aM���EB�Lp�gV��ژ%��:�"i_򍗢3$�S!��p��CXu)8"-PzXp�l�T0sf����ʪ��M�䳇�
@���0u,BYN"�!�m�����Rl��ةt�9m���b���w�&�Ȩl\�*Y�* ���� �d����DI1 V���d��
���,c�e��;f��zk����޶��~t:�Q&Ӟ'n�=�(��z�u�SHk�I���9 ƺ	�v��m����B���aL�΂	Pe{�HA���u�b�y�7[��vO��ʝ��Ʋ��MW�V�4�M5��t�5ڌ��;�%h����NVG��
Y�$� g�Tj1�+�� ԕ;��0����ד����2��h"�^3>��bf�w4��1�S �:�1p�h�\��Kv�#C�9�H�\�(�-qˬ&S�8�?7�6��:.v����`�n�R&FZ�a!�aƐt�[��C�H�w�^��=�'�y�7���E��D6wPTŗ%��
��27����M̄�M�l��F\P�t������֕"N�84�u/�2vy��?�g%6t~�&�<���h��S�3p�K���k.-e��#�ױq`�3t�;����E5�N�
NUs��m*����J�3T�*/ुg���JC�@�8���O�`�����[�,U�K5ۧ�*NU皕@�y�sxN �j����XY�﹥��յr��%�Y(8
�j���ݹ�钷�B���$z��I�L}S��4O��[�L���)	�,�X6G��=����$�Ÿ��sb=Jo
^�Y�)Hww䐘bj#1h��ୄl���1ݓ�� <ZO�w��7O�8.��}9�� 4��AΪ���J��öf+��x�$9�y�8���YS�U��������Fu�0Qډ�H�p�s�t�6��v.4h�"�]�hQ�{��Ji�|��HdrJ�Ӵ27��z�����|:j�x_�^��;L5���}Ո��I����0�8���qGC�j� Yw���_���`��"�l�q~��,ʡ�^ړ&Q��G&��2$d�̷�(�/8-�Qhb ���xO��t����xFU5Y���?7�a÷I�A�~n��g.��L�rH���Om&C��QwQT���Y��h�>�ʱ
��g�?3���wb�E@�ߴ��ݺn�wóJG�������u�S�j	���>~j'��]�f��-��"X�ѭ��W�~��q8�e����u��BjH�<<��4` ����H�y�˃�m�\y��g�7a�U/؁�d�c(:O�b�%�|���eV���[���Ew0���W ��Ɨ1~��B_o+��v��p��z (gux��Z�>,��f<`�,�1� <p���Ǉ���Z���.X
=�GF-�#�ߴ(�SqR��O��qB�k�`���T؆�i`���(����Dg�a��s�}x?��I�Yr�����(����ŕ���\��z ���#�V������}$��u���/ ��J9R�$z5����1�P��F���^�;�Z�'�ڞ'1���O��\�Bg�ƣ�CG����N�jr�N��?����w��s��&@ �P�I�l礼�/��k4�F=�8t͵���i���\��wSi��5��?��@\c��0H|in4�����ޡ�ș"'>�����e�a{�MB�μ���|*�L��ި,aN�aܶ��Yz|�ntlh��1�;�8�����-i ϔE�&���:���@F�����D�^5�_=lN8�U=�1�i��r��'S���u������I�݇Am��Љ��6̎����1d����#�ޱ0�p�Cٺ���F�M4Oƥ�:��������~Ę�;*��ͶL�q<H�`�{ȧ��קWP��5�H͠�:(��ӛ����ե��%z���.z���N�Ɣ��� T����^Rs��KK�w���ba��E�4e<�^�|�b(X�U(�?����W#�]0���1��CnvC�A&�E
��Y�Z2�H�ѡ�>�ǲR�(-�YL�*�;�Y���X��i��^�����2���Χ�U;z۷Ylgzڂ!x����Lф,��o�� ��o���o��۩����9��;�J$��أ>P�J�+$.�F�!r�T�r��P�{��b�~h�FP��o�F���l�_��E�<��� l\�E=G��䚺����k���i̎��P�ՔX(���֚X�\�d�_�X
�]zg�x�i�p }�V?�7o�,���t?SG�l��v
��o���3�ڹ��h"���@m)|�H��K�cx�� ���l�k��}C������7l��[ي����)N���@ f�۫�R�W	����?��*"�$�����ʂ�0���?����:$�b��7i�D�c�7"�m
��l���,�����{����T�h4�_�I_h����%<`�V):������K�:���+�� �V�n�^R����h�i�P���W
�R�d��e����1� O�{^�d"X$J쨂F��0[�~Ц��O}�� ��^�Fױ�|�J�ᕎ�I�r7�2�c&tؘ ܻP����3���SE��Ek�p�n����g���`��	(7�Ͽ=X6��ހ�br��h-���u��Z<�B��~��	D*��\�h4�W��$�{�z5�/޵DvU&��s�R�u
���z�z%���{˚��~Ux�&r�7f"eޖ��B_W��N%���2<$�Y_���] ��zb:�/��9�O�D�c;ONڶ5�e�9/>*����"ȭ��������˒���#��,r;��E/�$(ϴ�_�l�x\�}��e"?R�Zs�,�?@��}n*��C�z���a{�	*��k	�J�� ��䊫�5Z@�~�n.�߳[thr�����0�b�	f6��! �?�~��B����l��*���m�k�
��4`c�P9�%NH�C�$R��z�ǣ#��D#�����R:{��R�\����(;/i!�d��ނ��.��(T(^k�����A��Xn��OK�O@�',~�_DTˉ�R����Z�9�B��*���#З�!���b�d�@<�����a~��Q�a����-��抃_h� ��_z�����{��W�򕅠����0zY���Q�C�����Ҝ)��}�����70	����O�I���P;]@j�^Vd'��'z(��P����*�7���d�w�B��f)w'dO������)9k�R�4[M+����\�#��Q3k�R�FJ&�u�AfI���I#���y�}��0�l������P|#�at;�+�|p ~W�
d([?���T���������Q���P��~EH-O
P{+�#����]l����U�=�n����e���ܴ?�؅Jĸ
�ya�?�,��i��
«�	�3�^�Յ���"N-щ/7�V��Q=�ŭ�ۜ�+����,����#n+��'P=��:��_YT|q;�p�*�x��&�܃<�G���J��X���*��5.�0��u�j��,�K�p�Ƭd��DtIg�|���VO^y�7:�?�	v�-�����m� Q��'�S��x�d��`y}l�F�q�[��.���ש��Ν��
g��B��). ���;m�x�\�֦��sg�2��tN���Mm(w�#T`�2hG`O�r���O�dO�˱x?�]v�
�[F�¡�	��vǕ��>y����Ǥe�_a9A�{��X�	O�}��'d�R��1���ÿ�5�T(_�XBٽ_
�����3u�I�)����W�c����-�]P�p�����n^�چ�"3VJ�kQ�`�}ۍ�᜸ŴU�i3����+�V��v�����{�*5g��eb}�+	�S�/uQ��#������	����|������ޖ�iۉ�6b��ede�0{�����y����j�ɏ5���Ad�,�q�!�)����`c��qA~Ћp#�*8I-�O�����+ p=p�!=�lMC@T���0��C���8�Lk���A9��XJ�:/�P��'���+x�t�y4g*:l�v� ���[���!A�<4tΙ]�z~Q=e|ͼ^�{�D�X�h:����b3f�Tf�d�v�ꒆ[�T�43���䷍�΁����H�?��Vg��Q�9f����uO�:Í&���&��!���#~�n�!i�3�Z�����:4��\�`=��W�0a��ҁ����i�޷���X`ټ>���~N� �R.	�O��#�K-#-�	��h��&Lr��:y?8>x1�K��[m٘�Iꦋ�1�᰼��OG*�/<���c���3��h7Nϖ����e�Q�8��z�+�,��Vd��$i���@h�uosO:~�=���xJ���XA���%�6�����Rc�|P��b,8�S'V�F�+2�ł�Jf��tR�"?x�� ��^��0��4!ɢa"rW�Bza�W�|ѫe��\�GA�%q�$ȶݽ1z3ɱ��m|2��� �Zf�@�`��OFn���c0�+Î�A����믻u�;t��A���_ǟ\�ʢ�Z��z�KK=�m�.ǣ�{h���md�^�PY��qǘ���fo�$ٍA+�Q���?�P(���MWq��;�����q];�\��c��{�N�ta+�<J ����	���,���|�x��ɲoC~^Zˁz�%ɽU���>2fz�obvúD���R�I���^Rt<��7��zn~+�S�<A�}�!-q"���#$ IH�`О%o�I���c"k�-����+TO��)�@�6���H\t�[s,$8 ��e��;&��K^H0�IW3��!����MtCr��w�kUr�pc'��hJ��/̍O`	* Y�=�Y�r�t����ND�'�x��a��p��,Ѯr����;k���VD��7Χ/�	�\a͔UP��~��6]"M��9Ĥ�.mg?�iA�u���s>�n��*�MBMo�u��Sd�T�]�N�th桼�	2k�ZCX�!��\�
�����xG�`�J����^��>K��\nh�i�Q`�3�Cԫ��ڊ��b�?�H��� �J��39��y�1]�dd����M������	nX�������zUKH�Qm�����	��l���X:�%�'���՛q�l����?�ʺ�tF�ha�ј.��˘��IC�_G��Ə��}4�vc�4cbuQca�aLI���7���N8�I�ߘ��*T8����횷Tt˟�4m�e� 
OM�)�!�U�x6�52�O,��%���@|x=s}7*�˝����w\�7'���%3t	�̏:߉p���`B���΁�`�98۝�b�IQ�\6R��vəT/Ԩ�UC7a`e�<:Ø����R�h�"+�tPf�/���+UWd�9��H���c@���Uҏ��h<�I��v�������'�h�.SyAS��`�k��LC�`oI�4/�8K1�X����er�Ү���}>�.���kwdŎ˛�>�o�����u���G��u_�^�{�k��x��`:f�w�oj�Q�C#|�J�"��OK���Q�m|�4�,#��P v���h�9L�0N_o8#�'My���O���Q �a�`
3jr�������Q�\Nc�.#��p�89��GW[S(xp��U��mXP&��"Qx��2���#��	,p5]Y�7�f�����t�Tf �>�j�qv��i��*e$0��<�b]���y'�ӱ��Y�,�>�g6�n����^�'�{_E���߱�6ڈN��:�{0fiq�V��c���T-�+�ūZ1)�	��b�mXePSV\F))�&۶�t�G�A���%�������!����)����]`��,�#U�qjB�lfS~ÏxC|i%g�xz{��L̨^s��h�ʎl��F���n�)�l���Xx� ���Q�|�1%-��T� s�.2���^�/4(6�p��D�0�P�nT���q��n
�����y���1ǝ����� 6�RAصW�����l�Y�~�hje�O�<Rn��\������{�x�%�?�u�W�p�KGQ��Yv=�?�2&�fn�`�E�9R��!N���?ύۅ_�u6�5NJ��u1��D3�>�P��F�#�j���=sݴYf
�`)v�S�[T�iԜӴv�S�׽C���jF%_���x��`IoH	�+�o ����S�0*�)m�FPZ���̿�Kg�Yf�^v�Gɟ�]�S�C�F�n��t���%(gD�X��o�[9��q�l�f��U�J�z��w7�ӕ���Sa��(�)��f�
fZ���n��6�>�~K0̰��۹��6u-���h�ꪊ}J�W�6�g���?n��BE+�%���z�d4�_�"*ɓ��yO,�Dd�s^�c(�]����㢞U�X�c�9L4�@���O5�;pF,7�0��6>b�.�͎%��vT�.4L/�}?2��7�n�(��>~,j�`͌p!WO+��!�p�tlyJl7�b�]Q/�Yi����2\���*$>��VԴ��2��yӭ��b��5�_�#;{Y�=��p�p&W�/+t�'&�u�Gi�"�֞��;�6��'��r��N�]4�or��[�Ж��"�p\�u�ql'	;���f�F�����<{}��uu�7�d{�s��eC��ӻ�t*��4���ʙ�(c{ھ
?��fIQ�$���DPL����`L�l�*9_l���N����E��k �#�n"���yJ@Q�=FM�'L�7 ��o[}���N��6�؃R� r�$��u���Y(:u?��@��=�rd%ݪ��Eg���A����9���;�� 8�2v�K�v�]�Վ0����O=EkW�kI$b�d�RE����΁f"�I�ON��2���ѩ@%A�M��X�S6���;O�r�S�{ �f���%daP}��S��պr�lښkn�Wҏ��)~u���{�=%�HH�v c�_;|ĥ��I�V���w4`@�b��x"��Z=\�o�;՚Jka�e�T�{_)��sKOI\qң׬֋��^�T&� ����s�;-�����p�ӆ��7���&��O<�k�0��v�J���&�Eixe���������d�"y��S�
�4�7��W����e�H�|b��}�����Ν��%��E���j<�T��k���HF⸵i�"�>޿�3�g���`��B����7��X��uѽ
Œl�_�*��
]���!V:.�V8W�0�������6'��xAk�Y� ���0�i�4�b�����Α{<Vj���^��1I1���t��*3qP_�����M�r]F���B8�������4�\�+���H�W���R�2��(dԕ����d����H]3A����4��NoQ�^�ПH9��H��k>,��>��+P�(|&�a8��ރW@((�A��}���ᐩ��cʎh���n�G���u-�Y����s�����;�'��w	Ǎ?c�o�:���XK�?uz��/�PW��k>\��j:|#�P#n�S2�^�0,�r�q��f�f8��7cX���=��J�������ɓGDM�������ЋQ�>�V�AosjGq�@���\�韎�;�����{7h)5�k��Pgf�Z��v�X0K�V��RK��4�>�P<���v
VD����S��4�^�s���{��&�����{�&�8����!6y7�l���K#���rDkr�3_N鋐h����E�� �c����7���=_���S!ѫ�Iq�>�l�:I�>U"	�E �Iغ?�]�.��r*���~罸_Pۻ��D��N.̆�{Ju�@������i6�%�/�f>�x�練�y���2Uq%���?����'�DU'�0���c�(�4�|H�9}T����ITb��r������w��J�I���I�&����r�@?��I�=Z��>Jy�rW���b�=�R1��a�����I&_n���F{��m
D���,>yZ
�������~����/�Ťi�%�~�j��7���	T�"����֪�R�8s��Fz�CO�.�#��bq
Ws�;&��gpN�~��`��"�\��,�t*�c��|�J�P���Uo0�Ns�z�ܼ��<~K+��6g!43�ۣ�\J�{`���ג��X9)��`/	��J�iਕIջ�M7�'`��k]H���Y���P��?^�L��h���i'�K}xHb�/��,X���U�D�w�C��Nם7's���_ޘ�b��29�\�r+�ɏJw�t��Q:���
ϭ>'TY���A��F��^|�!^\�ʫ��X�W��5����.w���sǡt�#8��7fOK�	��BH[y�#�K�Ȝ��u�jh�	��5	]���ja�\f�L�c3fm�U�����!Li>%9�a���"���F���Z���S���ND�Hn4s̥���I}�z� ���!�B�-47�Qu���_��η	L=�Y����j��k8���#�+�O�����	Lhl�n5�#���R K���d��ڋ�_:�
@Ш-�,����;[�t���1���(C�o�xqA���v�=�DVԩ��Y���ÙVն1ǉ�x��G�b1i�2�jg�]�^Θ̫����^����y����VP�ҋ���!Xh�T%:�+�!M��|c�j��2zxC,	̲�%�w�&$�C~��jm�m�D,#���	��Ȫ[�e�X�
�I	�'��C����L@��[1��d����@y��~�	x.�[�v�A���Nʷi�v��׀�6��!��ź֡�8�G����Bz9���6��q���hk�8G��kD-�qD_%F3�?���$�w�qv��*5���F�#gե

���o6n�ۓ�����B�So(�c���9�-��w(;h�:��}��8�MyK�n',=(�3��a�W#�2���t'�~ {���%�t.�\����6'��=xMS�B��i��>xGP7�簣�6��G���6\��s"`�tE8�?��{����pڝ%3�6�#Į�����PJ�=	 ��D*�PqM���`pk����y��B^(�S$����J��G�-�m����\r�F��2`� SHqlթ�KtX���[Խ�ϳ2qa�w �^���}�\Q~�)Tj�u?L�.4���� �;<�(�B�2���-,�`H�5��O��/7j@���������R?ȭ*L�c��Y��<���
"T
�X��޾a(��{��eO�]B{�Y�,�ߵ1m {��ݎ�um*����H�	4�@1�y |����Ձ4*��_��H�k������?�e�URm�àZIC��|fl_��0��6�������.���2��/�|�\<L�׊n����������%M�Bn '��揃�-�C�RU�����t�P@Fa2#a^D�-�S����8q�U�ԑ�d�#i>�:vf9 ���lU�c�B>W`7e����K���|]u'��7:ֱ�y�vF�4��_��ֳ���������}D����w��//��&0�3�a�$��`��V�
� �[���Ɛ>�Z�#�͒琗JǾ'���xěx�f���BC�=@���>� !Z�p!����pE̮n￱�s�4��rKH��BZ\�O00�R���(�N��7�qIji'V�$�g3�F>�����P�ˉ��t���3�)Qs�[9�\��T����F��kKQ;�8���I���m�(��Z�{YL�-���/�M�:��Y��Dȧjt����6���I	����&����D� �J*}p��b�Y�í��R���s:~� >��A0�i؆#�PY�t��HGG Ȇ��]Rs����EV�=�N�^��P��h�)%�8X�­s���%yb�H3��w��W�Dt~����V6F?��ԛ��\��C=���K�)��$[&s�pJ�L<7.����/
k&�ҳ�1k�,Y�tj��<�Wa{�]↹`}>��Ly�*�4�f�U����� S���>��+�i��rr��㉚�/�IaZb[E�'���j��s�öHBm�v��!:sT�2�.���0���|y�v3�yӁ��tS�W��vs��{!����Ɩ�|� �������z�N�ni_�<���>�e� b2��e�\~ұ��.���v+2����GR���آl���J=�@�5��c!k�:->����2,��W"ZY5n�Vz ���;�� ���~I�F�ݚ]��5��s��y��� ���Cp��/�ݷ���	a�OӺ�y�5U3��/�jZ��J��C͉�4��R�	!�I	���7yd^��5k�&�	^�6�Gm�C�U�d�ұ�P�"P�+�J��ޕ�