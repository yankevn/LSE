��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U���K��)`�c����P�k����C����׻�U�(`�-�B��H�0C���)Ck�i�ο>mY���w@�^���G_�_gJ�t��$�\g�L��Һ��st��J�R=Ϻǅ��S�5��E�2(�T�!�����;��
f��W�(�G*۪b�r���@�!�3��B�{q��8k�*/��7���7g|�C����4���<~o��pE�>�B/������&]�C��A��:X�*<����\��|<7��0\ʅ�f;��uqu��}��N���K��dF�Z� �mև��^����k_g�D���Ar`{Φ�P���^��T�N��~h�={�r�L[4t'�fT�V>��{�/�	�XN�������-7���z�+�zq��ߔ���:v�/�7D�*�V�!���E}��W�2N��K	] T���1��V��m~��&CTНE�M�8{E��=L�]�<]�P���RК�u8���h�.uFKk�=)x7��7���5�Fie<������A�:-����竡���O���h\�<��A�8��5�����<���	L�̨�u�E������n �՜u���ct���!�3���� �N�)�Q�8G0e�C_�(_��Xu*A�#nG���phP�B5lG�\7O���ON��:��_��aU{��ٚ1�)p#N��: �@�h�H��>��Ww�~���q����o��}���6C����{�ap^�3�A�[��Է�W��������(M/v[�5ҫ�Kl�~��ʯ%�x���k�
i̈́���4��\���蠛� Z�Z��x�8œ@}�%�,�_ʣQ*{)4rx��Qຏ;IH0��>��Գ����/r~Y�[�rN��W?����h�����o!l�Z�1(�|y��w�%�ؓ�<�,�7%���MVcXe�!"@V��ap�&�I1h|�6M���5��n���o���i��h;S�8Udw��<�Su�Wרb1L�2����:<�A���mu�����K;״�q�w�>���.��^ZR�f�.�ɖæ���>��Xr�_4y�X7�F�P�Qؒ�	��Mg���S�ܯ��L�9���)�8#�tV�������@�������Ƅ<O�Es��E~C���ˀC=�/Mq7"���t@Nn����m �f�ts�\2�GO��P�UuDĬ,�
Ў5{��P&Ղ�Z5�Q�8�a���xdr}X�*�[��Z�0V���?����.%��wM<
���86�ڜ����L�ָ�@���z�+E����A7�y�*�Ǌ�{�|��mS��Y�]�`k]�Q�}YtC,L3��V���)n�7������t����.D��&ޖ�ah���*�xj�-e�J$�xr��;�8�U	뤥�\���ʸ��z9�^k�����0��LҾ����	ʽ+^z���n��Hy��o+��6~cyi�:���S�
S��r{��#��M���HR�ƕm@U:�E�F,E���W]�]6��෰�����?yQ�F�;�Pإ�e/h���CfsO9QҐ�t�	Ǯ�e��P����}rY!����hZ��A�?�����5B|R=�f���E��V�d8TmɛK۴Psw�\��H�RyB����[�a=h��B��c�;p��`:k��U�Ӝ�ty��0U
j����2ݪN�3��p������~>�P>q�5m��K�������^[N�R,4a������gu�]��{ٷ+p�UE�.٥�h�"7.q1ȉ�	�@O=I�3��O��|$����[�UZ<y�������X�Y���A��Veʉc�<�J��Շ���e��������o��}��J�-	�,?-�=���t4��������B<�:4(��uLJ����n���.��!k(So��)�9�x�O�a8���u�
���.~����j�.�zhֱ�ڊ�-A�A�kJ����@co	�T���j������~A8���'!B��cKQ��w�5��oT��g���u���2z%���[������g���
f��2Sz��w}��Lc+
R5�C�9�Q���L=�N��+���2y�Z�S�u�m�V9+t���#�@�]E�_���]���@:$ӂ�!j�?�����@ �_������ ����Y����&��8R�|{e2�0���  m���}g��E&	�%�C�U�o����v t(�i�|�/S֪�|-1��N6�k��l��>I3W��T��k]��B(S�������Wt�P=H�gdn�q��( x��
>u��m�P?�D<x��@��^����g|����՘-p*�5y��Wn�y8�WzL�=�`�x���ڣq��Oc~�R�q�g����E^�s�ps������f��X}���|=w��4ki�a �:���y���W�gG���:z�1�6ȥP�ΥZ�Tcg�<1����ξ
&�~�˹H�O��dm]j�z�aT�햭uTΐ���/�;N.�@O=��{s�6;��(hX���vB�i�z]v ;�߿��F�R�>����n�s|t�7{���JAI��p!=���]� ��v@(ݕ���%R�4������]4$����U5αZZ�
	��������q�q��M��v$OH�r�!tzdg�y���MH�����������Oo�^�`����j/��*؃�G5t�g7b��(%�����.�db�^���[�l,�vd�	N=?,o^td�S@E��O�s��̼}�/Y��f��I��������*��E�NqŁ/��2������f���}�I	�L9�?�	Q��fU4�4>�����~��U��?x"�,.__�S���Ԣ_b`�[����4u��NC����Z�)FpTԶ>�#��D �N&x<b�.�2��u�t����+֠�!L���ʯ�$���I�h$�x�_J��iy �H��u˼��;��-#�i&����]m�E��C�,t\�(�
�.������f^X1���)w��_�v�.;2�s  1��u�s<~�&��{���\�3�Ri�2�8���P��iQ�4�� aj���r�Ҳ�Lq����^H��pL��a�!Z�x��c�n2�b��� {����=um:�S���hAV)�^�1$����G��u�kn�I�I�y�2X��.�k�dc-G�n!J���6��)ɾ��0:9��x�\��f����Ay�ɓ�L��c�x1�Q�[(�);�-�)���;�x���yT�y���Lm�I�������^S�ؿ�����Nx-w�H��L@Y����ȩ�B��7���}U�Z-�8M��gs���b]���e�x���g��0���&��4r�c�
iD��djZ��Aސ�ɓ趞܏o�^�F��U~!������=ג�yUq>Hz$��Z+T�m\FN<�m�2 d<�דa�lq6�-��d�GZ����̡�[��#a������'�/�Tk�-����vp94SL��:~s��Q�@�#��=`�1zKɷ���a�h|R���{����@����c��t�r�4����	Iho��g�4�F:$ٝY��vK�;�\!}B.N��b�<~6o'6�}v�'��PJ�B��>�ٙs聯��y��hY(��SN�@�/����}�ᲆ��M(%��p������\��m�c�>k��uDR�%��鶦l�ς;~={+s������.��g��Rk����y�#��Tn���Cr�����ܸҎ���_ņǨ^6�
�t�n�֖[��F�Q.��@�?���9]![&C�Vp�T���v�~�mm�SX
�1DO����	�\��kz X�\,S7M>��_C0S�}ξ�ԉ�$�P#�)�*%:��K���јDg � N4 ��|�eЏ��r���d��>EIT�{Չ��:��{b���O�'f�<�,�IM���p�9M7�=�Ys�Q>�S._�@��w�� �]H��֋6�.�;�}�8��{��ɸm)�ё�E5π]L����K� ��z���$���.��p#��E�)���Ԟ#ZC��~8�ٓ�Z5v�x"�Yx[�_��?�y�|�	˄�G�y9��v�Qə�k�0���6����ɵ��2�N�O�����܎����[��4	�b�#�bA�X"ʄ�s��ek�	�[ZNDn�_��!d���v�~�c��n�"���*�W+ .{�5`��B94	޽�}�brQYxb�\�l7ݯ��wT;S.�0�3mOf��ü4��0�b��s���c����(��#o��0Cg�л�k���Fy���G�<fD���$�S����Ye8u�/����\��"ɟ�X�(*�D$ֈ�i�L��c�D���ѽ+wtE�<����S3@���Ku���T������	ā�$�T�0ɹ�x�\���4��+lIC��At�e���u�&��*��38FI.$��T��rS�<�`Y�y�(E\�/����^O�kVF��A2e�
�%�Y#'0G�`Q��}��y��m���1�G ���S��Ӫ��w��vk��$Q���f�-�n�AϽ�`���:L!(=z�nZޖ�%�S)��Q���^A�L�8&?؟��ۈ�ފz��%���?r��%+��	I$�.'Br��v�MPng2�՚}O�"q�U����>>ʻ�Dv�����JIu+i�OMwI��< ����<M��1w�nV]!��j���0ȫ9Mq�Z�ӔVv��fp�)�WR��ǅ�۬�Л��i�tX.V��C�������~m��*�Q�"��dʒg��R  ����(K����5d�ߏg�� 
�:q��S�r�/�.S5I ��U����w��ipG���J��W�Ի�����gr���¨ʞ���rj����> ��m��8�>�^OD���y�^ڹl�u�PC+�6M�y��%�)���l���R͝)�;�:�����fd�2ځ�E���(_��
�� ,j������%G���pLAح
X;H?U{-
TU�¾�dꝠ$sY/{����Mt�����Y�S�/��"B�g��w<;��i��-�ī��1��S[�e&W	�c��)�3����֑����n,GMl���v礔�^���4���69�/����tn��dy��X��9O}^V���{0$ẖ9�ژ��e����׈��n�S��pw8g)�ZPi*&�ګH|zi����Ν�P��"��������j��S4O�2@ûq�V�}����6�m�Վ�|<�~G;	_0M���#�<ό��A�i�q]�`̪�J���֘v�����a$�ٱm�1��x��]ρ
�#3 /c�~�m��F-�ٯ�`���y�9�hX3�A����P*T�?y_/�En�ƣ���Ih ��
�$�5j���g��""㴸:�G�<�WTA�S�(�>}�Wx*yχ�"x�2�<7
wnf���+딉��K-8�hiy"!Cr����{�����w�<"h�>�V͟�3eC�	�3�Ę[%�[��������S��<�5&
-	|�i��g(����0�c��r�^؝���Y����O�?�`&�{���y�|���� �:��(�� P�y�k�*�W�Q)�ǽ��Y���m�{k��6+�̴6x���Cъ��k��
�a&���Nύ'���z��?�lܙ�!��]~�8r�~�D�h��@D0*h{��M�}=L�0U���ڨw���M{����M~�8%s���3�>Jk��}Dv�|'����m�j~��.���_���E���Io��&������$sL۸4�2U"��XS2<ũźE�2���V���Dyr�_��c�6<�Ne
��*H�#7"EF�H���mI�*�4��+8ûcӼ��}����>�N�%��|1#̞p_U��&�V 搈�#*wn��rn���5!l>.D���-�x��~u��rj�����Lx�Q48+��D	l���MTo���i�`��uYyZ���d~��"��F��Dm�0/�2��I��$��$��~���M���|�`��ʺֱ�<�1����}�����4XYQ.�pȮylu�����x�gʹ떀r�����7'�Xʋ�W�\&yr)E�L�a��E�-A*Ug�]��$q�"��Mj��z��(�1��5�Kp��o�^V�>%h��=a��
�&cə��ێ(]G򮘔L�d�t��n�Â� ��+���ൗ6�����,QZ��Te'd w\.A#��V��?���!҉��(��� 8���̭D�1%��19�O�5�?��?2|��(�G뻣�])|�#<�P����z��7aG*0[>��Z�À��co������&�f�g=7�p��N���0��8➔��'�7���@�C�k�x-ω���c<�w�eI�ʋL�yxjC,���?x� �U�_F��f��~Ζ��	;h1K+�WT%�O��m?HHN+�#?$�oT��N���L�<�E�i�xܬ���L���;�IP�����b��S���3������wu��5�ݘ؀�^GJ�\ىV^�PuX�!ʁ�JM�4�A ̾��)�i�ewNA�k~���rO�|�������U>F�hə��� ��TE���)�o�wRiJZb�W-�c֟{k���X͒L�XD��^����>�'�@�`y�e�mxe���:X#���ハ}q#_�!�ͽOȁ���7h9�;���5�@6����N���i�|�ܞ�KŃ S�f�Q��-�B1��'�� �ý�k�j�QW*�U�(i�sXڰ4�庆�Z�y�D8 I�N�~�FQ0CZ�r�SUuB�>���6{��zHmZr|?V�f.,z�W��ȇ��M�3`����9	ï��P�L��Mq���������@J*b�tJ�+B4���5����lz�+�-�*n;����	f��Џ�T���}����ɒB�Z�Y�QPm�࿥L�,w�KS�
p�u(�ԑ�%ס��3��f|�=:���i�"\�,�,~��s��d��漋
EZy�ou���RТcM�	N"�k*I�5Q	���L�n�I���j�7��:S�G�E��֐���m��+���G���l�ӗ�g�@R�	���ؿ?��.-��^�]���V�ճ-	�Cm��d�;_�N��������s��j	p4#g�:��2��}_���n<�	Jk��	jA_���������}/�l(S��:��� t��h^���2����w�j$&m>ɥWA��ߛ�g�v��\���Ԛ�!���9������O�Y���#�Ok1Z3���Q�f{��4�6�#"\��5�	
������m��#�b�-�_d��r��ӕxm¢~J����#�EzU���A:�����fő�ip��
Qb�`�XT�&Y$���if��Q|���_\��P��U�m���a�X>{\�P�$4U�p�qd:��N�a��-��7���S��]�ٱPXwU����a�G�)��xbr�˜�s���?��ɳF�@�ܜ��/P�q�Ǘ�&A�:6L+��X�_�l��&-����޵�*���i�%*�a0)���5�p�LY�/��`�]�/��/+�9�qki;-�Bq
?N�.��Ϝ٦���i�<��ɕ.��I��<O��a��;�IP挜']��u��ѠQ��ǻ�O��D+(p2��r���A�B����rI�=g��xMY�R�
P9����g��O!���tϘMޟ.���������[n_����oZ�[��}@d�ڋjҲ�J6�s��E�(7*x��ǘ��G������:.ڼ�Y�5ic������YUT2�TĢ��Aj%�?�@�8垚/�a�Ħ�J�C4L�A�O���8s�7�2 �v)�hЋ3�FM�ש�Go��v������j�?�a�q>��� r�=�Q�.S�魝�U,45�9|�N�4�_��?�~U2�?52֢?�j���y���^�D����H@�p��ϧi$߀������CF��@�z����D���%��ݹLS��G��)vB���ݛ��⿪߶��=����x�鄈>��O:��)`6�@�3�GM����j�r��t^K!���}����(	��`g;�^���@�H�|�;�A���s�z��?�S��c�.��K�U�4(�`b�D'���?�=����[�ʄ��[��eK��XMx��u&|�3n
c՗5�x�4����Fj�NXh��8�ދ_�	Х�$��6A� �O���C�
g}`��cL�S�6���OI �n����i����z�<Df�4�u� ���	�;�ci;�Ю����,����6V�ej5�U>oB���3������w�=���3��I~E���Sau;"�5��l[��ʘNwT�	!)��Ge�G�h���q���y�}(���I��Yp^ami
����OL�id�%Q�kQ�.�t`���Uw؍�ԧ�.�)��,&�YY����~�cn����f6Lo�fD�Ib"�
��E��&?�Z�(N�(��j���Z/�J��?��;��5&��U��B��e����79e��٬��
�y8��G�^�o7z�/��~[{����{��o��@e�h�8�7\�p�72�h�h�p6O&�c�b.�9��'��)ֆ2�~��#�0���U|	�[CPW�'^A���u�`��R�B�W�d�etq�Z��uT�Ʉ:�2���oP��ظ*�h/�Gس���鰶���}�i��8�ʚ��m)�����ho].ʑ�60^�!L1djY���=��. �������*5����
C�����2'*+Het����C$�t���ʫ�W���.!/����B��\C��oI4�N��ޤ�x5�u'R��/K�g�%Ŭ_m�R��kX��O*-��˶;r��ԟ(�ȍWi�c[��~���<R�;5�e�4����ey)qt��L�I�����(X_��I��:���C���m�nF��=�2e�ke���&��2���#���y��"�1�����iDpp=U�n99]@wD���$=��������k��h����	�AouW���$hr)1�Ռ[�{zF	U�l:�P�c�L^�~�Ҹ �Ǖd&?3�<󉴤�.}�hm��dzvf�D)~����)����+�o������ǝ��)�)ϝ�W=��Cr����5l\�d���cyiD|P����W�I|oߎ��{���ؘ��])���Q֌,����	,H�8��s����6�Ed���xz�daʍ�&'���q��ADm͆�m�A�]�`�>ݿ�f$C�993(���4���v�y���&>��mM$�|��~��Dd��Ё$�DS�i��Po�Re�������x6�'֞��;�̩�����-Ds ��t&�4�q��Ar�znbm�T�l���8��۹�$��lO�>�2�޼�rP���-�3?��iL�FDCV�ϱ�.ŦD!�3�#j�0q���5 [A�41˜*�?G��S��v ��O�3�Z�LVz���G|U9*�?�,@s��ГB;/aI�53����C/s�%~J�+G>�o�mQ���g���t������ɠ��/ZO�$��|,W���$ �$xI�}k�^	L=�
V�w�CxxԱ>�uq�+�y˭]�4P�./8�aT��	5V�p,�C��>� ��gכ/�Dt�Ӄ#�1�?F��=�^V�HJ�n��	ۛúE%�^6`��Z�'�x! ��E��^��)(h�ū!9�T?�xV�4SY�*˖�H���GA�����#Fo>�$�@���o;cW"�`�Ǳ����HK�����:CN��VC�	�������o���Px̏�1��S���� �/�KR��y����V6A��i|Ra�1>-9}�����oN��:ԕ pp��+HU��!Z����3�kY���'@�숨8��P��A�P؋a��6��8t���;}	f���9eq�'�p�������IY�������xV��WSt�zin��3R4���'�x�w�+�ъ(钕���9�=/����"I������w����"L��ʬgP�0 GU�y��*<`W�v5/��s�DZW��&�%j�	(�%��'0�Z�:"��R&2�B>�H��%5`4
�>!�����H���]���9���V�}�;�E���	ζ�x�s�R�]�kX2�D)$���|ϸ+���H�_	�̸�uȊ��0�?($4���0P�Ӊ��;��"����1�����!� �������h����t�}X�{�����;8��W�B����ka���O �oS�N.��-�����Sp_��+qFj�N_Z!	�\8;Y��Q��7m��s1�����%��D��,Q�-�'l4+2��	� =cGM�j�G��UXu�Ԅ���f����)iN� �~�Bv*#>1�Ƶ�i,d�����32t-.NX�=J'Qj,ࢧ�%�S�Ř��0�i����]B�~�tP<��ѵv���r��o'H��� ���roC;]�jO�3�΀ 4����?���"�=��Z�� t�d� ���k�eˠ�{�Y~���:e��E�"RQK�]������P*y(����D����#_�b!o��u��Y����;� ���QCFe��1�?��:��R���n�E(Za.2���WI-A�`fa����'fD����\,�:V��0�@��jC�Y��������!�51�L��T�����pRo
~f� C�3�f`���C�PПV��*�a{��J��!�o��[ܖyJ���\H�U����ɬ1a���l�߬Z��u!���(��u端�@B��v=�N�!;��� JJ�Ug�zz������m��
�0�3�:��b@"Q����(YT���W~�צ
#3B��	�G L<�O�
��f���t@�r��DXE��|
îE�]�I���9��?�=�+W��슯��?�R��v:�ib�� �b��)S��53�:�D�;S�-��h�>�mL����]��;�` �/��K�m�h�q�ñڲS�1K;P�Ǚ[eyK��u�s��$On�>�k ����k�$�4CDH	G���$�:�9���h5oA�ν�7F/TH��-c8�:���dϓ�g��wT6𳧛��9Tgwo1¬�f����Nn_[�d�����S�^	o�	<<��v)+�T{cY�RM���?;9G�Y'`�`�I�s���bˈ	T�xȧ8�ׁ�����]JG��Ņüq�aL���rG	t:D ����JT.�P"���z��x0^�J�����)�����>�����M1WŲ���늓�X�
Q�CA���my����&��/�g���9��;��[�+�G���� ���]BN����Wm��W�Ǒ�ԛ�^Lrq%��@����y2M7q��בl��$�d��ì;�T��y+��`i����nZ������ca�`G�7�s܄�%�jZW���t����3��,q��'[�(��>=lЫ.bZe�C��Q���M��~	/��3�m%!����4�����{2�G^�yZ����wE(� �����qh�P�`�Od�#�ҭ�%����i��TE2I�d,<H�D�`��GF댫����6�Fʏ
�l��z����|S�ecm��ᓩ/Ol��0��MDe�`P����T����R�c�L������ţm�%���%���#�T�/�_�,�g��ԋt";+]Qa�̒��D����2��F?ػ���5� '�joY����/��7
(Ep�ڝ�Ծ�9?���<lOi�QUl�E7��A|G,��S<a�P��J��cܮ��N���<�6���ɇ��N�B7���30�S
�$-�bw���7�ղ� R�I����|؉Ɋ�r[��׵S��2Ly�p���|(�U����Mm��>}��1^���Yg�����(���cS����!D�M��#�?=Lq\Ȟ�!�]����U*��c�7"�ўڏZ,�! �C*O��;��ű*l5�w ��xʹ�º��j=}m,��^��xP@I��f����`|�n ���iM�e�T�q#_�l���l#7q�u��,���_�k�>mg��^~K��da��̊/�W}�u�R0f&���J�*���N@N���S������W��O&�-d�y����Yފ��z)�"��L�b[�ZR'S	|�G�Ƙh��4g��Q�D}���kϡ�<����kG���5���# Y��P��.�S)����_#���q�I�7� T���HaX�C!�IȞ�����w�����B��x��	e��+��_d(��|�^*t6Z��^��κk����MFm�tK>RQ��o�:h��S���A�.��_	��zJ�H�ids��ѯy���eFY���|FQxY/��e�d0����_�}�.�s}�綥�a��a�e�� �8����wk�W	�^"~�rѓ6H���i-EW�o��^ڻ�8|�Q��ah�&���(���`_�����I�Ҟ��ؚ�[[-;�0r�z莾�e�ӲӃ1���R�Qbη�Aj�P�g�:�A��Ea��E�zo��%�|��x�-v�؁\�HP;�\y�r�b^�<���"�o��j ,�|u�#�$М��Z?u<SR�e{&NKM�J��QX��ax��,���,O�iS�;5y"��"�q���dT���>�[�3�Oȯ�(�G��&�S<#xI���-���u����Ђ'KO����PJ|=@ł�Hi�?ն�	�^�ow�J�%�
r8G|��ۙ�㓓u�J>#��lW�I��(4�����I���H	�p���t�0������+�2������:�����֩���[塴#Q��"�"�:�zT�]���:�E@V�@t��3�OT�s�k�[�I��%��+u��f�@y�HK5��B::���I�-,SI��)h#p$y~����"/��"9r���g��?Mm����"�5����j<�Fc/��o���E8M��Ya�2��)�������hX�I���B�S����W\:����6�ģ�y��=���_3,~�gv�,L���{��T� %��#�n�Wc4�c�)���H�}L���%нb ���T�]vq��'*�ׯA\��z,���O�g͢V�)Y4PN���F�F��k��',����/C-.��ռ޶�����/��ޚ��hG/\;��4��D��`r��+��'�<�S���0]@*�V��M4�l�����k��m"��" �t�֙�*A���=�[�q��(đ��m:�/�v���(m�i=�A/�~S�k3�@Md֪A���n��$]�����7?S6��2�Q�9]�R�ht��+�0n|-�i��6���Xs��+�2�Zr��kL�N�;�A��@�����;���������}
�[-Ź0�^�-�A�(w���R_�`�g���X�?^֔�!��v���<�<<�Ð��.���;����@.S.ݗ�t�*���^ӑ��c�`�V"�#��ͻ��;�4W5��i�����n��矻[�Y'���4 �?=n\���'�q��
���۵֦�^�3-���hz��V710��?Z5��kԉ�Ͱ��q�E2�7u���]jA�� 2K9����A2�ʭ�(���xշR�YF�eYO��U�/�=�@A�I�&Ɣz[����6��Tk��A��j�,?�*����2͓xPPck�щw�\���*f��#j#:�j�$�� �P.Az�jhpۃ�W}*��n1�%�@�t����1~����<�u*�<J� 5QI����Fa��_lS����_P�nY�rR)�*@b-'P6n�TY-N4��9K0�6��P ����}5ަ|V�uk�^���W)���㼝�����Z�3���:��C�׆IZͭo�2,;�0yo���Ϧ�����fD�}�9T �,A�F�vl����m�A�!� �"^�	۹m^�_L�ճ��'P+�+�������	`+05-L���e#􈢹-���=��r� #�::J��e>�dGVK�R�֨� ���GXmHN>֦��e�E�qZHdI�j_��{9RQcA����؜F���8A�ԃ���K��5�spA��6F��;�����0,s��V��
7��L+�=Z�΂n�V �C�2xj�T���`�L�x��6_
�+�L5��U�;7�T��=�w%