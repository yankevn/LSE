��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~ !�s5��<��P��Ҕ�S$�9�%,���2}9���]�?P�~�k�=��[�`��c�ω���M4G�Ц,��w��s��1������Cl��'�N�>D?�� ��Tť&��ަ��k��A>/�����V�v�J%YbN��1��kT�9g�8���הT"W�G>�ɪ\�ŉ���:�/�FFkZ:��<tA�֒@Uϡ�M��f�<�c�bj]\�ґ�ǟ��&h{�������/�Rc��'g�AD!)�,2H5��i����qq�I�2�)�E4D�=/�����w D&!rY���O�W(�o�@�:���=q-��j�u�d���\�E牬!�4{�p�,1+wZ���qZ�>��d`Zyq�;�c����8i!$��*,<a�����>�_�gaw�L+A/����$7iy��� oӊ��[M��FY�+g�.`���[����sZ�I+`���)oi4Z&�Z�k�4KS�`���yT��w ~�܄]snDy�g�D_lmA]Ju��.���^���v�ӷ�S%�%^��ЗF��$����~r�Wd2���D�]?e��oQh�Ƒ��E1�/.H���{6f������!#���TxX-m?�=`���e?v�n�G�"��/�-%4�֍��M�R&��JT�3��.z�.<�J�YN�6�U��/'i$#�x!�?|Jf�3���\)�0��ص�B}c�xUP��$�Xk��1��G�]�~V���؍�,�	���mB�[#����X*����^�����Sm��
ӄ_�x��E�^X��F�!���.8)e���a�e���2�����v����2qy���7����͑U
4�c- �5��`C��t����ֆ���c��%�z��͠��&�5)�(!�Kz`,�O6�6�s�%)B�(׸,�"���V��c��с�i�}����c��c����o�;��*�
8/�h�օQ�UueCU�䵾.Z��� �7F��&�fN����*���*I�3m�-��b��_�R��kۇ}�k�gJsi���5�|��ʮ,�0y�dà0��E�x���R|O��-�
�ъ�%~\�r>{`��I7B�t6FÁo1����VE�	ЂϞ�w����)�Qw�d+��nm�.�ɻ�po����,�`�j�3r�� I<�Ɯ�X�3��S�汷��H%��
m���,Vm��A@|�PZ]X�!�B�p+�ޤ'�4c����f�Y� �?Du�tS�
4�%�Jv �����.�>K�T�T��ȏ�����e������3���R`^��i�C�`D�n#ݐ>��Fh���&F��2���6@����
aG\YQiZf�Wlh1�����DѪHXj�&*���ѡ�o>�����IwO����9��O �7��\��Ie�6��%g<�����/��0O�r�n�c?��)LN��#�����(E�-�!
	�=%ˋOE��@�LJ�Z�q���&0�9�w'��%>.0�X1/s5��C��>��+|s1�J�`��ݵ'��
��	ʆ�4Ğ%�,EV���X�k��7ē8'2���7z_�7S��L£�\K�Vb�&��bK8��!��.��(�v����1�e���R��jF"����Ǎ'��o��u%��i�^8Fh�*�d����f߱���;�f�9�F���k-�197�����"��)���7��7�X��~����Ƥ
�NE�� �{cB�\����=K�q����B`AH�M�a�]�,`O{�EƄ��l�ᐲП#I��:L�-��[�#�l�M]y
��fWv��}���v�vڣ�!2؟L��b��xQ3�bΉ�̓�[2MWr"�	�7+�&]�X�r^+���^�)"6����H����R�[�.�T�����G	��x��}k��.N�F�ҬCg��[�S�I{`�n�>YWU}�(���a7x��{���G�' ́/.�:�];�z~��u�� 8b�kD�:j$N,x.�'�
q-��v���K����>���Y�8�����{�C�����Ng�[؛��]��rN�7^��?�����y.��C/d����x ��bv3׀�T��%k��5M` ԓ%D�7��g�8�
W
����[WK_�	��6 �������<{>}'�1�%�b��2C\� v���h4�?[칝�K|�Z&����G�}����XM�IRy�׽���m��k���;g'��js�UѬ"�Ϡ�נ<������Q��V��➢Y�	:�M�D'����x}���r���;ؐ	�A�F��Gk���4��nא��������4����0b�]Ns�D7����Xϴ �kJ	&>$A�3�$cŷ�핥�p�R������ �C3c��^�"�j8�2}���p�B
��7��D��4�*(��:��m�;#d��	�� z��2-gzɽBۉj\�O�x�
TR���ҭ8���"_��|���*����Ni6���Q�Go��͈��DP�p\�[q;U�M�ܻng��iAc�3 o�nFp��p�ؚ��\�:osWwd��m�DN�$S�M��6�W:����e��8#�<b_>��YSP����oDĥ|�ר�~�#���0�f��凘���i	��+���8�0�5��u��6;n�F�5��%�+pm֕��k��4;�j��)��7���	h�i=�"ı���҆�s�K�˙�,�Z���?���h���1Ŗ6��%e٧��0R�B��뺊Fl�#��� �)8��������d@� ���g��{�~��3|�|����q�t@S�=�-@+â��_M]���ڟ�s8�LC���qp��14�Qܡr��;d�\�Ӟ���v	���P��	qh^Ǜ�̓�{�N9�S�����i��ru����ϖ&3�:�4�}����ĚW�a^�LE�p�}U���*��}�E�|q/�Q{q���>z���%�؂4��FA��z]@��4-RT�V�qv"{��e���raT���@��E(o�i�w狨o^�!p<%ǹ�J�&K�HhZ��F=�����dCO[�G�?8^��ܜ"�m��'�͈�������� ���*ά����SY�<+�{o�O�?d��Lz4��mSihe��M%��fCm��1O��GI�~g�?��:@[���������p������=Vź��{�2�N�$�3���D���ˌ�X4%g4���;KP��d�̇�3��?3�U��b�Ԉ��8��Qww����W}g�ⴣB�*��,ĉ�+N#k�Vjv\B�b2(Ckw8�F��dX�(��7�
��|^[��g��'$'�*_��ho����\}�k���H��k�h�!�A��i������
�#OM��\��E]��vm���|�Z�}5�$ GA^�1w3n�}����-?햙'fiC`3��o\hu�AIX��D��^OT�&�H53P�Xm@�p�i��S�%�UDJ�B�ڵ�]��&�DʞXu�U��ǧ�6��U�$��`�UK���툼�s
�� ����
L?���z���/��ߺ7咚���D�M�����JT���g�5����8����8���&�#촞3���0��� Y�$��s�:�4�Ag�F�D �b#wހ&L���Um�B�����p�蝏<n���^2gNW�}q<g]�}i���B�G\l���V��m��z�r�d�sHQ�ց2Jظ8|����;7��?Y�yj}�����`���.Ⱍ�? ��BO� %���p����&a��S���)?X��$#K�*IV@���;e�kM���v���(35�c�4��N0S$�ܷ�=�����)F�v䛜3����Z�����0�
gW��#n�R��M�a�O}�����y�
���y0�P���+�m#�T��`��
7cq8���+5�����@�$	g`��[�dE&)KPd�~�Ж��a�.�OM��p�"�i�����I��܎Y���X������]���/��D���I��EH�8H�������r����>�M��&��R�g#�/�WB0﫲������סs�"`���5�?�?_�jf�b���W7�N�.�x��K��s�D�����L��}b��Nγ�W�Kiw�����K�nD~�<)�K���z�2�����3N�Z�b3V:S�:�lS-V7f�{��-KK����oĠ�]��٣�
�qK(SIÑ���4��sHU���e�� �5>x/���ʠK�:�.�xW���+��
��s�q�O՛k�^��R~{Եxà���4�����ݨn�0ZGӼ!��]��V1Ӕ$����em=�Hx�9r�@2?v�0�|��8�S<����̯&�a�c���J��/-Z��Q�{0������E�T��
�t�iЯ��2y!�.�9��oGlt 	����"�ctt�q���j�ֿAF̞�=��	����Z[]������aB��[��tR�Y� 4������|7��~�-��-��0p/}5O��G�)R��G�["Q󬇲��G��!��Z�Os���x�;�o�ϛ�!�ιl޾""?��t�N���	kI���~��9M�X|S"����J"�u�	<�G��c&�)�j*vr)G�gb�lg���M�W�j�Y+Ed-Д�Yf�g%.�%�c������n��� �O���#��u�?-���U@�x�M.T�� [����(2����	��J}9$)���lJu$��`��_=���(nal�9��Z�����#M7���xw���d�l�j�E��m4WQ��&'l�mz��`��i||��R���FA$bc�#�Y�?�@�Ӽ�IknrOK����������m�d~wpDF3���..G	#F~��.��%Ѡ� t�,�J�M�r���A\�@�zCl�K�s�5����9���sݶ\吘Sz	I�#�^��!�'�'CeޠL7tQ�a��u�SO�f`��T�����"��T�dv=]�D�\k���Q�5a���C»��q"���=�H�:��@@�`��@M]����bW�/cf��3-��K���
����G����x!����Ⱦ��G���0g$��dI��!��f���xk�d���U�tO��{��Ҁmը9��b���S�W���~�����ഁ.���
p�M4R ;����M}�g��)�\���WJ55SE�Fvy��)1� ���ϧa|o���ȡ�y6T��q�����<�g�*�-0*��͒L�#n�Dzܩ�y��=a�d�D6��5`NT���C�o-b��[�����&��E~2�~�b�
z����T+P
��H��1��� ���
���p�*�.��V��[�<�I��AgX�S��y�!��y����5��g��Ŗ�P/����+Qٿ	"/�WHQNT t��b�6e�D$�]�E�ױ�>K�g��[&<˯Za#e�Y8&�������`ܠ���D��0~��J
��i�:k�]�e��Le���yL�0J���#���G�x�K�.!kt�" ���9'�M@#o~�s{jHz�n�%�;E(��o}Q>²���̞��l�'{0^�l+'r���y���UB�&�"�;�����?D�ʅ\�g��������={��e��96�V��캊�qZ��dr�ھ���w�Z���5t!ݢG�(��o����;
���^�5��"T�I����j�ۘ��W���RZ6/�gVPoi1��'V?H�+�1�cKeЧ2؟�x�^��*C�3ʛ��������E���Z�j+�S�u� ��s�а����L,���F*��Ӥ����t�(6�� ���&Y��,A>���f���h��=�&"��4�뢙�a�;��]����X����f����(�����g>�^�f�r*�^0E���0F��+qϓ6��zm<���z�����Oƻ �<���B�Ü���0��s���y���?�6L�/Ŋ��{h.�["���`����e�Sj)��9W�I�P��\f���4�f9�D]$���<�0��Q5A���=C��|؁&�S��H�!\�t�%|.(��p�Pp�IX0���IĆJ}Yw�����QК��֭�q�0�!�j��4�0.W�6q�R��=�.�يy/���3*�W�CSV&����[OSr:�G\2n�+�Vwa ���f�/	cK։�b;��'��/MƸU��`����ˏ�UӪ(�Mp���/b1)��5��������G��|_\ m�5>J���˙1"���wBaˮC]e�{��	�9��Vj GD����G�.W�YL)~�]Q�&x榺�3$/Vp/�R'�;�	�4C�F܉:B��S{N�pv���[�����Xۣ��y��݃��r��̽��i�|O#\Tp���Sg ��T��"�Qqv���H��(��@{ab�ũ�܉�0 s���$/Ġ���,	Y��k��qv�+�zů݂�F����$W��c>9��A�X�u�����|)I�[�����=/^��K+hyZ(��u��D���d�[ꥹa�3̔�1�S0#��lA��i�<Y$P�W(�|2����)J5t�5��oG4å)	{��Cg�ϑ��H8�\����Ir�c-L���l���0��6�q�r?t+=����zV�/gy����r��D�`��C:Vч.�$��y�q���>߻U
���=�sEޥ䤣.�K��4
�I엝58PR�>'�hz0�r�[Π�-y��E�ے�'qy=�	�⢭�U��@x�fY�>/�:��M0��;
%��c��|�Q	�N�0�ND?$
t<.����VSGڱ��d���HR��l-;:'�w|%l�`�*��r�<%��j�f����!cO=��Mv/�FQh����Ay/���վS�A����#�M�V���~B�=T��&�#�=0��D���y$�I�tu�?��4Y�L/x����|N*>|��]3 W1��u�5d����^&����l<���f��r�W����N��Q����9�n^���N�����Mǀ��k
%�]V����� /2���fL���+׀� ��]�c8�xo��V���U���]б~[� �6N6_J�&	s�,��T(0I������e��=�2��Wǽ��T��\.r���G�%N��]�`�5R�i��5h,����,�wb�XY�ثx��ߎU��~֚E��̂Ώq��{����3��r�K���v���s&���1����L���u��\VA||�!�,���_�oh�Oc�Ŋ� �b�(h7�5G?�-a�
���螗�'������~���}��Ѣ�h�(�Ȇkc%��{EX�D��m��lڶC�i��d����
��;�cKח_,��E@��6���]�����ZX������YgG%�G�p���!���Qߊm`��q�1:����Q�4�P�9�ʧh��]P�:��C��<*�Xs�O�7rv���K>RYI��B���l�bTX�w�66_�[�d2�k9ћ�I�!q���yE�1��� g���<=r�
�i���`=�[�X$9B�x�퍹����?1��P ���x٭�u��N{�������x���χ��y������IbKznnݢ|�u��]��B���v�E�幱3��e<j��m��{���ĺS��c���ny�鈄'����O�^���6���A'��#�zat� r)��#�d3, &�Z7��k_qe���x~
���c��(D�(IU�v�߸���m�1�r���{��� �ÿ�!��+s���k���Z��p>��%2sD�Yޢ�J���\@�\�������G t�Ru��#Y��^X{���s��Z������4��Y���!����+�wie�ȰX���P셜e�eډp �>p��������[���%�t��0��,��	F��҆}M�B��t��X��+���הg?b����}<�ZAr�t[��ҸR��5��S�#�ʺ����R����!� T�Vkr<O��Et��f�=�T.� �*Z.�[�
-1�͸�*��Wi%麗d�x�����=�CM���C���6[�\F2�i`&O' �ci�lB�Pf�+PX�7�L��o�4�!+��a�����B����K�bA��M\�,L�)c����xj���>�����4�+��+�T�>�r�*Wv��lM��Y��9���!����nE�!��x�D2R�mi�ĐoQ��	�� ]��ǖ�G�=�=�I��Ȏ|��g��F�7� �⬲��Z,~ݤc F��5�[��p��G�>�S^�>����� �v���Dʹ̲�VKD9 Xn�U��Qe�6?�;�_}2���Z_eXtKL�m�ǌ)�.�ˤƩձ:	��F���I�ȵ68��Ҭs���/x���+�Zp�<ޠ]�	��K[�������R]�:��DG�*z��K�U۞�7�ψJ��ӈBh���*���`� �&�'p�k��ɘ�@}�jP����ʋ�˭K��3����v���qB���4�����C^�H��hq�4� K��c_X��8��m�?��>^����F~2����@��Dp!�l�we�^��-�7}g�%��=�/ۜR��~�H���-U��sF�Tzih�3���tzq���:l����ar�J:f6ǖ��On`�R���m}�=ʱdcIބ����Zf�i��Ǉ�Iё
>�;8u͢�7�(/����4���"!Gj�97ߥ�ʶ ��/�����ΰdUY�;��r��Xˣ�d-B�e����]�b����ޓ�J��7��_���j�h����U��ذ�Bi����^��7o;w w�\	�څE��}�}/V�[� l��>U�������ܰ)B���	H+�c�%Lp"eM�vB�)=���r6�	j#8��T�->�;����ADӸ�4Τ�X��p|Y:F����IЊ?<���X�V����FL��U�'��� ?kfM�RT`�z!'/��l�'��lar���7�rEˍo�Qfn�Š�'��9]�*�m��X�ř��M�I��e*�6^�@^�wq�*O�EJ���\�F��{��~�����!��M"�����'OP���"3O�-yQ���tx���w�U1�$*�3�;QY�QOAq�>��bDWc��r��2N�9W~�վ6�Q�Ϥ1,��M�2Ѝa�!�+�iH҇.vf�/�d����k'�Cmz�V�JX��=���8ޤ���ā��d��+Rh<�ճew�+,�x������L�]���N ���<���rl��X�4�Q��L�}������C���1�k��>$]|��]����q�e[��Ο�t����2+F��.֍�4J��[�����)~�>#N�ꎣ�t��56�r�
���*(�D�)<��1Zv��?��H��ǩ0R���ť,�4�<���FY�<R��z8ȕ��	��I�v��5�<���V����ck �S�a�ӂzHNn�����Z"��� Gӷ��5����Еh���4%I�݋:�e�qG9�M�mT�S�h`>^d�=7w��dD3��h;�0��˲rw2F���w�� p�Q�Z�Ecq!j�}l�lk4Ö�m��,�����-������4G'�:_�gmxH�4�b�5	�Z��:��&���'ͼ�vV~�&��)9�d�zA ���9m�x��ņ>z'�pO�$ڞ��Ǎ"��L�<��|6�����Q�蓩�"��	v�� ���
rY�o�w궡޷��I*k�Eݽx:�u���,��]Ë%�����.pN��c�Mw���uח�h��;Cs��wF �����*�~�R�K�c��V��7'k��:e8�,���4.���܅n�t��y��>����w&��zhߵ;WB@��<�e����N�����eK���bUkt��1Y�mx�#�_�o����f�h��I�+ÁH5��D1�����=?�S��{*>9,R�����P���;��:HKC> �r�}�fMg��v�\js��fU�S�2����&���`�����5�+az�V�H�k�"��zɸ�\d�3��?'��V��龖�����Ƭ����K�����J�뷴/��b{��U���ƞ�b>���0��͑_u�����X��0����WAwp���m@�pQ�M��!J��!�1\�o�!�$�۽��kE�+�*�y���M��s��ى���d�b������e���18��@���.�{=�|�䭀G�(�������#��*���ݜ5��P�m�vf�4qG��~��[$�,J�5k��;��F�a��J��ϻ�G�]ޏ�n	��cWQ��_�<�r(!`�x8�͡Y��5��?�Hc�0_3!�������ݒ=������e�?Z�2.�3���3H�9�f�9�
PUd0�=`*�L[����Y���{��݊�(��WU���8!Cc
c��IgB�G���%!��0���..}�BM��JZ12�f�S ��b����'�����j�RU���o4�������^sUړ�5oؼc�m�iYd�®�!~ι�l�vCq�,&&�����	rzM��$d���yZ��ڠ�5���>���D�d17�w^�cx�/�^і���,�~���ϳ��n�ʈ%6��	�7~nBWݞ�����H���vt�&N$�Ϝ�XVz��	����1��x��,556��&;�bHU��S�|�E�f�U T�+Ӈ���9LHI��߼n����X@������A�gnlU�Z��,n�|r���q��
��ȿW�%'�n:>��>�QȶLa���u��r�i��pt�y��r
�^���m��<bd&%y���V��C�rw�P_��+x��Gc%�����;}|U��I�^	s�H/�R�@>h�t>���D��z��̺�Z��q	lv��9��S�a@�cx�0/��<e�^u{�]k� ��,ͦ��o��a���X1�QY�0���6Gq�s��LM���B%��d5s$�����=�A�kLp7�N$���泝���C���f�&p�	1�=)$���t��B��>��9�ɖ&N?���7#��\[��:Um�;��s�����9Ƭ�W}�Qjӑ*
�(�iW�7���2�E���S�������+.�~9|m�����R�U�Eo�
S���܂�4˰��6ES�_�ytNyd�㋒/�-o(� �&W�CJ�E�RX > F:SC ��)a�&����p�Kk�h�y0�J���5�V^��23��nM�ҋh>��ˎ�4�F���Ȟ����j�IzC�ҴE[I@02�=5�ϓ����� !;;���ȅ��E/�ԍX�-5�h��#M��5�m�������6Q͎���� �Rm8�F�x}f�t:�lx�L�̂�Tw�y&�ቺ�]�qJެ���`�<1�=��ghk 2�3l�ˈXR��=#`B��[�~3��ζ�m��Bz�c�3 �[	�����H�!g���u���(�PX0��kC��	��������?\)�x!0�e$8tT
�@��'��"�qZ�gm��Z�GQ���K�q&'T��!��f�� �G u�1���,�}����o�fM[jY��Jı�5��Ծ�I��"� �|��Ƚu���z�n�k�%���)	�l�E����a�����m;�;��g���0Gm��Wc�|�H����hUQ��ɨ��6�X��w=��}���
�� l1r��-�=�)�sꑋ���Oᕒ}�Tu,ڷ�k
n�?9{N�c������8CQ״Kz�e2�~э��J�a�#>]\3h�Q���P�t��잝����|���f��H��Bg��A�H�pa�[����Nڶc��CL�H�`���=o/)���"� ��+E\���E�)Gյ��Q䔙�$?���4"��M��F�UY
!beݙ��1�����%�G�7�u�TkVU����d���rX��:����t�fa�z��A4�t�F��KME�1�m�:��� �u�yrx����P4�֗hr�*V%�_慚uu�U�/�gW���2d�z��Z��`��a
�f��Y����aqx��6h��R`�v��^f���4�ֱZ��^�)�I=�>R{yCu[������U1�q�i��]Ο��8�g�&Rz�?�H��D2�������~�t[�|?�
��s�N˽�J��Iq�~~iD��Z�{$ �{#�&+���	�A�k��͘T�nM� �K wũ�H6%i֥<K���f��I�*칝g�˅�hL��=|g����8�\O)?S~���4�0V��Mf����~:,:��<���b��RR���K-P=����3?�:�������8���7�p��P�ݮ"�k�����=F��Lz�ZF�ڜ)H'��-N�d��ߏ�sW�g�Dc�Ҙ�{�C&����_�||�pG��RI׌�C���9����9u9Z�_���)j92���jC�}ŗ�X@�U3�8��i؋S!�c��X4UOg�)�,�s^��^ʚ��}7���E*;�91��(�=r�� ��bT�x���j"�ܺŀU8�0§X"��)�^�4O���y�]�X	p�e/�pY�	��~N(�j9�,�G^�����������9A���VG*ζ>�:O�"l��lZ�iy�mk�1
���:h`��p`+�����*Ӑ��-r7���� ��~���3��E��)z�0��k�c��:IN���e��F���Bc�W<���K.;`I����~�Y~v���V�p�������:$�<Q!!�q#2:�p�n*F�s�=<n/: �=���Ii�`��/���G@ҁn�Y-�����V�����6�5�E3b�q[�9��k\������㗊l-���[�\a�e�G�g��^,�t�fD�2�qy>_��� ��j�i�az�f�$(���K��pH��(�R9B�m�h}��k����	�0n�U���Z��Z4	[�W��[M0�l�ډ�+T��zI�a����l�����:�ظuB�t8����5����Ǻ�@��d��r�a�Sk3����������p�����S�Y[����"��U0uw�oJ�w�/�6�Қ�b%�5��	�`j��2jCz 	Ai�^��1��
3�M��\'4ƕ�mF_My-�ѿ�7<9��ȝ�M��4 qm$�/0W-��\�|ؙ*�R=��l�keXS��:�w=jG��{6"]�P�����*�>���&J��-���-����J(����8v晦١�o�0�ԝ��K�ZM'YaQs/��Y9?
bD�B[���fn��I;�1�-�>�͹�)�K�P���6��	7�G���]t��0��݉Q���J؞)a�-B�A����@�u�<�� &n2�Lncf�`��&�v�P�|��6m�p����%2Ё��V�ǿ��Z�@뼍s�j��PH�7PFiOp6uC8n��$��v�������.&�{3�%Mm��/�)�t��������C��wa�p���t�f��/���tԽt� ��+���;7�>t��E���96$�;$�����3����0��LjF;��µ�E����ѩ�/vrߛ�(x�1;�@G=�w��S�K���wQ-��KB4��>��Ĵ�*5��ڮ���y�4si��L>`�j%]�:�G�R�NDW�^�uH�>Ϙ�����;5��-��#��,�B&���N5��^�|ߩEd�CQ7�5�����>ꠏ�5}���zS���hYp�d�_�°����&ȍ�i��t��.�Q2&I�h�<�����ߝn΍�wK���7O�������gyg��cΐb�)N��w{p��� �^^��$4����T��M��:���e@Ϣ����@b�fb#���Z�������9B�3^����)��y�q��=Њ�ǿ��8�"a�MG=;3M�tO;Eu����Kި/־�z���d�G�$��ޅ�WC�l,葀B��q�yN��_��(V�~3�6�(xӶ�R�h�Y�"3�C�?�L�ѫ��;$+�ns��$�Ml��ΐ����2��q�/*�B���v{um�)ƭ��[�������H�5��I�=�?�Y�����Qwp�����kD�~\R�f}i{�x7[E:��4X4ҤT���	��.s�ceBm�&~G4�گo�y��G��}��ā�C�Lg]�=��Q�3wʜ���!̵����w�ݓ���^ȴ��)�.YI�6(��03���|�A�C0�|=6�l�I�_���Z���`c�"V��U�+�AMfq�g���0����ߝ����$M���P��2b_C`4$��{�2��Ϲ6��!��.��cBA��./\h�'��Ɣ�Y�\�;?5<9z:��pA�i��#�,������m����-��G*7�'���Hď£x�7��j��FŨ��61��h�"o���rQLh�S��gHwO��8O� :�`p�����l�Y���rV��ݯ�Ih�������0��	�چ��3ǧk�L�[1��o%=b]D���B�o�FE.;X����s$|��XHs�P�n4��E�{�Eyq��4�Ng�Fz's�_��eo�'OdFS�X�i,����( �-�ukWҝ%<*>��-�Z#��ۂ*Fx�M�UIw�G���,��b�/n�� ���?j�(J�k5!���0��kN�����V�nR��!&k�ؐPE)� o���?Vڟ*rQ�1��<׌���.�
�;=�H´��_�P�(c�Cp�a��9�#�4�����P7���+w ���sN\����#C����O�)��e��o�a�vV�
g̶WB�F-8���,�.��R�?Ƽ�z��Q�>��k��zc�,@ܨvj�=D8��Kx���F�KXF�Л�C�pf�nL��̤��Cn��"�����|��C\+L)�GU��:��H�*jדd#/�u������8޷���9����X��(p8vՏּ��Mx�9HQ��y�õ	�����M}���?a����ar�9s�q��dp�gm�ef�!�� X���$����Q��!+m�J��L��9�N�O��SVa���:��S��\�2Aク-��n[x�7[��cG�}�L9L��$ �������b:�^�(+!��� T�V���ߪ�3/m��NQ��'�0%�9l2>��BBN���]��X�c�^?�"��j�L�]0 ��^7�v���=�>m\B��'Ѧ�g΁��'��o�W�+5I�ŋ���Rp-N�Țz�dY�&��b�[�Ca��������(�&|Uul�s��D��0�n�y.���$�snJ��ݹ�֑V�}z��dX��.�01� ���ѧHo�����ahI������5�Bï�R�u\ 'Nl%H�F�-��������Hf p_��l�12z��`���+��_�*�����<%�<҉�,�݃�xZ�Nn-@��3�������{�S��тm�������$J�|�G ���^t��yp��Ր�'�3�6 �q6�����A�D�)/��{2P��\֛\:��@CX��x�v��V�n�@,&,[,qX[�X�˔�ae&���)�ث�~c�"�P�����F�p�7�D	�f9+m#�����9�{���*S]P+��-�7�?N����Y�e���dm�6-Qy��0�l����vW�m��7��Z������
L�|(��"f�C�l��H؃�{ �����z$���Ąo���X�=?�F+r����������l`�>2K$H�c��N��=}luX�k���
H#-W۱��U_r2��p_�_���z-c1%5
P
�[)�UG��1,Ե��� ��F.���r�4CF��k0)��;�����ݪC��I^�'k7�e�y��5���Q+)x</�!ҡX��4ec����(�x�px��R+�q�-{�n��C�9-݅u+e����S=T	��'$C`�|�m]����-4>�< �Fv�"�c���->α��Q��a��p�wc�)���ӯ��l�c,,2��An�F��Q�>&�l\H�Q�r�=�.���T���Σ��;j���W�G>
�Ɋ昒wȲWn �_�n��;hݼy���j"��g�':ɡ/}�5�s��cq���#�d�+e�ZYo���� t���4@K�-�jb���:L�.�lY�E��V["C���ԩ���5~�BCMOY�M�~93�n^����'=\����=�il�)���k����p���}v��,N�|i�����V2�=�@ħ5�2Z�a�"Z����^�G���<M��u�
�G����)p�ujC!��X��a��W���">-fv�$�eY�S����3�~�������J9\�����2����sb�q�X� ߨ���>1�� {���`��Z�z9M�~�������6�V��Y��bwo��6R�䰂��4r��D�P��&E���>TP��o�q<�"���h�:�Z����1������u�&�� � ���۰���a�|2&��+r��ǒ�{�d���r��_R�6$��狀�Z�:��3ω)��2��%u8c�Po��(T�w+_IX��Y}��D}���qC��%����l���'�M�j!`
��q/��E�����w���!�0N���g��ѨQ8́�)<�k ,��i!����;�N���]|�w6ߢ�ҜO��`�^��ӻ�S�}�Z;�i�������������6�K�G���U�J��3K�A� W�݀\%_?��|��Z�,��kB���PGR����L�r��?��NNzV����qH�^�3��E�.+���� ����0_�}���a.���7���y@n-G�0����5}ؤ���kGi!4����]\.��}��F�V�K��1�Z,@��y��1����} �L���ΚiɮNo4W
"��:{���;T�����8�V�{<-��0���sI�&�"9�t6���bC!<U���%��^d�]Av�X��#�o����ٽ\�9 @�,��Ē�?%,�G�(Ƞ�ƈ+����GN��IAHG�{
'���+�Q� �NZS�>�ŉ��{�?U�l9��L���w��D$��K�!�I4HK��8I�
��Ev�!��t��A�E�� �O|_f�II��J��$���R���t�h�,�p�����:��B���k��"�Y\],��p������qk�P_����-cS#��e�D{��u�&�bCQ��d����E��!MX\~��v�'1?��ҷ���у����y��4XP	�����q��xdث�!Q��Ϛ�0���=�OP_0�I4�U�hOf��n�i�)I^�3X$Vȑ��;̖Y��r�#gzO�2�
�9�"O�ЌT�aN=�>�x�ӢL,���Z��s������Y��d���ԁ;b�N���O��<�),�@60���rw+x�2˝���ˋ����i���H,����̰�<�ͯ��A>Q��l���W�a�W�dB�hq�hh /�0樊��tַ��6�����K���VLb���8C�,���=���\X,�}��+��J�6B	���kn]��3��7��u�mذ�U��E��������hλ�����z��y	���T|�Փ�PQOt��u3x_���qp�&a��n�D;놴D7'dQ�{02c3��[-����f�����x�g蝈��`�+�M�ż�3��j�ML�<F�-./�a+�联;!�Z��{�c"aЭ*�~q�N��>&uB%\�d�4T��{���N�o�����Ӫb G���a�y�*"�PG�|��iU�-"U;L�8y*����E3yP�������@Wj��Q��a`����:�Y��W��gc�������%��؀����a�"i��=�Y]�9Ѯ��5�7dzGV���G蚦R�{��.K�~
qlݶ=�����z���Ҵ���lR�|���=����Nɵ"�������l9zZÌ���$��t7ƿ��_3H��	��������w�kX�����,9Hߪbյ�=s��z6�,���~*^�/�6w�ޞ䀝wɉ���awW��e�V�� �f�1ƆQY��Θ���6+�r����Y� ��Vμ5xK��D��]U����>q4��[��� ��<�qwXP�A�P'}^-\��un.2v�9��M��<�Z�
 �yp�NBM�j{�%���q|:�f��6P�<J��X�3ւ�ˉ��$K�a���M��\�kDG���QF8�y�)\.�F��c���b�&��^��Ao�cwR�_����mX4Ƚ���@o�:&)?����ҲW�ogwvG��/䲭��!���=���vJm�҄���V�Tv�/���Yp*Os2�v�8��bj����&���g
!t�P3K��0�NY�ǕQ�B�ƃ� ��^o����kB+�"����ْ��VCV��Qh��Bًp�]�� ����Pk�ֽ��������ɽuֲ������	��������V�2�f�ボ��T5��L�cH����H��m����a�[6h�~D_�9zݞEc�;��9)+�