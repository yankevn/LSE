��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�	5w��O�̽�]�ɽ!d�`���٠�L�3��>�TI��Ft��"�e�3j���!|�x�����S��D�|�<���2�5���cBQ73���ƭ!=�҂M��|$�5u�Ly-������a��^���r$���M3d�n�Є�g9�SIm(�|#�7e����6����a��\��P&�9?��Z�y?��l��M��;�X��ܽ�7�Y��9ڤ����v��R��{z���e2!d�p����w�����?���h�9ؖ�3vV��:!!��˯��q�-������$5���q�:������r1�/����"DM<��~,@]�"�<Y˶�����l�ɒ���\z�ғ�b����H;	W1/�o� !c9X�� �!��S-\���kI��i�Z9 e����; 96�0�OQ�sĒ�E��O�*�W��p�ղHcӇxϯ�^;��I#8N!�Kq(�۔οnS�o_2�u��i�����cʍ7��ݔ��#�������.��l���/�%/��ez[�\1�2�2�'%denìp]���
'�k�������r�r�~گd�O�Kͣ^ �9]d2�Ct�?_[��W�Ȼ�QD
xڽb]X��~R�p��(����*4��G�4O~lL(�>	~�]�`��E5�&����o�s�%O�����`�!�H%L��>��Q^r���w��m��*�K���ƺ�ر�d�`��}�������^X-���C0�����XC��R�髐�RcKԂG����}�D���?�{ߴ�q��~�vr�>�K�y�B��,[�dE�G��p~4P�v�d� N�=\!��mC CU�#2�TC���8����� �ׁ��p��G�6���Z����q~UMn��I�-�|��B.����7'1�(�q�5�1�3����a�T��� h%�{��J�AwLR�j0􇊇Y%**���u���Ma[kR�{�������kY�����6�]=���WA�m��S��&�\v�qx�JY�I��8Q?"��Ɯɺ���yp�&X�/��r!��Q�q�ڷm	�#I&44%ʿ�qZ��H��c�x��x��qM�g"�dƙ����X180$�#�i��k��𴀣�:���V���F����4���㎶x�H���~�+P٘y7G�q���YL]$�eX����V����:I���p`*X��<8��Of8�rq��Eaf�}�0����{��s1,A��Bu)���Z�l��lI48v
:��jDnuoJì�������kh�1o��A�b;7��ڴ��J�I�_�Z+ ���k5��?,C�u������8P�g�Ч��ۦ�<��"3��˻�_9F3�0Z�+�H�g�BDW����Ƿ/IB�`W
���-d~��W'�o�!���bP�;w�נ��tj�<d�4g[^�����$"N�]N M�g?W�?��h.��'�M�Ȧ��m�!�5�i-���FplUs����
e'�9w��Sin=>^Y?��,,7OB{���s#,n�rBÓ�=���;_#h��
�?��WK���!ûm�I�D �k����"ö8�V��ܲ�,4�:����U�ղ�~����ﯨ��a�l{q煅쓱L�H��1��w��ꝑ(��?^��	���zӽ��_Kw��L��S�6��kAͳ���:V�4�=70���F��5�=���b�tqPQ������� GtaƊ��9%�	��K6N�����k�C��̰Q^؏S!>𤹎�a��}n7m��|���{��w W��̑M���Y��~�\��B*�o��,����"�Gj�PH "��� !�����0OPb*�^t�l7������Ќ��!�����|i�QP<����M�-��:(�Tn�XU���h�S@�>�[�o�z�i�jJ3(6�=�����FL;��m�O䑴S4���C���f_PB��C3��Dq{=Otp0#� i?_��`w�ZNc@��[�a������t�x�z�Cү����R��x␋����>��AE��ޜW�������Ko������M�"7�/Zt$�Q��*�8vڦ�����*|�L?�o	zW��*��/�'��IL���XJz,S,���y����sMi�u�_�V�
j�\ډ�hώ8�{��q�c��0���QՈZE�&��Z�?ʡ؀���]�$y!�O>��i��VC�����L����u�@�&���c��;�J�Y�d�QbC���N�t'����R��bM0��D��1�1��҉`<�';2�z������d�?���a��l�f-�e��ڤD�ݔ� ��Kzr����޺�(��^O_^N|�.��~]j�9j�G������d�Υ���j3$�)�������/��p�\:�}�XL���"J�vE߻͉�9� [����Eڍ_�F*��&*�v\1�Z}Aq�s�BS$�@��_"}ҧ�!�g'��溜�����V(D����
T��S`�����.��e�	��O�=tE�/��!۵&�IS�V��&�����0>RrxO��� �Tc�m����?|���K}s�ɸ��;��@��i���ǘ�����u{@ya�����׊����|u��`cx2�>�K��g�=��o�k��!�c�kwzd�:2��+Я�U���"?��}#h?��h���2�E�'����:E���o<�HaH40?����A%�9��q�J�eP֠hy	���l��f;�0�H���ET�hXp�H�`���S����.��(X�;�2��'�����rQ@T�<Po~YI�6���Y��,��a&Ρ�>�'&���%VΗI��(�[������6XL5�����g�����S���<���+!������Y-Н0��*	3�p)�,�.t�3�0���CX�j1(F������]B_�/s>�l���fꏄͱ���%�$%�Q�@Hy+�� ҥ=�M�0V7j��H��\��:�����A����o���.u�<�sФ�� � �koZ��Gy:�g;$�bw/�c�K��cO��~���`���Q^�J��#F�h$��}��L��R��ͤ�h8N��I�\d��b:.��F��N��:��L��Qu���B��*tk�]��U��nB��q������~'�'P��Q��]��!�q�~��)���'y��q��D@m�U �k���ե���!
m��I�1G=G�o����s��p�&I�O6w�)�/��؃�޶�o������ۑ�AΒ�(���P� �w�)8�C�]P)S�v�(�LVCL�B�.�?