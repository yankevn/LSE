��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��E'VTEB��A)���7W�9_�ľA�}�����+A�iȘ+6�[���u��y�����9g���hə��:��e��oKBm�Q|��P��2�5\�xf��($�z�Y��L8&*
������ЦU��C���n���.|��Z\�5i_$�������D���T�g� �UZXr2��LW,E4���i�f��o9���jr׼��o��sd��{���+~A j��c�|�l8�e�V<��^�?�"v�2�[���5��L��3Q�p�\������G�6x�J�έQ��y1�O�NG33t�M�� �A��C�م/aH���W����NSS(`���֙��)o���z_'�c��k�Y�+i�K�j7���&l,� ��<>j���H��F#�
* �J�����Ȱ��5a�绡(#U�S��Y��4���j��C�=ov�MP�)���7%MAh~c���*K{�Rfv�^W)�  ��ъn!�ߙk�F�уm�� ��m�J\WL��{�g�s6�qĳ]���^W�0jcx�(1�8םc̊�!\��pɄ�V	������Q	�*�?�8����ߎHb��#L�`q��h���b®*%��꧶*��I� wR�S�-����z�r��:*���>��T` ����',f����;z���C�+����߻�#/Mæ}J�U�C�/Hw9,�Y�:8ZÊ鏸$����cm-�%��$���"�Od����e`D��G���0J�����}�!��E�*������j� �*�T���z2��<�ܼ�a�X��jK�E��F����ۗ���H[���a��ӥ( Yk��]i�T£�c�}�K	\dʹY��ޠ*�c2���i}��� Ɠ����}1�(�{Eu2����`��,�ew��-+{]Bv/.v̏ώ`A�v=K[Y@)�ϭ���:1��i�ϖ�� Ȋ\�_��H�;��$����|q�-���-����H��6�������IU=�w�(z�C�OG��M��e�[�g�]���-ָWh��2�t���}2����k�o�x�j���b"��fٵ����j�t�0$N%:�'�з��6�\ɳ�'�.�	x#uM8s+�F:��?�)�W��j�=Q�4	�r���y~s��>���Z��a��[$�8�KƐ��0��5��(`^W�_���˂@�q���b�3��n'�ۇw�0��Ce�U��8��=u�Z����
W��G$���O����"l]��� ��49�.����q�9DQ����爮�d�
Avc0"��.��q���P�V�O��2R�}�ے�M ��������hR�۸�s�׻rX�|���[�]^\^<���>JP.�KF�41�F �X�g{��㵌?�ʕ�j~U�m[a^%�{E�/���N�.݄�N�(�+��⷟�p>*}����b�0؁4��!J�ˣAQ1�(��>��,��@�apq���i����(�)�Mq�����W~ԇϤ6���7Fc��zC�*��m>���S a��a����	5�'0������j�b5�"T\��f����n��V����&}�
�@G疄>>�p*�=Q:|g�N�%����!���ew"�Lݱ�#<���m���gW����2� �\߷� �4�l��:I�h�.�Q��t��1�.������f��ׇ97��f@$�vQ�+y�*(���.ۜO����UΕZh�=�OH��:ǰQ��}��x1c*��h�_��[�G*�a�� �o~�g/<��[x�F���6o[@�L)]��̱$�4T�蜨�E��W��1TO,�R`��
+���)����oQ6DJ3`B� �0Qg�U��+����4�X���F/ӎ�}b0T�` �zu����%��>&��]y"�$z��;���Dã0[yE��͐�;�м�C���BhrF�Ms~_|�Q�^��4�pz��t閁�T���Z�j�n�t��~AA^�s��u^��~�K*��`{ڜ�i:�L���D`�2��V���K��T|uLyࡍ��Ξ�E)��54�N��}t��Jj�O�{B/�w��Ë<�k:��E�)�줎t�=��;e�*�SX�x�?��wn�f�P���%k�.֟�Nw�{ˌ��{W1:$���;U�3�`!f��8�IZ���I�5$rO�4^p5�������6�ۖ�;aU��"����Rn7ȧ��~���U�,p���:���I�Hpט�T����Ȝ���=��r��������1��ߺ�c�O�(F�hW�4#24c
������cQ�J2q}�$dj���Z�*��s|a��t �T)$L��}�(���I�
�y0��/�b"oQ��˚k�P:�m4t�'I�rGA
LG癥���nELX�G�Ez���,5(_�" >!�߰:zv�h~=ۍ������g���WX[	��Z����i�e��c��O��'n�(�N�/Ő倎�?G�(x_U��P���4�\�Ө�M�c����o�E�E�&RXt|y��&�<�-�
cQ��V�r˽Hs�U
3��i'ŻO�����"_}�w��!�#���ǃƠx�	�?	~��zر�����u���m%5kN<H���\'9bS�Q?������P_��{�ٟ��5��"������a98�j�4�6�!te�6=a���6�ƁWN$U���x�����
7"*\��4b:�S��\�76~��7�8�O_��{�Z`���0U���8l�}�PJ��^�-A� ���-�������/pa���k}�&�ͭ$kXH���Sה&�4�.|��,`G�o�/T�̥6�J�Ӥ�t��Sp���U�\�b{���kEi�,�AyTҧ��2�ҟÛ��$	>��J$��K�Z0�B\���Eq��	�0n����~�]`$��6�CM����3+��BĬ3�$Iȩp��Ɍ�L	�����x̳��X�˱�;�%x2Hz|_����u�ah�/j�FDY�B�6�ٳ�?�0�u-�/DXV8��NQ%>�uv.���X5C�ؤ�0��I��E6��p���F׀Rs����ԧ�!>�x����svS�1�_'+X������<a'�y�k����w����]_��Wɹ?����3]~��dkx���ۈ�@�W�5N�V/θp;+	'�	���8a�q	p��R,Kq#c����3>
��7�x��*��9�dC�=k� k;��[E��Q��s�^�{ ����q�a)2�G�(b"��wR���@�~Զ�����R�Á�_���Ԫ��9_)�y�3{�dS����ei���;���$��~���DZ3tx�0���c�Q�¹#�;���	�Sv�ο��I׋9^=��0�9�L��	�9��B�}�x%�|�=����jV%Z.���oZ���!9���&75���ɍW�OXu���G��rB��ط�w��΀z2��[��l�o(����p�W���{ݗ&)��d .��MS�)��w�8-V���gq��sh�/$*X<`�7��yqa�m��3�s�����(���?�[��)�p��6���!^�$Bvq�ĸ�\W�f`U�x���k��ȝ��i}�/�L�C��?��%Vb�Tg�m~:�Ӵ�Ne%glM����h: Xh�hH�%���Y����a�=h��ѽQQàD��b�����/_�,��C��)�Y2/����B*DŎ� ��d�e�}N/�3|v�z�FYI)O��c���p4�5�?;l%�U�
ve�"��������/���(|�0E)����m����R;xԆ�R�q?�uI����"nr��
�R�%���D �a�Q��Q���K���6.	�5\{�UA�*�5N����P�?*p{�}���l���:w"�
�#�Ԥ���*j�v^Ҡ�Y$�\$���b�X=�q�ȯ���e����m��y&I���ve�Z7�
��Y��ծƀ��Gq��,0��'pwᄊ-�8J�낭�z�F��ѽL���1_��rƛ����~�4�zN"��� D�&n���@!>!�o�����]V�ݡ��ή����3�j�n� ���ӂ��<��ԑ��k�0.?0��1���U/��uVSE[�2c9�'>G�	�.7ƽ����+*�Gl7״}�h��C�Ju=�I�?j�G{G�Pɢ�/�sK��������3��)e����kS�u
�	���´��0BBB�fs�dP�L�*�B��v�������X�Yh:#�v����?I�
�2��/�����y%�K�B�"����j�ا�\�*� ���� �sq:Z�rwT��.���y{���
Ш	�~����� \���S VN��/"
+����S;};_b1�YQ���/��2�2b(�mBm	C7��L�Z?x]&�
���l~��h� =t;.�ce�H��<̲V��D6���h@�r���{f��@��W��N�i�Q��[���2�LSa����� �7��N��bJ���Z���Om뢁�hڐf����ĩq�$�(��,��	��`ٴ{��}o��\���f�*n��*��RlP�>fGq&���}���qw���na#�w�a��=~��xUSw�V��e5��f4ڡ'>����0�/��>@M���L.힣v�$[�YL7Q2���@PP���TF��nѰ�~��<��ꖂ��3Nuy���x��F��Y�˪�kO�Ab�I�)�(�MGeۈ�k�18�D�����=d��zq�x�.�3dK �r�}��؎2o&z�@>��1c��N�%j�ՁoI`���i�� m���I��Q�m�m�Caܴt����N�w�o��j��m�랐.x�SC̷�.Mh��n�巯��ۖ�,�1�{N�$I��j��4�+Vf��/B�m�#��PC6���N�M�t�z �N���fXa�6n�t7�C]�����A���O_ߌ�w�U#�ʗܲR�b$�9�;�^�����H���]K]��H�۝��!��=Jqԍe4�U�t�hd��T7D�d,j���h\Ho�|��	�7	2Y��_=�$��qFi�����k��� ��*%���TnTLx��h���\��A�XJ`Gė@2^l�8���~��.Rs���$��q�,]֧�� P4c�U����d�J�Ֆ�h�f�3h�A�z9v�$��J�?��0y�T����1!�nx�C�f+���b+LQc��� ܤ+6�<~	9v��� ?�FJ��>"8>%�,����}�q�('�K�w��Yĩ{���o.(3H|:cQ�S�`���M�m��܊�W����<��I,�E�n�	�a���Q�Q��Os�U�S[*AM�D���d���B�L��'`��x��L:�=D�E�IL`�\.��Ų�� g���c�ܡ/�X;��/�%jsH�}������+���n�W�Ԇ"6蔡XȌО�����g����C�*[��rc����&.Fd����Z^b�d�*k���L����.����M$)��(�E(�*�Qs��O�Dt7��o#�ƀQ�R�H��w����ź'�yJ'{z��H|<��Q����Ve��]&@�)�D"2�>��(x����4�@��΢��e�h�~��~��_�PZ'9�h!�t�*h��Zy��x�N�?mc#0p7�4b�2��>�$d-�J8[T��[�
��K��pV�$��d��`��dd��jfQ��X��ܩ�|����|��1ς��s�|aY�ʔL�Vk��pL^?�Eo#�0���*��4�g�MBh�v4�T��P��=Sp�RP�='?�K���I�����!�����J6�4��_�z=j����;�UO�KvA��o��+��/L�'����{�-�L�u|��7�'W.1>�3@���}�}#���S)4��0#]M�\Y�9C�$�֕3P�8���ӞHm��G��ޱ�I$z�E���Cq��FV�b��n�k�%��ʗ�gO^Lm'��{ˏtᘠӃc�B�,,�vN2��=�F_��e��8���\H@��8a&���M4m�it�c�� fU$%U�V<���ds�ҩ�����Yl�=�ǘ:E�N�w��\M�Z%e0d�[Kŧ�B�!���7��%��p�êBMD�Y����Nڸ��^n�J�k��
ٓ�3hբ���|�_p�TL�u�ѨH�jo����H��ej0�%y����?���@qK�#XG�X�e���A����^�4N(I��+�n���� _5�
��7H"�f���l�.}�@w��#�l���p�Kk�a+]���[d_Gmm7U[�mZ���V\��e1�B������L:��ĢW�M�$e[��M+�ݾQ8ŋJ�q�6y2Z�QRA�
uby�q�mK��a?���J��ڬ&ׯ��ͣ��VH�_�Vta3�=�4n�|�S(�@:�%�j������M�"*̩��s��<t�#U��m�*�C�Y�������F.-O�����e��'ϒ�&J.`��C��}/�HY�A��Ou\d��f�n��;I�5��:[7���G��U�7� ��G�b��[V����R�<֫v�p�t�L�Y��@�YE$�Rh�'P��NSaGj�?�������^�nH9K��D�;�>�G���d���rJ����e��нĚ��.3^�]����=�Ȉ.j����ET?y�'�9<q̤S�����6�>>
�`4��8P4F���&��6���T(,&��U�Қ�� <��TUbi2�K��C���/�f{z�d��S� O���0J�W�������R��_��#��\��?��@�#�J�rd���[eH��`5��&�\R���ҷ�)��]
���m4J��ֶ嵩#q6Xہ��(���tK���PJ���7"���p�7�1YW���pi'���ˆ��Q�R�g���:5�G�^F�&��D��6m�ʬ��w7'lX�s��"�6�%�I4�����[�V���l_�h�Bc`d��(EM���5�rpw.r�m�H�h��kD��vl��d��7���?}{T����
��耛ۗ���zlSL��@�@ɬ�B�a�sf��<��NI���x:���<��=��t�O��p��)�v�Z^�M����&�{*�� �K�ۭ�+�
�����|�<�Ix����/#\�3�?�����c�oπU(�z�q�w��\IV8�#���i"��b~B���0�ъr5��������Mcْ#�fa,M2�s���im�/��j(s���X�oEܷ�ԏ1��(�:ioD -� ^5��g������9NAÓ�	}��%<��h)*��p-v�K�� ��p~�m%r5�o��� �=��(��Y��-�h mkG���/of�Ա~��]�>y�\�D':� �
nHVxP珙�+؏y�}[vGQ9����������RV����^-�n�ɝ!��I��x_�A��[�z�gXKX��3m �a���^�8r3�$k�ث�+��:�y�֘��k��^(�̜�����+�ʚ
7U��[i#�oR=\���6��!�v��0"#�ӣm����ZRz��0a�5�ؕ�t��i�P���V��Re����ֿ�գKJ\?��ҕD
��G�5.4��s'�a���H�.`Q21}��
*�O%�����`S��\�(�ҵ�������yv�k��ŭ\� 錷����H��}����������R�Wc��}w��kM�z�7����<Հ�4U�g<�?��Lg�2J��!�Zs;��=vx�P�*^�.P��m)��0�"�2�zj������m�̓?��PkR��ttWz�	�Bg*3��.��n/4�����cPz��jT��A�����d��udU�R�i���3'��%.S��32���N����3P(uZ��@b�b�'�QbC�>B`]�����y\��������^`F'
�鱂��d0������^Ue���x�ː(����&��-~/�dd��:���U�C�9�
W�Y��J�P=��K���l_���#qc7��Mp~8|?Q9J7{Z=��q�v6�yG�j��~��9Ɣ�뫟��"���Υ�3�n2:�f�Zz��dY+�>fvu�WdP�NAѣ�d
�Iۭ�+������'~�
�a|�'�;��*�cr�V/-O�'beE��FJ�?P�`Jٓ7o"�>뽏�Vt-�.��b(Z�v�|�gX�ɾG���M�eF�M��>	h�`�-#'P09Zi6��#��/r�4!�<��Ր����(	����"����������I�@\/�������>�Dne�ǘN<y����J`�+���:�AW@}M)w�ɨ*�Y��q��2MgC�����]�~�&i��3)J��-v#�.rᬓd�,^Sjَ�׸¼�1a�*��k��K�
u�Z��g����He�=3���,�|4���dSJ�]���	���A��l -����zZ��F��{@�r5�����Y�˭l5U�j���B`
R��*�9Q�5�٨��a�G7 ʡ���W�c���U���?�o��(w�L@W	�qEkl=)�N�1T����d��gpD&4�L>��GI�(=R����4����v!Bޑ0%1\�Tc��I����,d_�z������r�P��Ĝ�}�1���9���y^��ߞ�"{7K�
簗�蓍[d�Z���li lC�d�����(��5|"�.@��9�j���OKu%?�J(�r�t*:+NO)�!R�y�2�	������e�Wۈ�.�v�5qs���l�D�d���;�8vt�K�ړ�ƗZ��:JA�)�<�WLY����p�abu<�^8������j~��iª��+H�Π�	cK_[��A �D��==���2�nÔ���._�{͊-3�2��
*�r�+�錄M�E)6�T4��J5E�|J��a8@]��E�"����Q)+�7���_};p�	����Ԧ3`�b��d7�(�S`xn�f�U�X� �r��uX/���Q��2���fSjQQD��on��1(3�m뀚�ê�ZB��\_�Z��,��~O_`��m��cB�b�����}��(S$��}5�a/�K4+�
6@ D�X0޵�0�M��^�����9aG�p�����dwqݖ��Z6b�8���~������ړ��`�(�A�m�ͳ��P�T���!�K� v�2s &W�C�g��e����i���b�@��&ϫ:	/��"ԯs�$Q;�/X��T0��U���Nqb>��*�*��،y4�9�"�s�[��ܢW,��/8��KgT��>��v�dZ0R�<�]�%⤷�O脌�>�,�p�m���_�H{���P�fp� ��nS:\���	����$��e���ڝg�5�k�ν�1	@ky�f�ݪ�\ma��_��:]�do�0�R�L��I!�9������x�6��I�풙�_V�4c	m���T�3[x������f[w�A�S+~��D�=fۛ�U�>g���n?��?���W�7�v�m���?�eB���<�--l� +z�^��p7w���9��R�@���k�1��9�U�s�|u�}��&mr���Z1PE���k��?��`,�Y�B�7���K�
}i���,�^�[.NϹ���qI����܇�����G��+~M���7��w��
�A��dJ�U��㟟A��}t��xt|>}�16��'Ϻ��#�r��k�+?l�"dY��V������1�b�����b���s=���E��?�
����$�����X�)&�n ��r"��wS�gn��xQy$�/��<�mg�������aaȫ�H��%�2a1MΜO�jX��T���w��[<S�W/�WWTn�h	A˕�G��]`��b1�7�t���Y1�����ӻ�1{ߔt�mܻ�M�#S��ƺ������݇ua):7xDx&���J��!~cC{f3��!�+�\7?������=*c��B��ŏn�t6!i�A�F���/��w4�\'ݘ!����;��)��~�	�)��Rk��J'�W�#��S
��k0�m���հle���|���c��W&72s���x����sᝧtq�7��S\B=9���H�[4n�c��wO�km8c�K�2�ӈ�y(Y�l����b-�i�����ꇌ�
f�<��o�9�lF�]̤_��9�:��3m�F��I���B�J�-��
a��lĄ�I\p��<�l#U]
��j��r˫�u�
�s<�Ӣ^��N�i��P��Ƹ����"�ꏒ=� !p��o�Ը3�e������g�r�g����K���	��IE�,<��TpN2�в����N�
�E��a��b�n���Ĉ�]�kqj�}o���H��>Hf	j`�SP���}�U����J@b���'_�
�g-rcm�qw�*�"Qf��!��H�Z�T0��"�y|��Ba}�щ�-U��F�4(Ē��0-4\xN='(·,�Ɣ, u+5b+f3d�����\�/�|'L	�I��H Gk����J���}�zzǉ��'��%�cv̘��y�JnT(����LY�d�E�������'��`�_��q*�"9�[T�S0Ï8�pQ�;��|����k|�d��,ц#���\d��H4��C��jG��:wcu���	��<�eXZ5�
+S �vHCr������M &*�~g ��ԕ-B�e2�Y< �\�b�oz�|��&2Q�R�	3ZA��+L�Y��^���b��E�!�z�d�XQ[�-��)˰���{��|�^��Z.��a�sÝd�����B
pO<���L��D��ouUx�}�L���t����T�ӡ�?t�T��6,�e��w�D����e�X߱^=,��n��QB'�:�M���4_,�ᢴ�=S�{7��qw3�� ��A$�}�Y9
8_�DU7�`ʇ���uƃֿ�-���ю��\��)@Y�}xzѢ\Gv��X���O��j�䓁���TMr��p�!T��e@�}���^��xYH����2���p���ו�?�e��������C:��+�k�<MȔ	�����q��!s�L�a���u��{��	�8Ay�j����WPӭt͎L-s�bi��Ĕn��?�eK��~;�D&��%CS�\`����F;n0P�"zo�]�@���!��|�k��H̒X^"
�DV��9w�ݍ�8��`��v�s�1�"~�΀��g�h�� �gQg��LF��w�s�8JX�g���Š��5ÍU�^m��3�pZ�� �`��R�`\�5�������J�F�_exkAqݲ��H8�h}�B���5K��5�d~��/����n�w�kJ�>��ѰN]S��*�~PTm"���W��j ���^}L��g��e�����Zr\e����<�KEi�ݕ��/��T�ʔ,I���8�K�>��̭��3G@;�k�m�g	*�o"V����n���2P2�S����3�PPd�M��p��V��=��*�S�t4��k����.f��ό�v����9����U�3�Cp���)�;�Wk��wӞ�I+��$"?�1���(��nx�����0��+T�c��D=^G�S`�3�j��һGЬ�du_���2 �8fh0�2��#	$�6ڃ(O^����E�]��}I�¢r�G.�����xŗ����K��G�ޡm3��rQ��X�����r�K�F�,#�:h0V_���)0~YE�օOU<A��Rq0͏���ɕe�u1�r���Y�n�Q�<��ֺ�3{"�ƻٛ��w�)B��h]jD2�!��XG ��A���G4A��/��$�!@�JKnc˂����t�,��
+��b=�^�D���a��y��8�
�@��N�kϗ��q��������D�ЯA�Ul�ݧ�]H
z-d�1�(�S��ղ1���= �����/��
Ǚbn(�F�RZ��ǗW��g�����}���1!��=� i��2_*!�������ާM/��x�/ !������E�0�gэ��5��~bڒ�|��v�q�eD@͢�� ���S���6�p���7.�[4��j.u��ȣBqt{��f�P���%5jKph��}� ���t��n5�4��ulϹ  �����<˺q��Y�w$�P��t�JW����'总� ��(������(JƩ$kBn��,$��(Fݧ�/�-·���L�*�.=�e�� ��s��[��ZI1#�<�Y<Ď�"��̖�����pE��DBJ���Eի�N�D�z�2䐲�x��°)��Y}`��\:Oǀ��\\*��kC�韽��?�����!�TQ��;P?���<��;Ǉ�u!��`8����`b�5���?D�Zj_7y!O���Ca��g��N��C�Ŷ�ܭ�M�-UxQ��%,���%�o(��;�y���)1���\�����楈����P�Ʌ �we�f��<�l����UF`L�s�A�z� �%z��:��l�$D�^��>l�'��v�ہg4ݽ�u���/��=/:�|��{>vX��!��,��<T5\�p�)�E��w�v���,T��M�Y�z�m��uPڶIv�SҨ��ѩr�����{�D6�/t��]�6�lM�XW� �Z���� ~�LH�nO�r���z�xʪe�t,P�%��O��r�� �����:����i:��[���<{�L8�J���6S���6�x��3ґ�v�EG[�e����?��m2���⮨��cSۺ��TKH-���
,�}��|�$u~UG�&��� ����$!���EB�� ��;��w'؇���{K�ϿRg�U'-����Φ�>�l������L�ʵ�d4��yf�������ݫ�P����K;}�/��| b<,;�,�̸*��*�IZ�B�LC���л�,M��H�n�G~,	�`��p�u�)o���[M������V���EܴD΅�3�9�%9����M�,ܧљ��T�}6oHh�P���E�����f���o.o]��'�pi~���e%鏓�#4��^1�#R>�󋏂��C��7�C�ɻ�E���K%��}cEy��7��<�r\�Ҁ�cƘ�����,�ʴ��y�2�N�%��F��^��N����"kIi�5�Ch
�N��TI� ؁wx��kP8o�o���;�O�i"�*�9D�Y^�E|lU���������)����G,�9B�x�|�D�:��j��m%�v�H`$E��A��Wv�LR�8M#",H'ߚ�d]4J�2��`�xC3�.�Oe�`�!z�c>���������h����K�?
�RZ	R.�d��`j�R}U�M��{�t����?��0d<��R����J�Q^��� {BӃ�o{"lJ/	JQ����7�ͅK�U2���@$��|Z�Q��/@5�$(����$?��_�H9u�-9���H��P�SJ,�)�<6���1nfza���O!PP��<���x�.-���LUh��@@v�&6BE3B��<��of�̐��&R�tکZ~K�v��G9_�'�3A���K8�I}��<�m�r:6�/L��*nv�R����s����[�J�9)��N y�|�`����`a|�=�r��&D�u�Ø��Q�)E�(��H�����+�^���ٝ��ִ( L�ވ�{�WK���N7���n�d ��}��ς�#8q ³1m���>Xj@��xk,��_.̇�{ 
'\k�>"Uތ�2*]�q�B
s�`>� ��Ϲ�h�\��q��t�cj�@�bN}�i���<q�*�/��\��֟����l�'Ƣ��5O
��|�<u��փLO���)�IZ�\+����ިEv�n[K��5���I�^�+Ђ�ޖ��J;�ϕ��(���bx�ɀ�B��SdlI-�DZ]'�Q�]�W�}|]����:!c�VG�4˯^?��?��Z�Ɋ�@c�h�W[Hc�\�+[��y��Z��/1$��� �ixjàu���/UɎ��YO��Mf�� F��%���-�.|#s�r6�lW�� �w��A+n�a��=�ѣ��������`���m1���:>�y6te$f�_f��]!�t��;�r���M^�w�P���1gi��$
��]�L�1�#�ux��$�A����Y4�@�3я��ϔ׀pau��eR�Oz=��:�"���u���ґ��%)<jn��A�!a�!ł���k�ƽ7�Q��t���ET������_nzv�.����4��O�eIُ�;E�ϤQ�k?�����7�s��sH�����
3�B�3X.�`�/��6.����A�:xJ�)�0�%��Ǚ�6)`�p}V�&� ?��8���e����Q�-�;H`�?ŝ�~��� ,����Lf��)���B$�؍�+���Vk����JDd䛇o��:�]Q�P[�<�P�,�{��9��ۈ���zP]�aB�&pF,ķֺ�N�-F�$.샼� �@��t�藗�ާs���g�nM0>�fJp��\��q�T�&.�$�t��-p#�5J�Y0N��=���`ǃ��}�_)�c*i�R�o䋣�齸 Ɔ���yO?��NB0>�g|qUN�����Ȉ^��|���ga��O$|�A������S �,Ft�9q��T}jVt�5	~�Q��U�����<~��S-S��F��3�:5<p�{?=�~d��Nt"V��2��x<����Y`c>���=L��|k�`���^����8ɝ��a���>3�0��],�)�c�3.Rv��7���]���%�[��6��g���U��b����}t�9�j~�����i�>�����i_�Njf�պ�R&1J��z"'����j(�ՓF�PS�]q�b�Tť���Qe�Z7�7�;���A����K�1�/g�)���.�4�܈n��-{���e�N�D x�81��^���u*f�U��yi�#�`#x��r��>�����%$�FIH������?�v�����Z�DZ�>ڡ� w��K�A�h��@T��5�\(���7�g����.|l1��5I�LϧwZڭ����O:佢�����ﰎm�]�N�2�#~�vʢP��48tC��yb�ivk��p�� O���"G�͠�~5��aO��������ƅx�Yw̢�Q+�a�3n�';�5�
�s�bM�3I�Ef�m=�H�D��Q�C�'0�&��PR��0��:��D9�����ǯG�N{R�pQ/\�n
��3���X��y�$n�w'
�q�V`������<�P�f�-|ǋ"����O��KUg1,[;2��B�dU+�f�hk�l`��T�آ�+���6p k����uI���W_��G��)�8�R�ډc�����L�%ʐ��`S����[nX\yb�M�]�9 ��U��K۶%B#��6�D�Kg�rY��:Y��w�9�����V@#�q�ES(��a�Af����|N,�����"��H�}<j"�nT�,�/��G��_2 ��y���P��b4J�1^�`q������k��`��{-ъ{��y���O;Ӭ#	��bK�$���71 ��q)�X�A��n~r��B��И&���y�:�Vn�1�2'�v��XJ��ȓ���q��}J�'�e��4�:0��3�_��Z�).����3��?��ƛmp3����A�4�)AݢKO9���/b8�Q.��_�ң%�ح��N;;�$V��E8��L�[�:wKVF�hL��,�Z2H�,z���F�ⷠ o�X�:�S�����c.���%��Y��q�`�����8��M�� S���K�ƒ���h�Ā�V�	�斖.B�?��@��Q>Xf;������r7�_0W�.8��{R�E�E}��`�c�^q%�g�ަG�D�P�����٪�(MD~ !v���w���L;�F�2FW����.*m�]LX�!�;q��~��Gu6�%��E���N=Y����;2�P *�'��/�҄K��|��X%8(d��'�Gm�u]W}ʄ���$y[��txb(4���p̀��f٭;;���#-(nօ��5������`��y  ?()d���C�v����l�N�I��LX5<->M��~�]����xԭ��&���n�ٲ��J�q(�ǧ����6��zA~�O3a����9	Ls�G�TS��h˺pjtu\>0�Ӈٸ�n{߰������ �GV'��H������Yl��h�n�bs�7�����;��A����Nε`Pi���`���;��wa9�gM���>tI優$@pmK��h��dF�/k�LOӇ�蓔���!5�~g����GYPt8d�q/G`��Й���{�� �Ay��w�g�Ξ��	�Xq���d����#TdmJ�TB� =����ȇ�7��96����3j��_n ܶL+A��t�s�Uz�V�Y��Y��A,��h�:<L�x�u���_<�몖�a��I�"Kn��0�U��I%5$�b@��j�wF��#E4+��=F����"v4k�ꊀ�_�x$�����~�߆s�������w}]�*�Or��� ��ev;�J �ֻ���>{�������`���p}��s�������W}�����|es�������q0�r�"S��fp%�b��M����� p`I g^q�5��������@��Y-f8~�_�ʁ[�9��kT��9�K�P�����d�.m��Z��yH�q��{~�7�j����1>h�p������_Ѯ���u#	���Q�;"�\��yl��j��R�t�a2��٘���H b��l�*p$�{5�c]�l���ϢS�������7\�'�T���t��o�B8�6��
/h?�£�*8���W�ub`#AM�-�'��ۥ��V�ZعJ/�`�����z�t�Ϩ�@l/��uX��nE�1��K���Pc���`a'x��Q��F5�5+��[�fJ���As��o��2\�޳)~��+�;Y�l����m]�`T$kx�	��io��K��<IR��_wڬSu�O�n��^���@�[��oW?fJ�LL.�
Pu��q�3� U�ˈ�&�jzV��G7�@����%��oȏ�aظ>n��H��%��f����-�Slٟi>�3��i�'�9�`������Q�ƪoҲ`������n����j	�l��PW7��j���p�;����EXo$��2�4�F�����1��ўJ��A��{�g�z�fl����a�c]�����8��$�T�������w�<N�4��@��}���-���h�C��0�����ǋy~a�@�66�I���|E��j"�8�)f�CE�[>Y�������ëe�-n�y�T�b�D_��C[�Qn`2��W�$�B'�E)�۾�*�N!
Y�����J�$�[�x��%�VkU�5#�|���'D[ֶ�j�k֘����G�,���D��瀜5�X�PPF�ԋ��8Nƭ��Q.N�v�:b)�#C�d��CE��Ԛ+�+��/�>���`�[��F<߆pוt�}%��gP���Fg��q����il�^�*]I�s���>�d�G?!�K���U۠�ք2�9DHH���kL�髪�l��d�mf.
1�;=<ԒK1�H��C�v��K1i�������m[2�h�Ne�G]G�i=G��ܝr�煈�=��F.�ן^'A���J��Έ�����|j���Sݣʗ</%^��Ԫ��ł��M��h8yʀf��h��N6��7��"��KI��*����(��Ѱ3Y]�Ho�W�"��Q����8iV!�s}�Ey�B�[|�A������YWÃe��K�
#s�s0W�^5�jܓ�B��[���X�e0DNS�
�Ŵp8�iDQծ]�W8�ْӍ��a?WH���~ryzc%�iO24��N�z�jL5=�!�]�_[x|�!��73�O:�֔z
����W6bx,Ԙ��th:�E��)�pGE��y�����_�z3u�h|�g[h_�p�����8��+�����y�S1w��b����y�����'��Xc��R��!��-��q���s����X��K������:vB�pO�7��-�lL���L�����o������WL���L CQ���4�o��� #��bn #�G����~֦����W�Sd����N��������׫;��Lpp�q�8�i����%��-0��Ş
W�N��#����� ɞ>�P��y�bCSx����>/�R�7rg��ysCW�>����x�����x�|}* �ŷ+g�U���;���yL��m!7�z�{�%Q�g'�"t_S�f�ď�/����<@	�lP*�oӻ4�b�e*�sm3C0�Vd�/bC'P�v�ː�gU�yVR�:����Hhf�<�8Ј��X��n߬q��ę+�FH�]'{��Cs~܂�ݠ�zD�nK�1��Ƅ���s���B�7�����ȴ9�V�i�bP��t�$i�j8X2~N6��}ZX?O�J(ۇ,փ��e{�K卺<q�R|X�42i�F���KD��u�a���HGMT�h:	��C�po�����	jT7�G��`w��%��p�F�Ɇ��@�T�<I�	�w��ʲ�g��L�ړ��'D���� �X'kJ-�o&�h�Q�i��j~v��-�ɍX�����f�*4b��o��g�������kG���B'���پ��y&<Oei'�̱ؐ�.h^�O�s��E_�f�������T�ڋ'�]XZ�lj�y�h룭��]i]��쇴d�|����*�	.�
q+�0«�A��������
~H�� %o�m\��C-cr&Y�p֚z˧��W�7(��x�n0��.���Q�s6��{�*r`�R��ϐX�[�|��MF��kO�Q6E+3"�f�b�l�V��ݮ�Y�����C�56���
'ZP9ƶ�N �5�@=l�Bg 0���1AIu��H���dƕ��X_��
u�u>ˀ�����*�0�PJ�:ᚗ���U4!t�	��Z����/�)�V�f��hZ���1�K�j]�'����6�]�����-3��N�Я�
���T������R�����9cS5��m&�gɗ>n�譢���Z���HE�OD�I/������X�TݽI��^{A�g�|�5I�������gM�ŊV�J�� �޿!>#�Y��9�pr��iǒgJjk��/A&4�+O��
�j&���DV��%g�Cg�ic�~�)�6$|�����O�U'P�<��c�(���O�śxk�S��p�ra�(� B���)�]ބ�;��v���^����X0B�T����!�!���CA4R�:�[U�/!��p��݃��e2�[�ҫ��~�}��z8����ֺ���5�v��> �b,?�!��!��\��6���֘���USx�b��>Z�ZT�6ec�($,n��|��ǉWS2��j�[�ᨩ�Ux�\���WT%T}=�F��e�ڨ�Gc��qNoe93�����ew��jCIA��B�!Y�!!S�{�Z7��9|� G��r�+v�8�PO>�m��eg�[P���Q�5�7�Z.h��K�������Cq�a��6�3Zl�p�J=m�e�x0�;��lp<��>Iw��@-��^�|.\?hz���z�Q.��o:R�f�����E ��p���lo��B׿TMY�a��I����!`�s7������^v{�P��.Ӓ4مp�T���,a� ��|�Ռ�QT��j��C��&�J��)��F���d&�E^R���R���7Ȱ�hd%�e�t�Ax�W��m�jo�kY���ݛl��)
{#��K�L��&��h�Hީ�	r�n�!� }�/+�V~��EA���X���P����Z�
��.�X��7x��	��)��������w޶$R��ˢ�3��0�e��4�e���ঞFD|ֹo��Мm��=}�@����1	@Dm��A���-�0:N�Ox��Z���?A����<���,�A���L�a%��ac=^��]`}�̂��0��RQ�*AM�lEy<�X�(�."%��ֹi9��p���@���*gr$b�������U��������څz���kݪ�_�_�!����B��Ϲ_��:�,!z��BGY+�B� �ǈ.oR�����_ǣV,�E���c�bu-p�@M�+Pr�\Q��a����[������zk������}H	�$4h3�sY���М���{dbb���ߗ���爥!�u?w��J9�DwSfy�(� }�[�eHSu���W/�`���^�� ���Qe#5wy�+�g�%��bq��-#`i$Ve�}���L�bD�)!�K�C�AХ�Hl.% wb�2a����{OE=%G�d���@�L��ηIc�s��v��˭�����k����UL�X>/Y����ec7Jj�iH�gt�i�;��ʅ2������j���nHپ�a�JAU�y�����t�3Z�p�ͤ�+i���F������E=� ���j���k���=�Ӯ�Şo��6��!o4�z��#�|2�AP}<�~�\lW�X^c.;�xA�+�����vC�R��9�:sg�MB���و�i�\�w��#%-��L9�l�"�tփ��L%y�H�~HSߝio���$b1o���S������TGG������uGՊ!ˑ�p�BM��_���΢�77��.<q�f��_�gKa\�#`�%-]/E��Y;"I�|��.T��\���)ju^��y�a(ַ��V̕�$�׬��`��P��Ή�Bz��	_���as��т�%5���)��A��"��/��(��H9m ,I5!L.*x�,�kٿ�)��|��v�̘5�D֩捥��f�E+��ͩ�m��Դ�r���Ip��Q�̽�Q��ki��B�J���!�+��[�~��1lmY1�@
�\F:p�`��"�������O��5���u�)ᗪR�� {�Ie�&�T��s2/1]D&T�X�=��
��Èn�݀rs�^�D��V�O���:b�^�:M����#���Yi{�����b������0��{b%����a�_0���'�D���%�� N0h*(Q3-�v�>	obR�#��R�pɰ��m�Q� (;P��`�N���6�����~�ď��(����a� -13^�i�{?�y-ZGzV5�xNv*ԞZ~��/�A��߲��ك�;)xƐm3.Ň���-T�5����u�B'�X����0XC�%]u43����xe2=5}A<��͠J�wc��2C~��0��n' ߧm=t�<~�D��~�x�}��S9x��O��ͬ���@�'U"(�&PM.Y�f���!����.��@5o�癟,���;�#��W��✃Ϛ��?��OIc��� �1�ABF�y�>�HZϞ=/��RrK-�p~�T	C/[�{A�w}�h�����زi�]b�aq�&�E�<��)C�=`�m�'�u�7����:=Ϊ�t$��W�?��M�p��Rvi(�	�
`��m<�= 5��R��ܭ�F#�P�Z��e;w�t}��=A�`Ȱ�Z�-@<):�ڼ�u�ƫS��k��ݫ�ea�JcV�۞忋���Q�(Vt�0 �^d�:+I�8��M1��1vz������@{����������=UWY_��PiN�[�æS�JS�s~R,�?��)�0�y�/p���N���р[���W.���L߱�������Z���=����[x����g�Q#�:�X��Y�l�9��sCQܗ���8
î��_gt��YL��c���R�E�9������]�S$S�:���� ����/�����2%}3I��2�����d�	=S��PP��r�>mI1�&�E��X
�}�e#��;>� y����X�M�$��#ؠ��z��[��lm�d�2v�a�b��=�N�RL�P�l捧G�d

��}��+��'15��/y*E:ރ�*R2�(��x���vs�VzXYI1X(�x�e���Ű�oӶv�@=�^�j��Jd���WJ��tW)L���ܺ˧�ÊgU6W�S\�9kף�����}F�d�j�$���עB���$�ѐCcČ�T����%B䣥�s�c�)C�tt�w/*�I�E��f>:�s�u]�ݔB�!�*�@/�_fS��C�X}.7�8�2��W�V��!�sw^0�jX���\��e^Lk	�G�#� Z���wU)��{@�����t��K(@ ������qq�E~�L������.l��T�u9�}�`��ҟp�"��Bɫs�0��������;�xt5BNy�L�e���a0ΩE��g� ��Q���.��*gV��^�&�������0��3<��$!Zs���K��]:|��dU'�$|�����U��kx�d��� 2���+G�h\|\(l�Ͻ��tw�"�:9���|���o�F�c	>7�3ˍo�W��
��d����^>�W��WM��yF�P��E]�f�&W%�_�'8�tW^���(zK9m��k뒃�7���&���L����2��uR�Ժ`�۱@�C��T���L�Oښ��ImB�3�l9�e��]D��,쾟W�o����I�<:�ŝ CB���\2��
�Ow*>H
n�\,����äX��L�#	"������(�\����l�;'�] ��:�y�]�ieG=�A�R��@f��0wA�Z^���'9�)/�q��2���-+�9�%�A�}&-W6�����p�w)~Kv���f��؁nN�0�0�9܉1h���~�'R������+�{������C`��}#G:�F'�HH �~��T)�J�Z��ay���
P5۷����K5�l������o���H���*�!آa��n�_u#�#��ۼN:GE�3�h��#�@!ӄ�!�� C���@pjL=�>�� �(]Ga��"v/�5$�G�M�{��ZVa�9.��)1F�ǫ��Z�8�l	��Y5��ɸ�k��Y�p8�
g�Z!0�(�]�S>d_7�Rf�YT=�:�������`��^��&�����k�t�j'1�$~�{��_�w�4��}̊9���*� ��]��ÑwpԾ{$	���{r���hd����e��Ņ$�Z�fIypډ�M�%��މPp��X9A_���M"��������8��|�'���92b)��LR�8aশ�9B�C@Hzħ��� 
��	�1��_�sP���S��CgQ_��=�����Ht���n�)�y'�a>p���[9h؊�unf��qz��؃j�l����eC�y�Lma����������Nu!�����Dwi����Q� ��`�ʮ_��3#_�晱�X�g�UXc�{��h yzfKzCB_UBJ�?�>Q�yy/�ȠȻh�@]����CG	C�)1fk*�r�q�0�o�8�8�Ɯ1x�1I@� 7�j�v5��@��A��&�.�8���B�f��(�x,I�!�D.��m(,aN���m�hA�5d��u�U�6�$7��^�����8����2�2AY�� �y�z`�M@;?�h}�[��$�b3&�`D�/�0ɐ�y�\,��|Ρ
����{^�v�E�`J2E9ճx]����ɦIL�;UaNe��o�|fr�Y���WGn+���<Tѽ��'�����$�d�"�*�a�_��tq���� 默n��u��^����ν�K�j�qg���wj��\�K����bd�����`r���J�������Tͩ�J>N�,��ñJ1��j���+�1�K�5JkG�u�ƿmQ&|�gFfܠU$�5@^�ؽ�hh���ς�V��+C�8Q��0�s�V����T���Z(��n���!L�㓬+��r�>8�Y�IZ��«5��1�_"�U{4
@�3��!���W��nn�]��؟�t�/I��і>Tۤ�}#&̟ ɿ�!@1����P��d�Y�[:%L}���� ��]y�J ��n0n�I�ڱ:[���x ����':�⸽���M�oj7��p������]����:�G�>'Q����\�N�������G0R	еC���W�}$$\�W� 	2g�k׬=�~��M���Y�|��ulʝ�\��TD��>|��J���L��`&d9w���*�&b.#0��,x��[Yu�:}����K�WW�j!]���߯V*�����r��M7r���p���T���
@k���J��}�˒^M=y�Bf�8e��<�QD�8�Jx)c��Px�1�5 ������rr���=���&ʧ��E�M$�!��H~~'Y�/y4�G����-�u9�C�	)ð��P᎕y�)׌L"���5�VQ:��>F^O�t�S'�v��g��cY?�dTb\�� (�TCټՠC�pUBʦJ�W�i|	0���)4@Ʊ����"�j����V������sSx�	*(Hذm��H4�z��*���U�K"޹|�!	$�Ӳ-�9�^:�6é&��Wd�Pu���m�F���ց���wBE�k�H{�1���v�t���RT�P��1�@��_�gx;iB5�#G�X��
{�B�v��h�V�Q���MT��nG��=��@�m����#���E���ev�A����H�g�-��'�u{�2���	ȯcm"*�{�,��(J"��tZ���o+�W�RE�Y+�#�w�����[�����t�C4��^[�r(�0�Od�3jϒK�T��j�:�u�*΋�i?�4����R�wĘ)+�ݵ�D[�~�:�v4��(�]�bm����N��N&���\D�(t���һW:�oS��B�YV��"6U���pW9��nG\b�1P3�~�á��Y$��Nۂr�`�P���l,�P�Z�#�8WF�r>���Q~Q#�[ �)��{�ѨB�G_�b�l �|�e�w{)[�U���*���#&ϐ��-ʃIE;p�>��,l��[��->̱�-n5�D9�!>fy'H7̈�Np�K���ZȏI[6o�9˰ӕ=SYh��I+݂�����ğϋhu�P7����,�3L��������>�Pu;f�]�]�OG�(�����9Q�@D)�6��:��a�â�1��?=���gv�5�E6�7�>z���;#N�i:~N��+��'�m�I�i�L�XL�B$�X�\5�*���tӂs�E~K���C����o�p+S�]he�5���1��X��_��3�9a���9�MQ��%!���j?�n��F.�36}92G��ݡ���L( �F~Pi��5D��r��c�m����~@�����V��O���E/��,�:��:�"����'9+Ο�l
 ��Vm�d�����hq�P�������C�����[y�^幫�,�d�C>�*��|Au�yMA0(t?��N�o�|F�`x�0�)QY×��GW�P1@�S�}���0N��|�-_�oF�Ed���Sf���V~��
i�X��)�v��c�C�6���g�6�J�3�%r:��
7簺�k��]t��t^_��~�o��AZ��F����mf���<����'���H_�bp("���i��ѥyv~��n��^kjף��a�t��Z�Fk܋58�~�y�g�k��<��vf������WvS�:�������xZ�j�Ò�9�۴�sT�*M/�
�o�>EaN��R��6�'&�)5��"]y�������撺�+#*�h�=���d<�{l^6f.��?6�QUY�Im2	��n��O����}ٹ~���~�����\�V=+���r��
*��8��E!�.;�nj|�0�8�����	>!�����Z%+��y�k��c�A��� g� �ET��I}�?;k�N_���-���TG̠j[����u��
b	���'&i�+5�Ys�q�i�����.O�-��d��j	߱��@5c�<ky-�b�O�b���N$�ˈD<�_��@�N"0�����ʙe���tE��9�佻�]v�!�Bv�*`i�R��[0���q�~����p~��c��9%5,�]nq�;�S�W͓��.݄��o�<��|