��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q���qh%ws����dު�����j�"�^!P!�P�<�?��_�x��4#��hb�teSV܆�=� ��(�kSx^~�^�eyL�iTP�Y[M2�;Jqɡ��2 ��f���s�����c)���\�)�Y=vScXNt1$6���X�S���qmTy�-��9,��(�z�I��,s\��R�3tx��i;óH��_���ZD*��i7���<�-���q�<�q��� ��
�!=^�$�n�9�=�R`�[��m��'ZK���º�W��ȀI�xt�g|51<�3G���vlU^pڝ~�ʚV�G���)C_������_�c�x�+NMӑ*�ԧ���5��a�|=��t�w�^�E��H�F�G6\�M�MmM���n�:���;�H�C��,�{G�y=�Q��+�8��5�)OG��Gy�� R�_��A['P�p,4������qR^� �Xo����:�����/g�����Dl�&�hcr�(����Dܻ�rϙ�RcUb�l#1���}u!��?��t���6�p�W`�Q�b�����*'�	��-�x�f!����f	��������Vݷ�塚`#͙Ɯ����e<t����^J��1F5>��_�^�;͵n�rz�>�(S2��@��P82�*���k[�;�k� #��F�L��.���!�Q�d��?�f�7�#��E*��d��	�J��Ñ�F�$��SYpp:U�bX
i�s�/��W��u��;���h±��-�L�,B��⿽����s��{%!�$ўE�.g9�x+��Z�:�a��/D�/����2�D���3����=sM���7C�K�#��/�uȮ�SS��C`�������|���PrM��q�U7�o���ah,e.DK�k����Wd���i��ղ͌o��C�F�hE&/�hYpi��{o�`p��oz�b
�8�.��KZ��0��/}C��$@OV�wP�~�������T�`%���섰�8	t]M�α2��;�E7ɔ~�P�Z�Q]�Qv��?�GMdD����>JzbB���R�aa+&D�b�7uB�u�b��Sk^v4U��-�uŚN�}�?A�Fy��窃��#�NV����3�l��]_�&x��y\�������,N��gW��T@������2�Y+f@��Ae��d�W�}�^���Re}���u�����M3V���LP�[�K�4~T+avQn�I�0�͔Hp/c�ڦ�ˣ��ܻ3�!�'�v�3E��9�H�rnmk�fMH�~R��9�^�N���Y%(\�u���ϡ��F:Þ�vv�A��=�ó�Mk��J��pf�R��D�����Ơ����zK��Y�	���릊�������~�uZq=�����0�A��sd+��O��"�/�U{͑n�,%iI�,�o,���6�Ty��;L6>~�������w�ж���^b͖��j��A�g���hl��	+�7�h*U�2j1��Ω�@56��mmA���T��}�����d��{A^���X-.!��X4O%", �u��N
w����(�&�����؁AFR��B���74�M��9��v9���.M*��T��*r@���	�{i�g�-F7'\���iD�9�n�� ;����H]�[?��q�^@�͂�gq���10�P�_cz��U�Dl6\�Bxz�/Z�4��T2�$��4��mꮳ��苖
j{}%$x�����Vu�:����1$R�@-�=�ɬ�f� ��M� ��6����&��>	.�iFރ-�JRz�oOu���Hs���f�%ɔ�t�]��`9'&]�u��L�s%�ۤ �t�1�S7�d�4��|�z�b4a-pfT+�s��̼���\@9���.�M���vU��,�oB��N�W@&=�f��,JC�9��/��w���&t1Qn�o�!��]8p��R�
i�P!rj@UDE���t4���p�䔽�yl�V�,�ַ����(����l�9ҽ�^��5)�W/�8�ml9��L-�&]IL&�腃��2}px7z[QDK6cօQ�|T*s�A��q��>(k37�Z�_���Q��L"��G1`?�ڏ=%�
O�˾X���������ǿ��zW4�"��8U��[A|�4���7�?�˸a��)RU�߁Y�a��a�����߿�����(�<��.� ��ڄ���|�A{��]�{'O���yφ�15%�-�`.KŨ��y��՝8M����n_'����q�/��.\]��O�w�s9cM$�]��RkRC5uA���Nڒ$B�u�י	�C��5.U$㢅Ԭ�ܗ�0d�����w�;`�>�!D��"ss�>U+�5�$'{2�rA�rU�(%+�L�j�������bERe�6<� ��݇�a{{*��"u��!�a���V�>\c�5ƚD[�	�� 1�_�]R�u\ٙ��//����W�|N�}���t"d��E�v��w[H�����>%�[;��+`�?:���sH��.�kjd�=�R�������������Ճ@��][j�t��u2�
�{^�����2�����Q�Q��!�L�$��A}}�qCm�@]���nw8�v�*�<�<felSq��g<����W�qe2X��jG�Ԩ'	̶����6}��M��Y䞼/�R{�2u�����m�x���5�-C�Ŀs�U۲�\l4$4X_�a�ϐ[�C����a'�9�:Uِ�l�����2�y�.��E��Q6��`�7+K��@7x��	?	S~˼E�\�^��~�S��m���Bo"�۽���P��w�њ��t�f��@����z�5$�r;u9s�'[�eZ�ޟ�\�ҩ>Z�E�b!~�	a�e���2A68�̒�alF��T��
T����ju�������0d�z����u4�C���z���	a3�)cz�����K�-��܆�K�7��=����\�7M(� c�0�n
h���X4����.`$f��'��*�}��|g���T��Wo!����/sp����7���>������"�Z�Pg���!�eO�q�j��*�a{���߹��D�m�Z�H3�S�4�Ev���O쀿
���k���1�|�u F&er��~��	�ȏ����!��=6�o��F[\�f��A�>�k	e�Pqw�~@}Q$`�=��іFz���N��~��OE��W^o�Ydi��1E��j��r��s-�R�ZP���;����2��T�gj�V�N�~��:g��j� �Nl.T<����o=#oqAY҇3��J\��H��-5��ե��`Z�w�C������$�J�p`ls��������
]W;S��@�
�Dcw%z���F� ܼH�7UOi<
���6?(�����SsT]����'.�Ѡ���/�{%<$V�C]�"��g��niD��x���W�y���\#�)3Sq�����F�e��=4g�*j��wvc�q�|�:�?���_u�cK_����n����0il�qO��ʭ���E�[�D�{J�R��)͂��+K���C����%^�&�83B���H��r����އ��YX�l%�jP2m�A~;r���D�����ցM�~�d�y_Z�qO�S�3>�d�vGf��!`+�]�j_<j�o�!G�l�,=��v�w �%*NQX`d1�75���Mi+շ������aH�J%�,���f|�-)#Equ��X ��Dj�v�n�+�4r�.j�Q��O5�p�9;��)]�5!8��uTJ���\�w��5�1^E8\��':9�=�YJrcP�2�$�櫷�޸)96n��́��(���g���5n+ ڡXw�j|��Pq�S���>�#��L��n�m^[��}�v���*���[�n��RL��縷D��5r��>�w<:O�M}D���ǭj��N����J))�>f�s �h��\�ntG �"M@J�X׾+�:��������$��j�^��O�˂�V=,�Q�.���0�K�%��\�O�Ն���i6��,��Q+���~�aG�ǃQ$����@JR���G-�z(Mu���8��Y�
9�������Ew�ã*��Z!A����N�R���/b
B&%��1�rЗ��(���/��?�`krQ���r��Yڠ��Q��!X��Ɵz��=��s����Q�YG.ڨ�̬0T�tF�y�ӎ���*<�Y�X��"Gw��~�<g$gK5B/���!�o�B�,���ƽP�� ��3H����b@hx�u-W��1��qS��3�>�-��Cb�E����vS����Y����`�[P��a����Ŭ��F������Ǜ1e@���!�ϹU�}[|©Rֈ�H�Q<�p2<�9��v�S�u����_tA���{��!`�
C��aBf�S_����j�TA���+R�.���������w��}���x�8A���6+>(���A��_{$���Y)�tR�:�r���KUEx���8����t�I�A�0�"���G��U��d�P���ܺ�޾�zx��ꑋҖuU�eK0e�a�\5A�@�ւ�'B��[�Ϣ�u��[�����ӹ̴�<����e�m�8�f�[6h����@=�g���ƙ�Z~錥Lx�(6/�Ȅ�i���J5�Vug�[��� �_�ਵ�z�(�>�t�3�Cw�=w���<�W�ݹAB�1�I��t�V�Q�U5����mSH�`�Q2�d)� <�1~�����'y�p��N0!�5:DH�#��@{�u�����x/&��ԸB]��X�8�w����\w�FNO�"�,�Mx�@��t2���v��I��/�#����y?�2�Gӗ����t�}�}OyeL47�~^K<�	Dc����!fP�(B����&/i�ZW�e�4��I}��q7Ӵ4LwT�z�����N��<�m���m[B$��Y�rn�,�zF�߭��EK�*���q=�K ����*�zi�MLMJ7��5�`�ߜ��hm��'#��d�B��1�vjoh��ui�)RH����K)�?dgO����H{��R�~'��,��0�I���8����<:����XK�9�m��р�[��BgV'���He=��x��8�$����I�'J}����i:D��u��̹H�P}���0�H�p(^.-XK�[6���5R��]�'�@!ȅ��#<Qg�mw��yT��&�[��ӡ�=���݋8+LŘ��uu�L��?��V�^o����6����"�pE�ܝ��T�Y�/E�%��냿�$!2��R��k��z�<U�ؽ��ڟ�m��uv�81�۟�����t�Hl�B���l�`���]�o_�*��d��ۼB�C_m��O�1=@�Z��Y��p� ��hF��3�b�|�Q�����E��n�[�����0� `|!@��c�ަ��̙�Z3#[����4�!�n�/vs�L�	GYo�uQ^F=ҧ.o��fݛ���3���9�aI]�Z��,ݩ�Jt�B��vBe�mԳ��@�[��E'V������Y�͟ >j���A�=�
���񮺇_���B~��w#j���	Z�X�%���ֳUMN\�$�1���_"j��1��/�������`�zg�iǒ�%���߀U��h+Qk `1Ӈ>�Hs,g�����{=��mK�Ԥ��*q��Em:^mYK�LI���@m�d�⅘�lsq�M�N�۳_RU)��H�;RGWu�����k���,V�RKК�I0
��!!���q.���zȍgg��a)�G��=#�V渧(6'}��;��Na��@)�v>���e7�P�o���}N"=�@?0��~tc`����{KmQ���&�죬�d�9ا�	��a��l�#�uZ�[A>-�S�i��f!�J&/�xac�6�����߷�LZ�cI.�ٴc�X���?�	Ww�"�NG���O+>W��23�f�@��?���aq]�&�����[Sv���aP�h*�Q�\��t�����\{�4�1��2�t
myt>؛�'����	�|Q�t�����,���jnv=���;�N�c��o<{s�j�+�U�z�����F��39���������t�]���I]��.CQ�1��ø�CAicRTVp��I>/;ĭ �C��ե�Z���}��C�>DX^���]�[W���d�J���/:����4�v?�Z�֠��21���?](3�޺�Ά�#��c�@��5D�M�\]
��r5�=��ٚ�15=L�%�z�z��*��T3�X>5��2郞�@��
x�J��A�4(P5Rp�s�v����2A�C��/�=�к�Uhb]�����Nw�� ����}��1�Ҕ��9�x�T���\�BB���������w��p-�8����)�!�Щ�·i����W^Bq{�d�p�6�����uOR��7�����m �6��Ɲ-�,!o0�ߠ��,���+�}Q�?��
�!���x�G���� ��= ^{G4�$���B��hIrWF�����*f��C�-�Rrz_�cn��qy�ל~����bO���a�⪰��T4�d�l���J���*���2UE�ɖ�8�!)�	
�}�(V��1�#{�as����EM>��ٸ���|�u�"�,�Wޫ8(s�!Av۶�������lcLp-��%@�ڿ��v[C��1Pmɞ�v��2���V�$�G��&s�S2��jJ�No�e�=V2I��:q�Q�Â�Q�������HF�p�)��*٪�,�_�K�_�6c���,H��zg�b�2ţ��(q �v�l3cI�MPn�RX0,Є��j$��K�q&��"�u�8�e_��o��+b���*n��7c�䕗���!_b�V�.y$�ǩOt|�}|ѣz#>�	����~R�=��;��D �U�Y��D"*Z�x���J���a@�m�M4��CjwNYS����G�;r�*RVE�������
pIő\�&8U�5\gP�%��;:�F~��t���_���`�(�=l�8�O�a<�:�[d�b}�A�����n�s�譭��_ތJP�U�؉�a:�l#8c��heA�8��9�����S�2t���~�q��+�i�ϥ���EH��69Di��k�	'�t|�n�sԕd43ϵz6C!.������1����f��0�܇�	��os���|��m
)��ԩP��I��;����c��������N�1�|wxX���ʶ��
�Y�Q�&:�ϝ>��jPiY�+^pOI���N���wV/{���.�[K���@q�#˗�_eCj(T��D��L==���%	�{\�.���M��n%�
�j ��Ƥ���œ�\��#$���/F�xX��s�;���?�A���QM�lKs�)�M�}�p����v���	�S�֍�NO�Lʕ	^��$� ���l��F�v��#2������9=��ֵ���Z �>��������߰�hA�nS(5l�PA1z�*��xs�A%ٗL`�6'��>f�T���}x�V�Oۊ��� I������$%���Ҋt��U�������]��#�y7�&��ՙ����k��#����gb�3��W|�p�3�6����	@{���+���9K�=���d�����|��U�#��)�~ږ4dή��)�� G}:�h