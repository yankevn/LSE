��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>�[3�W�ry�cˀ�
��$� A!�J��^4�<��(o ��ڞ�yW�����ķn���_.���)+� *: �N-\�z*R��h@�e!Q9
�}oWio���r����m�顖<.��J܃���b|>�c���x5Q�>���[��'Z#�����x>hQm��xteu��Fʱç��Y���������"v\�,-�1���)n]͝ˁ�#&��p��{�E}��ݍ��?ah��}����R,pe�S�t��J���?D�@�H�`�Nܕr�-�l3�מU�%<O%l7��r�,A0k|j?�+�E����a��^T�/���k���C�mީ*c�xU����l�1�b��	����1��l:���ӻ�n���b5\G��"��-��v����r
^��M���Q�{ǌI$���ߟ�Uc� v2�eͅ)��4�T#��0�65����do��lӯ����G��o�DJ���8fi��mZ�'��p���#��'�U���/�5]g��Q��j���I��e�k�^���$��0w_��A8}����5���|#��'��h����;s�Yjby�3��Y�@�'����]~��>�So�茙@���-Ȝ���+�!��B����JPJ�frl���+�t����-H�����#e�6+��t�#�?,�����vm҈ı��3� �q�`¹�Q$���IpN��o��3�]�A� �h;�n_���F}���.�J�->V�䗮���p}��8OI����r�����h�|���Ϝ�/}N�x)�r��c�/�G
�C�<�9X>n�5�-�X����9��w�"�D����,6�ᐖ��M,'@��܋�~@s�}ņ�xQ�9o�yfܰp�t���|�5�'q�8ʢ���#�v��Ԍ㳾�7։@I�2W>n5�=s2ƃ�b��x�!p�� �d<3�N����>-���9�X�eL�]#��״�Uvb5��x�-c* [w��Z/�����+X�e�@��A�Sр��}��b6;[}z-t�{�CXtx:Q�vW>��+RŒ�k>ĩ�zq6d��Y"̹4��iM��p:�	,1ħj8y����b[U���(�[:�xjs]�d�x�7E'�Q`(A��rvT�x"M��w�3�e�O2F	ĩ�����H��2&�-U�F4bx���4i9u��k��z�i�#�ͤ����'i�|G�Yx�rl�C'U�=E�`X*'I��ApS2���q�o`����~5�Ov�	�H�6��-g�ΜN"k{l�p��e�ў"���qu>b��2r��|&�K��(Cx[����G�jIf�P��#j���ms8�p	��0�tY8��n�ܯ�8�#3�g���zJ.���C���fKWa�HW0��M�S�*�z�����F����^�v$�)�z`��T�iE�4?�$x
͉���r���*6�1������#����ER�x:��g#�O��:W�Ġ����a���i� �Ǩ��&@��I�/���i��h#7M܈��uq��	(�K��KR�  �9J���� I/6d��xCf��=�@�WoN��z����tR��澐"/�+�UU]���Q��@�Xw��<ތ�_z%~?�p�j��Pe�ƅ۴�D^�7�7M@�.�ӳ�9�5b$nW���u��{���˺[�h%@��ii�k��2�-$?�J�m��R9�-`�n�����#G�<J*J�c'a��p[��k�v�VOs�w�$˰���~J�#�v��u�U�n�`z\Q胰�׮<����K�E��f�+T�mz��h�e�v�h/�%�s���_-*<�C�jt�@O��j��Ϗ�^y�0ٴ�~5�̈�L[+�6�=�-��ժ.�hΞ��-/�d*�F ��������~nQ8�Kw���=���&R����E(�3��}6YOE`e5��fE ����̄+���z����7�>�4<9�TB�ֲ=�����L���I:`a�4]�5&1Keߢ�{���_s��*�f�����Z�	�>fK��c���=`�R��n�?�$^�XFa{�)�k�h��8�� �
u�������ǫL����-6���y-B�nKh;�<ưY� o:��P
èr<�|Q̫�ʲ���ӹ?����p���}����k,̬�\�`@[=؄�R�a�s�����N��P�X�w�p���F��=b�՜Bw�[�j~�y{�l�b�uL�G4��b��g��A�eQ�+���g�,����5�(��4�x��U(�|���=gֳ�ͺ<q�0��I�h1t�^�n��o�m�	q���pR��\k2��������=�m%��4�FP��=�^�a�[���F���a��Յ]X������z����a��������$=�3֙mg�R�)Pp
N��_�L�m$�V�rƙ�vK��!��@���I��O1��������i��u��0Q
�q��t~�ƭ��{�Z:�5;pM��j{r�n  :}�V<�}���9�2y��f����.��h�Pȋ�^���L`|�.��(r�@q%  ����> 4�����l��v�yiWu�1(R
,���)�ܨ�{ƙ�"��t�}� Jۉ�O��'�+�D?,kŖ���i��������\EԽa�CqAC���2��L&�ϟ�ͻ�Y�o<�^��H�RՍ�/��0`�v��3�"^�Y�^�� ��I�?����x3�IU�ʍ�J)eW�� ��/l)�x5#�L[|)�b$��P䍗N�Q"�?�2C9�S��2���bveT	�t�@�Q->Lk����^�1����{���<}k�+�v%p4x�����!%N���5E{J��<}�}ۚ��*
'1�.��+qc��cO��4�-�~��?��(�=j��>_=	_���,>�	��a"�{�M��1h��ش��,�*���[Q믮��z��.�@�}T�ȂK���q�|�	#6Z��5atmE���;���
��]�OqCq=2L�zǵ�a-� j�W�|�����HÂ2�F�j׵��ދv ��G�k�!��t�@g�����L)2�Vʴ�$/]��3�i���`lV�!���8 a��/{���Q�V�(��*vf�c��Zݢ�#�ē��͞RڃQ9]%� ]��E���v��eU�q $��7@ˋ�IR�:{tfi�b�f�rYd�d��?�]&�t�M�:��ٱR�Cy;ӫ���{b�Y��0��j1��}d"���h�㛍��g�u��&��0��_Sz�Z�!{iA�U��p�K?���.��X�i��Y���<wōG`�2M)f���E]�"!��[�\D��sBK`��P�kw�"v�#<����o��+bh�ii1�nL�%���yS�̴�1o��'|lo��|�����${��DA�Jo�UG����k����w_����Nl<��z~�!g�2/P���}�_���RaJ{�k��4\��X!:0��5��{�ً�@r �{�J��
���<�ĂM(��f��|�L�d��H�>�& ]��&1���g���]m�c���y��a�����J]_G6�K�dUUK9&$�k'獮�֠q�/v�\�U��o8f��G��$�Gj� ����u�0�� /H-�P��h˹?���+�;)i�h�y�X�;��b8o_s�S�� j�EYC(�ضEamWy�.e��Ss�1��óz�č�G&g���*�W� ˕��ә��_��	֖�� 4[IU�����j"%埦O�ѽ���1I����PD��}�
�D�<q��]���4�}�����h���	��"{x���$i�p)X:H�}qP�: