��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�7�Kۺ~���t��z7�; e�?!�C�#�In��E�[�Y��O���D���g�	p�k���4���Çh{�n����^�QVho�\�^�6��i�=���?��FD&�����M��:޺�)bo�)]�rx�-s��Z�:v�.ma�m|��@^�I���Sc�a6+J�n ���������{�����5Ĭ.�`��p����&���){b�u��/�X�ͼ+��e�?���< �Jn�jL79 4Q�qM���z��V%�"�Kf�eR��^w �p���OՇ�R�@?�|\<�y�Ӛ ���ų�a�/ߙ��S��_����c���HR���	gNa&�p-�2l�M����Z2�A�y+��)LyɭO��֧���/��	R"��J����t��c������{��WW��!&��'t~��n�>�J��%������i�qwnP;�SG�H4u��K-�����4E�5=$���Fjze��@���y��L_�:�1�2���-?�/�4Hܫ����Zv���Z�}���8����MVF�ܚ/p�91'pO
�U�]4�>z�d�1s��{��fʧ�J��i��J��<8�amw؁��o����h��p'�r�m�����a�W�V��-�t�"��$f�h���n��p@�<!��ُ�� _"�5.��;�)bxXV� C�b�{s)ӎ�\Rt'͔ݗQ	���[�ڼ�o�Ɲ���7���!fP4@��V.>��$�}E	����fda2)�D�^�l?&JP�61A��2I5��h���0Ɗ8HIb�"���B&���h=��˯��q� <ذ��e��vʡ�
��1wS{�|�_]����!�f��,�~��A�{��fJ}��֜[����0\-�P��A��G��E���`&7�l<0�\������y�։��w��B�&���b-�=����y���&a�����3c�Y*�uwEA�x ���@N63*/j�6�ͷL81i��,��g6p=7�p2v(`��s���8�j9�&��]�C� ۈ��	1�@�Ѿ}J2H;���HP�ws��c��z3�2U��`R_�4iN�٩4p�RZ��zu�i���|1�Ѧs���V��m�h���L=�mh��$C\
)���E���~G5h��#���g�I��Pi���3����5�%N�%m8�"f6��s}��I7)�q#���ȣ�	#N��Tn��������c���nfU�mQ�	V6�s���5睑�M�-FG 7��4Y��3B�^@I����C��^�S.�j5'��`�������;�^�nvn[��pUx�	��56"��]�x}�8v�{�V��U�@�p���9���V��<�J�'Z-b��Z���H��E�w��Y���S���
&�����4~%�����m�z��T9c���LI�!�4��Ǳ����Vj������Ű���Oʕ���ߗ3�I��lݕ�*#U��-���1̔8<`^E7��W=3�-�8�C�����Ŏo�����.nt��| ���L�|����
�)�MϨ'�}N�s�7V��;�$��,~C�=x���n�����<�����9R�9���~�&�'�����ӠI{��*�i�qF��+*��s]����i��!x����NC�'p� w�ɴ9���2F� ���A�8�>���:�<�l�qOך�VyYqFwWQ�;��9R*̜����#9�z�ݜ�����2D;�_פ�:aܤܪ��AԘ�.�$�\�m8\�t+hY��!Ѝ.Hf�!�g����0Ϝ�ِI����M�M�i*a��ɐ�}0��OZEBCO�K���Cp�]	ֱ�<E��10+,�\�n��&w^U �>~��b&�k��g��-�]_E��<F��JH:�b�]�z�'+$t��|6�0�۱�jg�ld��^ߠi���޶�B]#�iW�l>�^4��k��H���A��V��sZyl9D�-v6@"�J�!^��� 9��iND�[��������I�1����X9�L �U��w�I�-X�F2d��w��Q\�.�w��5��)n�������z�!4�uB@��ɘ��I>d߅����ItT������r�(��8_�n��E��^���R&���M�XN�ɦ��ǮVOй��]�bl�.�-[�<�{NNm(�+��V�`�d��R��?�}h�R�z?0҆ࢽ����\��|)����e�@8w� �KȺ6��ĸ�L�����$W��\�b�0�h�)p�ww�M;{�9�E��v$P���
���Z)�K��e�C�t!/�,�D3�0J^�{8�	�^�rh�4�������A�O����3o��%�(�L��Δ��03�i���)�T�7����8DVI��ѿ�&��pL����6�'�1�j���*�׈��0~E�t�#�[e�h3I�ɤ��x�*�h����0tgлĴ#���e���G}6l��!X(d��~զV���:D���H��}Ӎ�R��:u�x�J����M�t�A�ǌ��9��!��i��~��3X�I�&MI�|���*�:j���[I��X{�9��u�*�?�=��D/?��$�	mPN@k6E, �0,�=R\Z�8�2��M� ��[�/����s�g6�S�b�r-.���d�����J^kޚ��V�o��
5�ql��e0*�a�L�k�O��T��<dB��B� ���|E�0��戃 G�T��F� � ��3����l��SD箓h����>[�ߋh/��_ھ���U��Q�����^��{��P��@����P��������urL,ap\/�Y���}oS; ��49�ɶC�h�|,(���� aXC�J%����H�.K�ҝtv�wu�����4E��|OUl���6�*F��`�MJ��7#���.������2����0�=	4�y��ۓ\%?�h�rYP��\ ��Yt�j�� Sm�Sf�a��y��N��Q�c\��y���kEH�mi���)ܲ�.�]��f��ɠB��)�ߤ�e��hI�*���R�Ǽ��J:�UQ��0�Ѝ+*���Y��{��w�ڴ���䮼FVOM{�;�=�-�fT��r�y�$�࿬�n d,�G�be*UY�~(�|T�cب�VyMÃ7�|C@�`�6�����)g0�@A7�RY^�=�"�&�y��`)� ��b�Fm�.�����b"�HHB���mV��u���P7�4-yX��(���0%~�}EZ�R��)ͱ�Q6���*2�e����K)M�
�x����gc���JNě��r6�Cd�F�R_º�)({xz��[<����K���j�F)��&�5�;���6w��rO��;Q��5�����@W��l����ު��tg61�sR0]�s��[� �#ܳ��Ψ3T�y�	������~)E��������� ���CN^+@���j���󯔺j�	�U����&�F��#�l܉Z0e`�ԛ �������A�������ݡt|`���Rm��n(U��1w��('S/����m `��K�t8�e�M���b��|�e���kg���`|Z'��
�*ܗ
��L���"wtK���\����������rQ���.�qap^���j�.�'uW�G�L�"�}7� �)�z�&Dc�&D���r�D�8Oà7�,�9��n��o��� ���1�[�:l���NZ���l��k���#��7�7�A�'����	VZ�Ϟ7�yuU���j�1}h�������ld���4���~����N��H��1M$�W�<�+��b?� &�:s�:�o~�>$.y�Dz�Ct�A��mj{�^��K�RI��Ơ�մh�	i��*7Hc:���f�����6Jr3��^,���z��~	4k�j��ĽO1��[ۄ9������m:�w>��a��'�*������>a*��oI�
��_��Y16ԣ�n}��Q>Ti1���C4n���sj�����W���C�v��s�oq� B[L�yW�O�?�%�΁+��s]�d��E��˳�����l�Q�\�;�
@m9*Pmc-(}"�_®$�$��QE�DQQ�ة����wE�3���=K�q�����1�%N��]>!*��I',�՚��U�3�J+��K��ホ(���)��<���O-ШL��������B�����r��?��9���~3����7�3ː5�
uԧ��M�i�)�V�kT@�':Z�ƀM(q��|����B��Ӗ�K���0SA|�h�]]nI�����"&= 4�Gݡ�*Sʦ��f
^�H��l��\�����b�kB��bJF?J6ε�0����K�	1E�y�нe��,&6�F ���G���������f�^�EL���:O]:#IO��me�~vѱ�z��h���nۢ&)����rz�rR=,1yDg�t��]1A󐽅�(��� V��J��y-�x�����!Ÿm��Bm	�����yȘ��	�~6�[�,r:�J�66�l�'�&8�g3�S�
�=	�4���IѤ��`w]�u��ڂ��פ�l�fR��+�ϩ�J*�2���5�T9��1��7ೕ��8�=a�.�C/�d|���s��k�֎¸��3�����x��cd�2o�!��T����#����ms�����D�>Y���5���WUU0S��8�s��6�E���VgW�/�IPkӀ�"E�:]��#�F���ڋQ�}Y돞��{~��5q��RVqbV{[�o@5��G����HO��S��.�ǻ~�!��m��1f'�R!JҌX��k�(�fXmQ �dPD$H@��t��#HN��>�Tm���Rc������9?i�02�5��*#��l�R��^h�[�ň?x"��P5/�X���qj�tt8�Ν�����,�O?��󻐧���$�����L��&�����Z�)!����j�i�(LK:�*~O�Rݵ^�cX4�S��	��nmh�T�O\���Tʹ_��k��ʘ�$�B��Z}=�	�K� ���b��l���@A/���~��mX�;�{,t��D��"n�Ƈ�}�ߚ�j�����f13���n���,���7X�(�z��L�l��lVZ&�$.v��`�:���ր\�H`U'��~*l����q�Y��ݾT���z�*IG߃�֎X<�Ř�-�NKTҭ3N���I#���[�����{���#�.�B��IB�4�O?"h)��[N���K�GJ�t�#F��e���pz@�B����0NĀ�&���l��iC����o�|G_�.�Z5�B!0l~1	>}�U�HJ���,u̾������"�$�3�:U�F�S	����Ƒ���p��L�7����	��>��]�4@�l8�6	`�N�&g�g�Y�0�E�^����9<1@����Ǭ6g��w�{_KZ��|U0� �ΉX4���:��굮j3ON�jE��-�&��ڕ�DӨ3������3-�ݫ��.BL�}��ļ:�(����1��B��TU!Vm���ԏ���n��)���S�"�`�	�9��Qz�����";&�[�0o2Q�����ElfeJ��`���$�q(�<Mq������:ۗ<�Z��V
�F�A�����!���C{~P�W�c^�1�Lǣ��ʤ������V����G��Q'����������t���x�&�aN���]�o�i�V�k�;ķ��i��^)2��%���p$���~؆�,r�����#|�I;ގa�������B@1�G�cx
m�4x��+t%s#2��$b0x�\�F�L9<���9�3�^D�YjI�}�	Yj�AC���AW����hc��9o�ju*�߮>k��H�<�h��m��D��5K��M���)ѧ���>���u+�q����|�s�\9���ˣ+��yՁgA��H�k�G=����x~�NOW�[@���Y�❶�̜g�j|��i��0s,��~�{R#���4}��"�-.�������Db=}�o�������ĵ�H�h�|��v������!5fL)s�F�[�jڳ�z��dc\���Ӎ.��(��9��k�:J�f�.lf	a��4��S|rcK��>0k"���S��Ɩ/n9�#M�	#z�!�B�5�Mg�D:�m���|ρQ��t��:q�ax*N�Ԭ"�j���P�N�N�T8�4(�����A�iq�/��e�^̈�¢�2�.4�-7�sOx�;��}�k��u�����i����(I�b�S2��}>J�:���+2ՠ�W6�#��U�`:ײ,�h����Ķp�{��o��:����r�H��r�)�L��dm�)x<��f�����bPA��
< |�#�5A(��5l�a��g������\���^�^�t�"�o�#&K����4-F�����7�A�����{
O8F���	�? (���b=TJ�-�����I�EU9����8�6^4w�G�U �˱�>39+���������ŕ��.&�X������K��Φ�9���/�@�N��}|��գ=��?�k�jjs_�kz��� :�$�X7�1'�Oz$	DgC�85Eii� v
 v*��e�}�N籺��K�,q�;r��]��,��ͻd)H���Fůj����!�	��r�E�&���:���+���P�����C�@FL��݆G�s_���c$$��l�������6,�(�n(Џo�-G��XD/ъ�%i�!mQ㳍ܔ;L���2�7�oj��0�4t����(������67�e���e���U<-��C�;"vfp�����C<�εy���>.p���X�Oצ~8��Ҕ*A�����W���o2�YG�~ڨ��G�����0��V��'F)�[8����u�D\�GY5S<u�����ș������]��뛜H�2\���9\X �x<I�q߹,hᥗ˪4���D� ��?�i�!��� *�$���	�Mz��tz�삧�θA"_�h�d�
0�h",P��`?6���-�d�@r�R�d=e�2'g���@�;�L��0Zx�C�gG#R���Q�{C���W����˻�-?/����6���v~B�+��馛�ul�v+�����gT!�B���j��b)�3��{�n��3묄R�h��L�%��`u)ȦF��$;�5�o�'z��|�{�y�܃�uKK|�
����|���E�g�Ga(�����4�0y�Nn^�^�J��E�C��i��O# mʋ^��`����B�Ҏ=X��\Eŗ_�d�5�e��v��kq���)�na�ծ�Y2������P|c�fqP׆������$���ob�*�G���	�|������#�M[~t�<��C�������AN5��Dq��I�����w�q��dy�r	n�����ƛO0B�Y�����}Ch�çA����6�t&���� ��U=�V.��y�ف
k�rv�m��e��9��� F�I�=��WqT�ܚ�
��?R��h�F��"�U~��`��ڈ@Ok��5u������Ӿ2��D���}q��o��M(W����ȶ�������:%�>j,F��,H��E����Z�@ֿ�nrC&�`�#�O2s�A�l�}�ǂ<юm�����V�iic�o�3.�c!Ba��2�Ğĵ5 ��2����dz�߲��Q���C-EϘ�5�����[�/SC�y�V1e]c.���2@�iYv�	ퟳE�?�~���4�;1�I+����A ���z�)�v�T�$U�0[���3x0T2VvL�<��Z?�&��F�d8����TSW���Ğ��� l����f$��&T�����&�|
x�),2��ާ�Qy�%��� �S-�?��ِ	LZ��k&��2yNT��m����3�j�
�1:�%�$2ۺ�0�p^��L`���o1R� �fЮ�k�����.ݟ64�)�h4���D> �U�����	�iI(l�Ŷ�@�xV�>ֶ�+?K�A�tMby&�Ƙŭ�cQK_QR��;��S��4Ⱦķ�:N�h��Ꚇ�"��.i�7MB��S�c� /���D��Eݪ���m�*�IX�3���gR���Jwv㶏:(%�	D�p� m[����,�t���>�$p��3���Eho�]����فHn��nULew��<��)�f�P�n�i����b��mՍɍۼQ�T��-TA4������#��P.І�F�