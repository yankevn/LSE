��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2X~�*���O���k�<Ζ�?
J��I���iR��eϴ�J�Ij�Je�V�e��JB^ �9�E�|�h,����� �������c���k�zbr���A�5b���J�f�"UP��"� ^$wW�1�t�Ў��	�/G>�ڇ�[mȺ��j���K�_���)ϕ��4�����k-�mVs/��͆Cw�$U؇�/4dY���J�=������ ��e[M����
㌞c��|?vNqs	U�{)�ic=�$s�o�����F�/�������.����^+��t�7I�ΏY}Ҩ��)E5��'K��z�F���40�m��G �d~��e�<8��a��d���J�A�i��4�[���a���~����Pz��������*=���{��Mn�Y2���}A�Z�R�+X?��
��F��1�
 }��M�t�ڑ� �-��֧iյ�A�kϟ���f�h	 K&z;���d�IX����"d�TM��{>4� ������C"��U>3��K�;�0�~˗DO(�8	7�<T:�H��(8���v=�yX���^
��>2�U/�����T�9�\�ԍz3�g�.����\ډ�L���n�G�\��F���ډNR�Uxǉx�.�Jys)��@p; 	�{��#2{�u�B{��<ӟ�;$������;2������(����������#-�L��	�3�0.c08ʑ�Q�`F�&������Tb��YR��c(�P,d�)�%Ar+�]8�4�h��i6����R���}�}�'R��D5ɐ%�+��]k�1s�/��z%F~�h���5��)O�6��}�ށ�TlUx@�]�3Yd@\�C��5���ѧ�
%�Á�H6\�\c	�C��f�b[�P�o��=���!��.	f�ḵ��V5P�p9]��|��D����Kۨ���W�h:�3�V|�g�㳤'(�YE1*V����L�x��G�[��Ӧ&լݫaIC����<�:���)#�@����^`�^��f?5�C/8!Ia��W�����Z�����7��:+����K2l}�`�LꚀ�'�Nt߶>Z��Jz�f:��I�������zJ�\��Jk¹������
m]�Ta���t�8��v^�F����؄�jd��3�����*�w!l
�i.�	p�Fv�� %ܕ�RX:>��E|D����_�"ix���|�8X.�
D��㥴j�8�TI���O$XܞO�H��NnÅ{��Q��j����KBf��"���� \��,"��Ӵ��EB�_�'�݂�%�PZ2�%V���2f�f��??�;#&�U�� z&��i�s��ƙW���0+8\F�/["�EN�
�yw �����Θ|k���0k���2@��?�V�يC�NZ�7gM�p�E_ �����4e��v�9��� `ޡ�L6��_�Z�4�6��1�)Yue=����罣��& �S�x[�3*LE���	wy��.l3��p���=cI�xǕ!�\d�8�v Tkͧ�s<�4FK�V:I����"�D�D$*QY[�v-��=��[��9h+��j�ʇ�0�^[}kU+3Q���խ�A6���AݘJ��+gڇ��٩5�Ib���&#��;%Ż ~S,�@�$��2��*�quJ�8IT~����IgN2��8HiͿ,�K����K	��TE���N��l���i���E����g��V�8 ��o� ��!�23V*�<��qC�E첗R��[B�sQ��M�Gu����I���g�d���x��.���o+����K���_i�E��-Cuk2�j�h<o�� u��T�?#r��D��_u2	�L�o�2�n��'i1(��цMP/�z�a�_MvN!�&�'x��/��$�D�I��9�Q�Kl�T\Ss�M����F!v�y7h2~� ��3J�� �L(���Mt�;�M�I�����a��E�8'I�����C�|F9-�,{��cQ�+���4�*i�K�9���bti��,�B������މP1���"���N�_I�p.�+�DKI:y#M�v�p��QJd�С6�2���>¨���M+)b�֚~�N��]ubk.ϩ�uE����VL�7"���^:\s1f��):%��Z�����*1���]E#���,��f��*bU˿k��h��6z�`+��(��ji:QZ�!m�S����ڊ�	��/��Pԑ���u9�"5N���=
��9���\��ʾ%,��ǎ\��1�����k��������31p�D�nd�&;��~4���}�s�3�/�q����3Nck|�.��)an�����U������⌺�_�;��M�2�(�z|�ytbX��d�7h�_�]S:�xy���Gctο�hy��.6�į�����7<�D�~(`j�t�����K#�kgW�(_Ƕ�"��Wy�޶���գ%7���<}���QWA\��ʸ�f��q�c�R�˕J�[�I���K%�u5�M��-�92i��N����)شf�%j2<?�f�Si*�,*���F�g�L���g,�sOܿI��C]�j7��?L^�����
�,$�4 �]Y&���v�&�B�t#b���[����p��FF>�Sr�>�E���,rPZ������>m�_D<M����ӈ3P~�h1P?'��F��G�%8�B[lJi<��4���G�����5yx�� �fޙ�/���x@��%�{j�k�B�1qygt򂖣+�cf�d.r�¼{�V���5�)y��(�Sm�y���n�u@Z;�Ų�+�&Y�(���z�=��҇�cT����^��G`�5�4 9�?԰�PG^��F�L��N'=�M���UY�����`�0���f\Qqdx��8�q6!���󊻠A���]o��%��(��z�,%(N�r:	���Y�n7Ю� ��Qz�m3?1��В?X�;�O�.,�=����:��;�J8aI[;�í8t��.�#���yK�`��n��8��uv�`'�E�tީ�N%?������!!��^��A��ˎ~�c Va�u~SqBa�y���ȟ���
�����:a�Ct��d�}���<��w���0��|�h:�ۍ�P��1/��tϏ���C����o��&\��]d7p���EÌ�$7�{4������y�*cW��ASX#l���/}Y��2�>Q�@[;�t��Kc��d��Ct�=�AE����S=]��y}\/�?x�-�)�,�"@F�6/$���kl`L^;D�^��Ad:�ʭh�G�*Zw�5��C.��-��u���{��_U)L��l6�FԵwr2e?���9����h�G��5��{�>��S�R�o����'�n�2^�;1�*<YT����_9/��IW�	�p�'��;OĠ�z���®�b?�1�V��;UI�����Ƨ:��|��ٌ˞_�m�I�(�ꅀ+7�m�<��qe��:�z��,bU�KĸUs�穚ʲ�o�f8���O�B(�)���-��^�p}�.H�爟�
���R�GK�)+�(L$j��Ş2s;)�G�B��-^���e�N��y[PPA�8�J�YBűDU�错�J5�c���^����ɿN��viq�m%0�Ͳ��ca]M��|��a ji��P��G}���q�;I�F�����;�H�������dl��0��j���g[��-���U�]߂������#7!�o`~�pE�R��8��J�w������:�g;Q9���?m����o$�<����~o{��£���8s�*Ay���a�;����1N�-�z:\�y��(��V0��C��y�eC��8�@�O�XR�TGSy��M���@Z��)`��mXӧ>�/¤���u`��c�p�!uXV�BdJ��,��N��d�'s:n9d�5��{y��  ���@d��<1\ŖI]�9*ʴLxpl���Z����GX�����aQ�xZ���Z0�d�o�~ᛙg���8Q��v�D�(�ե�XWN���]_��I�����9�]��i�1���(�C�hEI+e���H�6���!!�t���	à?3EX�I������8�Ux$0|H1��bN
-�'�<dce�Y�C��m���A�����(,UG$䒓�6��Ď���$��e�Շ����1�m��@IZ�U�
����;��F{{�(��(�]��qw�_d(=�u%!��Y��2O��-ҝ�͑ i�FK^�#T֦> �y��̙�������AFi2m4��3�6���g���՜;�|o�{�r�Q��,�\�-�I0�x�x�Hx|�&
��.��$���5��Y2['��iS|#�,̤���	f�K�3��J#K��x��K�J]dC�K�%�6Ax��숁�l͵:%`6@{H��A��v�����lmf�C���oW +�M�\�����v��W¨�V\~&�d�1/0�&1�g�@����D��QR�3�QF }p;��ן���;�?���ϥ(�L�ib� �Օ�AF��!?�b}�mkEok��8_�����H2�"��e6�I#���dP�b�*������.64���]b��J��⥱2���&�ǐ}+�A��x_��b�FVMAM�rwe���:�Vr�y]�����4�P���� �6Ը��X�-�����-A�H>/�u	�a�F�?!��b�ɔ��+bɰ_�Iv���
D� l�;��1�7v|�	��~�$K������_� �!�a���uL߹ĿR��uyB���?+p:6��H���.�Wv�,e�8�tv�S�
�����?պ-��Z{t5f�aF�%��'6��`S��TP��L�H�����(�=��Vt�`�}1G ��i�vd�N&�$($gJ�w�=��\f�-���>MaD]m)�9���]�l�F,ۡ�$q�=c�Y^�|�}Mv��<u2�T�܏�8/���n��.�o@ˮE��}��[Zc��kM�"D���H(h�:mYH;�����8���:_���&e H�.�w��|��2f�-��Ȕ��u���?�B�����7��)R�ށ�+��4��d��I��G���!E
q�Ps;
SL�p�,�C���J{��fs�*�/���Z�7��������d�2`�����Q��>���e&���&����Uܲy�S��W]
2��i��k��[���n����X~��<��P�&�������#Yl��cG�ݽ-ԗ�"��_u!�6�*�k�Sa�]��|��CNQ����Ƅ�)��J�2|	��@�B:8������g��B{a�f�x��[A���4��@��g��#wqm���L�a"0,���Y�Na�پ���}�����*�������}��w֢��AI�\�;�8�52+Xh����Bf�� uϰ����7�G�:��k)C�r���y;o�"OsG���R�Lߕ%�oIL�s|@э����7����?��	ýt�=;��g�絚����4�A0�$�	��d?��։�be
!>��� ��MP\:�#$���o 6�AD!ݛăg�I� �`aj �P.>ѭY�������U'��!�Hʼh�*pd.h�\�+��A��\��9�'���fr��\A���q��������&d��_�D�`;�� h	����T�}�Oy�W9|��m$���V7L��'K� 3[�M׳x_ʧeoB�@TVU�mg�t��F�ʯ��q��2��l�A?��JQS���=q
U����ĭ��O�uW��$��n��0�',1;݁s�	���(�c��9��n%���	��Z�����5
AZ �*����g�00�u�����tR)�G]Cl���}2hUVJ>>�3卺-��f/�f�Li<��Vxޖ��2�ч���ı.���c{/�m+k�zS���qQ������i4W���qM�M)�<����p�ҹ���.��ó	����y��w��y�	��[�2�2 �X�B��'��(�֬�_f/X��x�G)+�F�LP]���Xu��՝������̀��<4��l��"nk�j������g�zr�ǆP�V�T&�?��O���p ��tF�qb�&�C���K��[B�)�ila�'<��Q�>:�h�M~�<^[ШT�	j����#�,��tu�#����gs�0���4tC��10�Jp�������:���aa��}5J�!�jW1^������%eeC/�ДE����9Q��2a��h����T���4|.���w4XW8��S���/[������r��ґR�c}��W>� 5k ����94uFN�S 3�m8�m:ܙ[Y��	�Mo/n]�z-���y&� ��B�+�s���ط���|���}+��p��̈����I�rl�]����|Xs����< \��|�*���m7��g���0jxp�%ɹDk����^a>���x��vqҡ�n5AMR���]ٓ�6a�rp09���*�
��7��%���s�#�V��D�b����(�֡�O�A�y����5���C���$!#���M��ԍ�Ś$:�'�F�=�=��P)!ck돾Y�n6)��/�z0K�9z=G�6����@����?;*��Y!&�-j�m�;U���ȐOӍU�4�B$���:� �9�k��%�������]CԂ���Pv�◸�VQ�4�Q�_zPI��8�ڟ�-|̠��mU������9���?�5�d�P��G�=ԇj��lQZJ�UH�����"�kD��4���U/R5� w��#����
���v��u���|^O}b褑�/f��)�5�@{������wM��M#@�d��-�ĵqŁg>��Pd�⭬g������������2��f��D�3J
�-�X�<0X|�vN9���mWv=ѾP���%�����l��i�W`oҹ�p����[�j�ޙУ<Q��
�kB7=*e)S��a�������A�@�-�-�WŖ�E5\�I���*V���u}�e�1��D�'���:lw�_��8�kcފ�e w-1͈i�S �*>��U������Y��&��z�Nj��N�򩨇5��7K�GE�"]Xf%���ͶYC�+;�ڰ#��1�xT�A���L�fO�t4�@��R_Z����<>AQ0\�̂ �[�X8�#i'���C`B��.t��.!(�A� P�����d�L���f�>
T�;K�ef3t�s�p3���Y~P��8\�!B���eM���:��xv��c,e7s"5	ì�t=z�<�?!#A��@���̵gCf��>�Z��'����fL��AJA���}�R|B���i��iQ�Y����$�
3�	\��jZp7�v�$e�_��?L�Ĝ���	o��,pid� Qߡ~��5��h��z(]��ņJg9�f�`��o����+�Cp͵�p3�t�v�C�'(j��=�e1�&"x}#Y��MK�Y/���ꙛ	%�:]�1�)�$���M�\�h�&�Zz�')�A �3مl@�D�Ԋ�.�W�8L�5���ᓔP⸐2['�Y�j�o��i(۴q��E�mG����W�YM��.!�'`?3G��6,�eb�VhHb(�$J�k�2����@̰�M��^�[�x��
���{,�D)��O/�ι�l~����R������N��9���D0�ZYIVn�"��|i�9��X�i�E50?�r��}0
�N�n<�y6��WX��+
f���+� d�91�7����xԷ,����i[����):ͬ�e���v��{J�(s��K�g��O����ء Ef�&h�
��>�=�a��g��"�:3��KW�"K���"8)�V�TLQ7
(se�����&�2��� ݲ�=�7�J��z�Bɸ��e�E�MqUزT����+4�g� ��$8ҋ@?n� S9�X�)��P�k�ZEW��:�ڹ�p��w��&�G!8����zOHOB-P��K���h����ѼM�\�9s\ɜ@�W�ЎR@�#��~�mȆ!�B����g}��y_��p���������w:uYN�'_��s3��3�z�/0�YA8+륉 ��[ْB��%��Oe��j1�\]�[/�Z�:e�����U�����n�i�e��T�f4�K�zW�)�~(�t�ú����:}�a�}u�uy����X���m�+�����|��(͉�PA6g�º�(���-`���ߗpt.R�'��f!��7wϽh��Ah!������r�ب�]�q~{dz�S�yY�b�z׉n�R��?�؜(b>����[+��w�_��T�d<E!pO�w_����+M��v��?��K\�j�;x�,p�[���O��>��ZEB'�jCt�\A�����Ƹ!�9AG�o�GP�ߋ:,�[	���O2������M+�V'#X��-Z6�_�2��\X� �M'�ҍ>�M
<�l<���bV�	�Py�x���F�?B�����1�xe��I�|ϒi�`��Z�.���iۮ�3��R��-U5z�p{�t`�iN��$����l:��@�����T/��m���܉A�d.	
m���#��m���Dz�B���Je�S�lTu��y�ᾥ���'ߡ����V�ږ.�y���ͳ �=ĈzL��J+%����ĺ`��?�l�(�eT!��a܄�����$��\�"{��Y����@�1�Iy�>-�m��P2;�X0�O��'C�^���s��i��8(^A�j�1ɹG^?��6�c�j��[N�qi^�-`����@�yL��)�Q����e��V�/���ꊆ�!��'=�䅘�w
�AJz�Кմ�� �H���$e���¯���q	�PY���
+^�?�JϠ�c���PP$@�j�m� .�׈���e	�eA��!G��ſl�R�'RV��uMGI�ѷ�E�̥.�"�{�47�xg�$3t�O*]Ob����W��z�����jጥ�	Q��c��*�l6���l}�L��<�>+�3�)-{Y(����_�jA���cih7 еθ>h�Ǐʞ�8��D���s� �����ܬ� ��"����'lM��~�v�ON�PȪ��g��V�q<.ݭMC��^�ځJ	�h�����	���B[O���A�u���!5N�8���g�uA�Ĝh
0拢� ���=����M�4��N��puVa���[M���t%�:�p���
��Z��v�E(ݘ��"�
�> ~���Y�4+/ ����@�D����`q���nw��Ju�J�6�����|��o�U���i�3�t��9�yx��y�ԱZ+���A�=����{hJs�&�PKe�ޘm��C���φ��r�[G`rKw��jK�q��hu�>6?�j�ʺ�)Idyz*l6S飭�a�����}�cЏ?����H��_E�tE5۶kd��o.����9>�gѽ��3��@�5(TaYy_瘬�K������!8���/Z�	���ʝ���/��-À���kTX�50��F"�G�f^9��;{[����m ��.�1gPS@���Ih"�4J'2;{��-M���G�w�?򃉻�[p=��3�d�p����F�v�	*���'h�M���BMFu�<��V=����C�p�
_��5����F��gl�m9�0�	�D�*��Y��)^?�. �l��7��.��t���mt�
��T�VML2wƊI�+�=�%ƶv�D�X�M3�����@��"� ��(�����A�,EG�ѯ�n�J��;Z���;���jl�*�ءQ�
�b_9G%-.νG�R�C,�î�I�G]1O�sc��t=m�Ǿ%��JHe���:��C7������7F3�ɔ�s������j��"C�|X	�CQ8�[>4W}�Z@����+�s�����7��:c����7��qx�\�j�0k�J��P�?{�+O��9C[l�������b�k+����9�@�KNğ���r?f+��_h�B_U�XlYÁ��xsL�(Y~�gc��&k��d6 �l��� A����k�BW���I�A�|jL�t�P�!��FB���}����g���Cǟ�OQ���>�7TkSV�t\�f�T�ϸYR�yTnQ��-�}e$��� F�J�ROYU�/�N�Lv.�sF� ��h��3$������oB��S�qS��� �����ݝ۳��g�
rK0��$��<ޖh/�m�$�?�2��B�v��e@��ud,V��J�Z�5"����<M�(�`sY��ź�>����AR�&)=l��ii���>���uPz���B�
���dP~�:d6<Ar
�W0�U�In��d�������p�dF�bAN�N;>N~_P�Q�]��J�Zeze
^��+�k�z��N�O���!w�c�wǑ��●�'ui��۽�)= Ns�xb�c��=��,0Ȋ}tA7�]S���N5w��;}n�F�@����v�eeK�d����brn��8�?�D�eF�[3��Se1Lm�ѥx���vZ��g��\8�0C��3��0[-An{=Ve-IGc׀:����Exd�� �h�6ԗ-NST f�u>�ֿ����5Y&dK���P����Y�c|.� �����P�ū�P"Ԁ*fS�1/���W�����sS�0����Υ��P(i0��� �b�Kc2hezU=Co�A��gc(�<�\c�?��rn�b�/����bx��)m���0i��,��+���~���g��A�sY������7����AJ��t!j���bc�;�Ԃ`����|y��P<�}���썛�Bz�H���w��p&��A�K�{�Af/���!	���h�Ofn���	Y��+b�_�C6�x]!5��EҟQY� E��� �  Y�-����,u���"m'6
���\KCPDa��3���f��p��t-��3�����y����}G��1��%E	��ע�G�u{�@);�f�5��Rߟ�WSQ����iv
�m(_$�C�[���U�.@�x��gPRt��0|��f�w�@
Л��^Y����m��f,���y���.s���ܩ�X���0�ֳ�������;Q�9��m��\���ݚy���|W(7�=��&TD��&Z����ps��<ʟ�^�ő�qe�8�k(����A|�t��ߩn�^18�PG���3��46������.j����
�e&G�/R[���jj 6R�	@��ܧ�{��|(��s2�`����r����I,
8���|���v[�<eW,dڃ�L��>�+�|����	sQf3h4�Z��{.&��νny#�1�1:�����D@ư�|��&�;G�n�:�t�T�"�Mӱ�D�DT���eVJ�b���J@7�t��z��ѽ�g�����˶93��.��A��,͈c�U-���t������qϑ���V�M�"TC��G8�ߕǎD761�e�����{A���� ��l���Jh��Z��y��v��WG��̕T��T���7�N��w0@ei�?*��5�/Me
9*(��K��wש�bb T��|� �x��,H��0Ĩ��x��T4�O�L��[���o	I���y��JzS�{.� H�3����~���G��ba�t�L�.��l�A�����n-���.8��R���r��Bx�/}m�i*8��ڦE���*؛���d�?�3��]j�0G��Rq�j{�xV�v��R_�/�e	�(�c�D�>�7M��@�Fw����Q�/�킍vf��Y�_*y�R�R%�e"�kN�v� u��6�=v,=��U�MP����FA:��Cc�؁&<�׷��P_��Kc�}�s:�^���.L��b9�ĦKu�������y�}��m�7�%������ܗxIp�|��8�����?fW�w*�/���r����Z�8#��:���nV���(A��֭���I�p7�7J�hXC����M�HtW�`��u��n�wϪNUU��bKB/�Nc��xYNz㸔���c`1�3�zi��Y[�j��2� .�
&�ߓ��z?3e/O�JPF�d�?���,�e��l�>���Ð��0;��S��˛n��5%d����m��.���&P�)!'����vɕm�[������m�M�I%_�t1����љ,�Ye��!4=�G��x��QE�2j�U�a�|ǳv# i�`��/�#,�#����������Eշ�z��{BGf{\g���@�.?�W�����WLm����kD͇#�3��CYy�>��q �zJЊa�A.L���$�_��\-&&MK���Em��lQ�R����HG��v
��/�;f"l�Y��IsF]�7͝�ce6R�`1�2��l�����k;V�w���\�V.��n	�����:�5�܁]�tk�U<�+���N����^��S��0����rF���g�����q��3��T�_����r K��x�<Rc�k�}l��*8���X+H�Of@g\X�~}��w���(bM�b76�M�͞�pN\y�w9e��v���!O�Y!F<���':,��؅g�"D�Q`,��sM-���-� i���|��z�?���I���^L1�Oy�?�#"�X���c~
]���ؘ�{/��0&C@��=�&!���� kQƠM�*`�v�I���H3A̰,�pjU���%�v��mbO_�B�̧(}����a��$�xЂ�L�:!^y\� ��sl��{Q/(=�41_͜�K	���5�z�>ҝ��L�V�+�{�����u^��>��WB)��ʶ�6�iXo���s��##�ER�K ��R�	V�7�䑼C�Ŷ�t�lrODh@*<���5&p�%;�kܤE�̫MK;���4$�}�O%t�� /S;	0뺤�RΔI|�G�����Tu���n]�L�ô�|�R�ᖂ�d����j*�˝
���;���v����d<*��	{���r
	�LҒֺi�6��A�l�6v����-���}/�\��ܣ�0\���nd������U��pFn�r5A���f3�v[&&�j)��d�sh/�Adk6lU%j�v��e)X�$��­��tc�b�V��ʫ���} >���84��	va�</ߓ,�(�����	�^�0����ɼ��"�̼����T������r��;���r����,�/�*�_]�s݂B�#��~�X�e��d,4:��.�Elz�Y~�`�b�C�Hcjn��ـ�� �&+�U˴%It�����ykzm0�B1d�x�0��-��	�Jΰ8�%�݅b=2��S;|�ߦ��3���V�g��G�a�{h@̒�&1<�b"rc�2����v&������0��!qX��LU`��d�a�O)���&��^r5�5Hr\N{�C*G%L<�*��3����ȏ�F\=[��M[U��S��X��j��ǆ��</��t��;���+�ٽ���O��5��GVU,z��f�Z
՜�I���W�|0��w�tm�x&��D��9l�=��j��?�"���?��2^��
�)_vU��Bp	�"MCSL�i�N���u����) ����CL:�A�$*����a��="l���[�S҉bo�*�l$~�c�<�ɱA0��* ��Τ]���Iv6�^r9s<��q|�z��]h)B���eh�����O^��z��M� <s�.Ŵ�*`�9��9��}oT�V�rdPKJ�����6:60]y�$*����k�]j�.�Ћ�30pA1�^���!u+�Ar>���Z�֚V����4��y�Pb�I�|��(�������A��wE _(��|�4�̅��yE�/Nn+�!3��A��^�>���t4=��^����t1Ͼ��n;c�C{��.$hUaQ��i��C�I�]$Y��'p�R��+�� �'{u����Ĥ�]�rF�KL}
�M�EE4�5e�vU�@ۺ��z��m3��f�����_�
�㙾��w�оI���`��E3UƿD��Tk��,��%��g�}��}`�Hr�U$�~/��b�ꕧ��J�o���iTy��Y�BhGm��CG�!�$܄���to�?Rи���B�,]Y~���x���cscN���� �$7
S�!��ڇ��ŀ?Ѐ!)�6/�@֕_{��@��c�V�u���g�>M�D�/�+$uyȾp;�$]�x(�`-�.,�*kH�^��O�I��]{�ɨ�\h:E#��G�Ĺ�[�#�������O}11'�� ��E2�gIB��ץے��m[�\�l�x{��o!�"�ه`M�~����U�il�mA0�[�6�K��5��@a����+xx�jZ�� ��e�gw�yʲ��vX�V�Lu.�
Z�z�L�"��&$!��.aJ�71���Z�l(g4�~�mj�w(�Q�MZ �.����ةɫȗ�4R)�~��O�������9>�Y^�#$�5,om�Jt���}ms��$�G����R�|��#'�Q�!f�N͑Q �aP�{��O����#���^�œ��V���?��_:���ե��'R�[��ʪ5uNp$����2��@#�@���J�O��>��Fa��������z���t�e��lr"��#i�����0�0\�(�6R�l���ĝ�R��G�]h=�5�SʴY�k#��y�.�o��,�3���
�aQ��l�>�]L�%���׷�a�B�X`��FCQ��l�4�6��nn0G��9��B��/Pb���� ��>�ŉ_rS3����-��e��C�M��yA�P���lfM[��T�{�>8?�Q)���^���a��������t��l+%�mpp!}�'� �{��)=�\��1�v�z�H!����jA�5��W��H�#vV7���U:����F|S,��(o�'�췓,}�N%����P!1�Y��J�ަ���݈�eՉÁzy������0�f"�2������c�����+��!�������� ��+�.���oe�:�s�"I޶����C���vɕ1��lr�|*Y ��0�I�Y1z�V�g�}�[�y�z���ؑ�R��扷/tUMG��jd��loi�fh�Bx������N׹x�u��:���Z<-I��F4c��+���2����′D�FW	ʾl�{�V�rA>�gn�oP�s n��dg�����w�U\ ���L�@���Ɲ�i�����<�p%ȶ<c B��>Qr��>�I$U���_Z����r�(�ᄑ�[Ce����|vԔP�$�`tL��^������4ek�h>�|�,�j�yd3%`�j�:
A��GrZ��r&�4���]�����cS���_����q����m��6�U@^�48P�*��2��՘)�w�������7Y�&��f��O F���X�զ{����?�R����:	ҿ#�ƦnWʙ$3��8�	�����Q��Cڝ���3�:��RdR��,���J�T&5�ڙ�]_����"���˵#�n���4���Xd���}h3j�|ä X��U����wi�Q��/l�e
����aO�9�h�ۄe֭9���^Ro��&�LG:(�m��V�xa,/f�;"�!1��%q�@����.V�mC��?��vpQ���	��8��k5Ğ�����ɡ�x/#��۞L��׌���%��
��m[��]�G� \k�Ux$}�e���`q����2�\B��ѡ2�}�uʚ�0Z�}��̢�����p}�A��R�ͤ�|�a�x�4���F�a�!̳O�u95f���V���hW�r�<}�Q������[)"�Q���[��?8휘�\W��!<����(��@`���Qxp��[�[!�^�`��Y����|�]F�JO�T�V��{V"���ėi
�dΛHY�P$V��8��ڏ�"�r>%�J�u�v�*|��I��q˛-�6p�k����LLX������;=�I�$>�l�����hU��!f���`]���s�sv�CM�âN�ل�����LL�6�Wx��)�O��wm��F�N�t�m���DZ#����=��we彉�-؆��Û��;]V.����	�#�D���/Bn�YP��Qr"�:�%���&��X�4��ދF(�MV2��n(C��;^bG`0��s��I��Y}���"�K{08��������K����1�ۿ �����U�^�>L����(�װΊʵb~�����:�s����Wq�g��M����8k�n�s�&��͌�b�#;K�H���ߒ;5'��or�5��=���h��;�����������ʗ��@���,�i(y�]����خ?�)c?c�\q/�~�~�Hȟ���%�u��5�ʷ��%&��+JY[�)��g�yѧ5�F�@H��<��ǁ�S�D6�k��~i<,R����gF�)��JY;�?e~�l	���췐�t>~jKk����m�0CC�����"&;lY-�Ǆ�0^*G"���O����{�u�|��޿�������)�(8gk��S5xz��B)Xr����L�,a:Q�������8�Ĕc�8��D����k��R٪ԢT��H��ݤ͔����WΑ9��,`V[N�,��?�1�f���C��s�/�
�%&)��b���Xu��	7��T�p�-g���ܠ��l)�Fᮊ�u-�o�Lsg�h�
��47�#I���yF�A���]� �b
^�r{,呇rs,�}���B넕vJ���3��C���1��qp�xԛKA���wɈ�m�̱q��M1�{0v1��VP�.fWݻc�E�\���O�b �m���|�[�m���y�V��va��u�c�'�!*�m��Fm���J�ʚc��j����Ti��i��R���{(�̾	Ͽ�#ǃ�_(<�m{�s���3��)M.�~[��|��#p{�Zi@�{X�w����U=k�Z/x����
S��W��=����n��l:�@V�cwѥK�n*Q4��r9A��sUL %|{H�P�7i�(��EA�P������*i��Цy	Z&��hVmI�����2��4��:3�������#�[�̉�XC�a�R����U����K�G�n��{���%ϔ���5�Z2�r��}�^�K`ލ��Ãb��.���g;b�R�<��ں)� �ƴ�#��V�e���0<�0�l:�:�\�I���s�8��Y�&�H�;!�Y)S/,���;B.��h�:P�@u���\e�&ƅ�>�ZqP�j�b�Kn-����a}<�'��s���S�/%!��I�k/�t-H�櫰����s�V�e�Y�_�&搙W#%]���5n#�� ��F���d��ƈ(�?n44�h��|�ԭ���"FD2��?�{B�|�դf���GD�z/��y5��M���G�H��\��DX�VG}��
d�니�Y����&�A�d�i��Y�|{A���҃虌�ӓ�!`�y N�0���چ���|����c�������ofL5A�AX ��m������Nj�St7<�Fs�$�V��V�2T�4�&=+��N-P	��~����Us�T�^�l��3/�\�@`�ƲjS�󏲌�qΧ��n�mb��ݨ� &�N a��z���V�뭃�D�2�0[P�V��:����\+f��vܱ�7հ�e���}\���Ϡ/kc���p�%�����:U���Zb�ܜ���S�װ=�@{1)���E��>/���t���եVB.l!	[�����>���@7�5/E����Ռ��%�w��DY4����f%8�����L��J�$~�})�G@��c���o�>�G]ʻ	I��m�{���]g��c~GuU��Ä"!�\���j3t�H�I.�4��۠�Y$��9��%��,Wܲ�U��V	P-Mg�C����Ê=YXώ��+h��XY�rr�tY*�2���|�Y�>��D6�>9Ș��q�������M�Ι��@��rVB䥩�_���]?5���K�U��g:S+��9�j?��^l�]����	g7X�x�m ��ī����߻o�[����D���95��\\%h;'R�	`���1Ŗ'�59$��	m�E�o��G�4�B)Y� Z��#VK��w��
h
��Q�(�&��f��I�Ea�S�":zd���c�w/�?b`�|㴁V�gFs��W|=d��z��j��@�f�Uߺ".e"��,��SթHQ2�J5j G��{'�)���gF��L�#�'˯
<�.U� N�w(k����&�d�Mc�5��f�/��ȹ1��t�����m)��:%���َ-���1LB����B����>c~�#r��ѓ���º�Hh��p��������@7��/ejt@֌��
��.��4���GL`A�_��-~G�����j{*Ha_I�%9^�ҥ�7�*N�3!���骆e����?2��N9�4��G�yg�܇&��қUg�zq�3c�L6-6�KJC��O�5�?�ƛ�8������x���k����I_\^�moޟ+�����eK��� "���1�f�w	�d%#z���AB�T�RTg��%��ح��ܝ��*���)Ȟ4��;�j�/���8)��n�p��s�`�G�����Y�B[s�R�Z�/�HT={$S�1��n}��4����z�;(�`��2�4T2fD��h����	�5��[�w� �����C�6�*��j?����
��brCi�>W�䉿J�:��{4K�]��n{���%��`l�~�0�.[hw�����o��e>�+�KX�����X�]�喝�5�C9�$�'�f�]�G��ę���9����o/��+9��/v�c �XX*x��RSʝ� �Y�N%x:�d�%$t�fʡ�i]q�üWh{���,fB�]>C�p�� `��Ce4��ki�2X�̎f��Ma�o�f'��T��m���z"E��c%�Xe��Qf��wJ�8���\�
I���p(O1c�ĨD�0������Q��B�8ϑ�7Id�m���gg�#hݠz̷By*,/N��T+��-O?�3Y�>"�?��pi�Y���,҈��Ti%J]0������� @���F�����jy
���q�����$�v|���<��ڮ3'���;>{_��	s���kB�&	�Y�V�̬fT���Tn\t���f��K��C>��̧~��r�o��7j�_��-��	I����:�A.P���^[�>�7����#���<�ќ2t�*y����"d�3��g��7�)�BJ�Ds >z������G��o5�d�ftf��Z(C8�}e."��:p����X����:܁���u�G���4���,��� e�SQ,�Q.Zl���/��V���n����0��%#�����M������pr�BT�����!�2���A%M�;ٷ~㯏�Y�oe���-*�{��$�|iD00�[@@W�J��������2ʝ9�RƝ�?�-�������r��s��:`v��3'3�	��r.��ȃFU�4 d.���H��L�+���8�3��ɝBn���|��T���Ϩfk�)����=B=C��1rt �:fǒm���1}$��O�?$�"z��W���
�#���Y�tk?`�/�>��W�j�B���	U��p7��1e�kD��i劌�?�~�,t�.{������VOZ$ �=��y�C���h1֗$g:�x�ckN\.,��b�/�V���3)�����e�[2(�@�8��6�:s�,��-;q�x-��ѧ�+J��� ]�OM�6&�ө@���FL�.�ى�ZGU4�8Zn5��Ld��^���	�]����k�g��C�%��&\�&�7�E�K��M�4Dw�ҳ�������"陯���k[��9�RI�ho�o�4��a*�W�����;����&4�/�!��{�V#�o��,�g��w�j,��r:OK�;�ځ�.(�7�7`�yN���O)�l�;�5>��jL��I��D����èd�Uh>W�OB���d�ѧ�n���89J��SHGħ��i�2�t�X�o'�u�+Yz���B#�0��m����/��ɹ�i�W	7kOF��p�,��<�����ѧ�V�2��6{��B�[�S�&>*3�V��P��Hb�*K���7Jq��F;�ʄ$~��s���?���3w6|�r��!+�T�I�� /N�R���qcS.j����:3�x^	��e��<A����:�_�3��jO%���l��Q%�p�� I;�;��d^јx����@�ggF�-E5d uXH�N�����$���0O��?/%���]9���`�`�S�����*�#�tz3#.�t�-��[���VU�G������e@��G��@��]�#�K�Q뒆��	dG;�`�X��O���Y7Zk}����yad�q~[q0A��f�3E��d-�*�V��0܆ٔs���J/�f�(��Ԧ�>����BL�e���L������&���F���2�r�U�[բю�qX�>uD�1���-�}���9�Ӱ�͍�}��A n��'W��TS{t���Ə�4|��]\�)d�|.!��V����/���	�^�N�^[�y]�0D��Z��U�b�U�Ɉ�Fx���G�?�G'k*�����չ	��@����Ux���1vp���aYg����wLI�֭m�f�V���O�(��{�F�������:\(;�zh�*&Y{�^R�p�8��?d
�%;����4�?�$�R�'�B�_�v�}��h6�[_B(�p�B�|�AU�e�_����
w(r\�@\~�"���y�sӅhJ����Ty�%�X!<�k�6�(T[h�N�Y,k�j@J>/ga��;�&�׮�HDY�j� hg&P�#��F�'
AwN*S���wT��;�|�\�v\0$�Í9ٔ�"c�߽U���{�;`��f��2�~�3Ȕ\nʵ(�ŖV8��[��Wi�Xo|������p\����d�B?�
+��U�y�ܦ���:i!&+}�9u�yp�M_~,@S��q�69 �ڴS�H��L����I$��_eQn��*W��4N& �>��{c3��DG�y9���j�oa���6!�\���i7�c�c�Ҏ.l�墬+c�%��%l��N�V�����X�|?�}�®Z���j$2r�;j��"(�!�ޯ�_�;y��au���'�+r�G>���8ꅮ�5Wi���[$��9y�rzW?�䧴 �h����"f��?8��k� ;;9%�//�y�%Y���*�XP�14k�y6�%X��1_���S��H�ͮ���j6��v�O���3'd�sV
C�,2k��K��R󸠥coho�2�SS�x�|�t ~���� 9b�����0�>�1�7�&o�&e#k�aq��\jg��
Ѵ��E�89���%�<�)OQs[�Չ�HB�K1�d�8����bJq�\z_N d�zD
b	x1-�}}I\�\b�gF��
и_�@�����g�������:7]�{&P�w�5�U�K5"� �R���&V}��.P��R�W60��t�І�����6Tn�����W�P�)r�v>���J��"�7Y��Çȝ4T��F�iY�vS���y�5�l�&P0C�4�˞�:�����w�Ų^��Y�8L'��b�`�����%�I9��L�N�p�^B/ie�İ�*�XT�c N�y��AU���(y~)3>��+��a���4\/W�ȷ�Qׄ�W����U����I���l��E�\�t`��{�L�wql#jª�.��Ĺ.�4.
d�8~�%詡 N�ύ�iS��\N,�K���÷k�l 7�/��N{�i@ĵ����ރ�,�}VT,�V�Ҋ��#Q��u��k��rAM��@�s�ZR��B�!�m`b�k`�ir�Î<'Zx:�{w�z�������M����A)�X�}i��izi�����Ǩ����:�1���ǘ(:Ʃ��1G���rP��d���^wJ�Pp�L�B|-4�W��������8�J���9�>�67���U�`���tl�ȴ#�Mm�HH�x0�'�
E(�wj	e46s1�+aL�����ď���E�a?3h�CK6��`��ח���[j�����9�3����d_C�m��<�	��j�.ۜwC��# ��l�Ɓ�r�:�"|�ɫ�7g�P��c�F�֊f�R��\� H<՛�B�g���Y�.�G�j]m��:��Ԛ-��ܙw����u�l��Wn�Ї�@|`���,���G�}���Q�	vbه����I�J�Cc_/�s8�-�eR�	/m� ��H�����~�@��%�Jc�s^�/��(�gG�;�_cm�����s3�!����]u�Bæm^�{a�E��1�ݓ�G������;�/�%�͛�'>��i�t��(�+k�2��p�*����_� U�5�p7�~쇥er;��cUnBPW�4Y�=CE]SE��a��a�N��o�*J�#Ȱ�J҃[q�>d��Ϟ4�{"��at��/����J��&�_�>�{�Py(���d%T�*<���c��<V5�KW�3� d�v�rr�.3��P�(���Ԗ����n��_#�(i�V�V%�[���E"��H3y��	%W�@{	UK�tIͥCt�G�.M���/({=�z���[D�
8뚬��jh���1��`7 ��0��n:Q��v��t%3ı*�����o(�0�z�n,����|֗3=^�?���&=6���3��x���!�N*0�͘�ʰ�c?����\�}��,���i�o"��Cސ�=�dc�Խ�j\��]g��ұ��j��|i�9�?����f�ud����0��9��h�s��y"#%��=����ġ�@n��qWd�{#���&�ynlQ+���u�2&-ȍ4�j��bӺ� �/i{�X j�l���ɥ�gA�C�e�_F;l0�Bij{K��e��f��I��&�# 	Vz���Hu�Q�$���+�7#e���_�=o�?A�L}�!KaL^��lifＧa��~�%���{�U�3�p<����3�DӮt����I �L�Ta68W�h�?#�IԒ�u���j�c��u�EH�B����[d����6��U���x.xl��d�G��]l�S'Z�wt�([t^��ho[��$o�.���vh�^����� ������'':5��RN	�F���-�`������m��u�|�����f ���3�Һ�-�W��}_����F���/�V��7<���f�r��Y;�e�� t�qQ�)$�{�Й�N�$G�'���n���*���|���#9�MA^��S�|'�(�Ɓ�|;"f:t�VgAo<UOhX�h�L��X�O�E���C�vo�� V��zL�2��?]��'q=��H��dF�j��h�=A#(�,\p\w�hF�N����W���|�i�ߥQ�h9H]9m���>V���X��]pZ�\珍�z3@��c���,�h��In
�y�'��z)&�A�Q�É���Ck�Bm����1ϋ�l���.6����u{L�8�Ay�\L;���8�Q����7�� �Y÷c㗪����Op��A*��A�3v۾�G��.�q���J�����cOԏO�k�ve�s|���.,\�fw�eEp��#?��t�G0��	s��[)�,�sƜV������mOy���u�I3���5:;p�a�s9 �@��r�;M�B9�P��q��F���� O����X-j[�2 ���'ٖ4}�}z�K�+�G�B|��ǓM�3~�;{�L�z���Kv���R���d�!ٿC�� X�ə�D~QM�h�G!J���'���#�4�2���_
l�?Ȯ� ����\fVfL|����I	�����L~�e��Ʒ��l�2���G�%~xO�m��:�=�;F��b+���g0+Z�����[j����1�a/�3�A�}���g�P݉u�����
҆�=�8�W�5`N�3�~�����5��7�hPsu���r˭~�d�F��Q����o��ad��+"~�w�;J��=@���j
5XH9��Mg?B��|���6��M7��qHS�!BF+K?���ݠ�뤞��M5��ɓa��^i���ڧ1~:&�ː�?�i��	�Ү̚0-c��bD6��pC�������n�^�پ�F��Y���Ml~f�Hc�2��f3%��k�w�v�+��n.�����u�zn\�0��T�{c�����M]s�Eb/n���H=5�Vl�����5FHnA�4��Xti�Z�p� ���8E����"��b���{a�4͐�n�<�A	*H�r�ɨ5�z�AH�1UZ� ���~�%>������~uFt�0Z��!���c��qRR*]q��9�3w�fWʮ����b(�'�xj�&m�TM��	�p�C�L[#~�fp�Z��-�S�ڙ���a�o+yF���R@��?{���U-s2����F�O���R�
�ς	���=
LN��*v�'x,|
.��Frݼ��Z8,��^�H��������0e˝)	d�6Tq�[��Qa v��tȬ�yT�� ��aH�iZ�2�f�.]~�e�4z-��:��e��魸VŇ6}Dzo�}n�P޻=�l���Q���FM�3V:�)�qn���/���^|S���7��¨�-���f 폠���q����?�7h'�s��0�N�1�x+Q���Sx5��ݬ���{��+D��.5l�v��`��l�2$��7��!$'T��ܚԃ�o<j��K�\KN��G�E��Cy��������W�t�i�J�g7�d����� �I�\��
�O��T(,���ةR1��$s�S�F���u�R7�d��}~�i��e�aީ�ڜP;��+24>{��~�;땦��8NT�t���? ј�}-* [��Xٿ�>�
���'��9�0���+�Q�?9���VV��#!����V�S��R���NИ���ԉ�!�ޫ��#��}AYH�=��N�B��	�2�� 50{�gK�{�Gp��~�z�$<K�U��I@�j��铥��By���`а���R�"��62��.�������)���d,s2�0��k"��=���ɖ��(w���������d�<z���9m���ۤ��2Ԃ'�HG�-28�Wm:��~D���~���,��xZS�y�%��,��w�_rӓ�_�s�IdAW�J�n��tR*�Q&��(ԝ�]�+���W�p��'�k$���g�7s�hwP]�R��\��o/�8���b>C����gv�g��>�P��ypw���j���G���Z�c#B1ؽ�(Iׄ�s�Z��D֏���=�[�UE�yxOD�&Y�B���1nP��qǨ"�8Q}��Do��W跕k~D�!!A ��v�����`F�qU�#�D4��N�@[�vB��Ao�&�$��(xM�T���A������ǧ�&ۙr�7��$��q���f����V�
�~��N��T�;+�ǖ���f������y�Sn�T�eF|-o�p͂+	rC�����r�������M�`�۵M�I�L3b_$���Q�_��+��U�ׂ.� ��g��w�`�Ĥ�ۄ��+}?�@��Ӕ�uWqT��D1�	����4~Ѐ8��y(,��3�Fo��3�Oì���?W�iS���{rٳ�/�Z��i=�-o�.$]� r�2��^F�ȴ:�\f�J��2q>�d���Nj2�7q2F��[80V���/7X��N���!�>-�{���)��d�S��Y�,9�'ҥ��f��A�N��
G�Hώ<�|;�p��z��+S�i�����v��o��2f4E�r���" �ĦS��6�]��?A����?hQ��Mu7���B0������[q��:��� 4P˪���av�q��&��w�	���Ǐ��`�s%g�˖D���Wx��'�@��z�ڶ�n���6����d&j���!�����K<� ^HQԒX��Щ݉�ٶ��d�e�OHEFv����9��l��}pKZA+�7(uƽ�����׭,�Tɩ�g?�'�����]�d4mm��F)+�gA1s�̪��f�q?hO�S=����Ow-�+�=[* �iC,r��� �����.�c�%�K�S�ȴ��m��#���5�7#�.����:�����x@�� 6���t3�ꯥ8a��F�XC"lܑ{_��ƠA_�l:��i�U�Y�m�KMc����K��1���ɰ�dokf���Ԉ�wg+4�u�>1@���>k��?����秗715���31�{O��yj<�HO�5�@�~�ʩ ����i�����t�J���LJ��r�b�z�1G~�^t?�����%5�q���.-3b"XX�}j\�$ʾ��,��{���{���q�򝈗�
���O���0H?v`l8[���"��n��2�5ù��6:�^�
	d�c��=5 �\k25فB6F1*�քًAYj9��I�������B>�"1\����9�(�xL��Ji��U�O�n ���sd�H�%B ��x|�����l�T�Kf��Y��VF�*�w���C<]���0�ڃ�Lm�RՐ�������p}�HpG��2�.���G�Z-ǱDws3"/�K�7Fzb]�X��R7��F2+/��L���F���e+�@9 �Ѝ��Ǉt����R���o��%�ٝ���l�����z__�$��
ǡIآd��Cx����5Z�?��H�����cP��cU)O���Lg{n@f�!��I࠙���g�w�uO�� �ͯ�]J���g��1�br�*!�g=�]�8	����vE3	H��<�!����3Ⱥ��Qs�3@�`ӱ Rq�:w�\��"��(��	��Ձ�-2��0�S���;�])������6�������)/�)X�˨� *��2s�T1�@VH�2�U$��������pQ����$?zF�I�Z�Ƥ'�z��0��I���"٘��F}ĕ6�sJJݠ��3K?qlQ�ꮓh܅�����K����d"�s�2_�v�M�r�m� -�+�;��V8?ZN.\c�)ܰ���+QE�Y�)gF��3{�B����QIX�c5���t��NHߩƺ����rm5�n���������4D�Rz�?��^��8�ݗ �
D���Jj�1������ i.����gMĔ�e�B�o�d ��>B�Ik�{ή[�Q� ӥ�ӎ��<�������y��ۖ8�K�$\�u�5�h�9_��,�)1�\�7�1dt���f��+���3bJG�!D��=�O},�x���e=M�{�\�aK�Z3
H��-��Bꅁ�0��˖i��m#\_����gc﹠��թ�#��%���W�.:H��II*x"kP�i�)�Y�T�1b,F��ohP��?U`v:AR�h�p?T
�\�3�$`���I���8}T�yE�-�q��[�E��r`�b�&�w���Z����^�D�t}|��#���l�cXh�6"��{T�����a_�e-��B���#Jq�M���A�ǅ�v�)v��,��;����H�h���<tCM���&S�4�8?��� ��=�S����C����U a��v�Y�DY��U�H�;�P;(��I{E����Yt�2�
\ �ҝ�[e��}�K(l�o�bڻ�EP|բ�U�Ƥ�Rײ.�g8��Z�	����E�򑽯'��
���S;M���5dS0*�TgS�!�m��U��p8_f����d^�9�*�eKW[ל9Qv��<Wh�f�.#u"?��zkW�lUR�CHƹ�e(�����<z��I�*:i���3�m��]�n�h+��t2�)�]z�L�/A���)�,�h�*��/���R��2C.0K}�^�uݿ#��w��n5w�Z\�����c,��B�7�����{Or!��@�r�i��qzh� ���i���Fe��J:K9�T$�=0�X� �-O�W3�/�(9zT�1������R뻐�~U�N86��)3�ޮ�1;��j�ϽOI��	�US��c���x�a��F�׷���:����@#��.0Cؘ
K��f��y]ۿC^�pӧ���h���Q�)dyW��ym5���̸ƱY?f�]T_um��Dh�{ƫ�a�ihk�'��R�-ϚU]�7��@�K�M�Q��K�or�ɝq�B9aGhЀ5iFW��&-zo�Lბ+O'���+!�lK�n �e�:*��G/�U;�4�ܔ�����Z°(��̡j�g��#oʌΠ��;ؓf���^�][��� C�x�giN��?1(�G�W<�	M͠�s�a�Vn�a.��Ţ̚{?�z>i��W����BV'�vbW�,}.��m��ӄ�	�y9dz�%�-cW���]���/}�;�SڴC���B�[���TJ���r�+�{�J�W,�JՁ�q�'�K�X\�{��xO���gTo��3P;f�S�=I��ۚ5@��f8V��,�#m�="��Ԓ�W-x�;�I��ak�3����9N���r����>��l�$����<4;Cg���6��vt��^�J☔�
[GY������)�:DMB0 �0Pp�\A4ї�O��@
�86�Js������T�7^܂�����xr�-�� �J������7m���uu���m�����A?�3�1�f�ٮ���z���ө� ^-�U�I����C�0�
.���zB��&��4FiRv�O��'K�S�_��Jz��I3���}����k�c��cIĸ�
���F9Z�>(� �h����_t���b�8�L�����o<8�U�m�Jސ��^q�v�p�>ՠG�X�_�mi5��H7��4�3��v�g��A�7<��Ε�l�(��>�l���wea�l|'(F �P׹��S?��q���Q�l��#�P�ǔ�LvwY^i��5�LMI�-���I���Ϡ�g��<eA��&Դqb������>����{jifE̖�'��/�qa���qJq�F��[`\�n|-u��./r�@��v�� յ�� �;y�4~0�����F���|Ir��?��'j�5��}�N���lz'��b�n
���
�;O�l�h�ˇ�ߧ��2A�Y$��9U���*0'=B��"���ɚX��mZtբUg��QM�9�l�8�1���ΝL��6���h���z̐��R��x�+���qC��ğMm�ðt�9�?�B ���8)\�<	���~��JF�Q¡�<�ΦccSt��1rz���#Ka�9��9�9?������p���toSCuA/��G6����R6�&��r,9l�1Ƌc[�X=G�V4)ړi2�ꁩ%j+5�g"���2O/�i�V�>�
�P���u�iO�j����^эb���4��#
��[�����e�|�<�gg���A�'$�U���`�� H�;��^9���)^�Hv.�D����#Î0����첼��f`����أ3O;į��u�hû:��Y��έ��8����%:q� ����rL�3�5��j4Ǒ���x����'SA�IQW�R�w�4�NT������ZЈ��L�k�n��|�<��5
���q�1QS����å��d��+�D8ǖ��1�P�1���"� 1�zܛ[���/�2��<�wE��5�������[�q��K�Q2(�6o}9E�")��^.fŮzՅF��J�������x� '��8�]��a����.�\�l@�$7����
�m�O�}[��0F!�
�[-R9���z��"5K1 ;�ݢ��	����b���V#Rھ#���⽄@���df��+��Tv��R�tE�M}s��2Iz'�^xZ+*^�~ĈRΩ�ht6�y7����6�0n��j5]}~��9�����{��Hˣo�N��&޶%&�T���y-���z{��K�"�d�H�f�`ݶ�K?�<�����s~�@�-���5��2�	�����$�T����#pڐ��r_��?A��.0j�;����zg�6M���/7�� �o�n"���:��/����͟��z��}7�BjK���i���Ɠ�+Q���Z�c����Ҫ�f�7AG&@єi�Y�3b`�?�3�١3�4�`[]�L{�$����Q�sW�L{�$��/�/��"���U��b��6���9OF���R��,k���z4ϟ��6A;/ L����1ݓh��Ӻ�����?���T�u?PX[��V`���i�EgkǹӮ��薎E���m�N���7�V��9��`B{�VSȵјJ�FZC��iЂ�<�o����X�	Ly;LK"1���Zu~���p����7�qO;�"|���u�^J8�P����!w/͞�ĝ�R�Y�Գ%"��[˴)>+�Z�tB����1����I#�����}����t",̎y����,���fr���n�_�����N�c�Њ��ӏ7]`W�#1蒵_�ȟ�A�P�X�-��ҧ܈/�'ޯZڏ�����4ޝ��š�
�����Kz��d�(rKFi6N-~��5h]��
�B��cH�����Z�,v�r�)iP�� �zNW��P�#�n=!�%`9�dF�3H���o���-/��a�_�!FE�E�qk�-����(] �(aBX�z�*|j���<�{�,a���:���0h,���i�)&V�d�	��6��+3X	1���E�E����F�A`:_v-X{�OZ-xe��cYok�,�O����+�.��G�h�p�ظi�JE�B�F�.���L������I%Ah��:Ȕ�U��^*��NA��N�<\0�\匳�\��(�QVk���~b��-j�\/���Z[��y����,m��GH�����GG&>�����I�d�PY�����>I��y\f=��*���X���5u�K��)�������s��������F'��ܵ^�D�33Cq}[�|���|��{sx� ���:�ufz����V�`���)!'������c�J�_d��X�>�8A��o�T�	�O���=�&����wgK�����{���}
��ӑDH���WKb�Nl�C� ���X�����~��X���ф��I�Wf346|�}^��}��/�!y�F�g�~�� �WA����$��ۢ���bCw��}�O	�!B�CA�� �>�Vɩ�^���V#�6F�X������/�W��R�i�pcj��Mk?����=��b�<�����;�:�6����<�F!���'��%�N�c"#�l��J�w�1/�U���iǌ1JW'w#R}��b=2��dl�Ae��"�8_�9V���g���ʫf���E�F�EnƂ��I��{rgS�-&��E�0�Ä ���՚0�I[��U}0z���	n��q|R�?�yZs�4�"�`���������x�(����B��6�n��<,ּΛ������ɉ��yR����4���҈']�ìf�9K�O�Y �F��w��{C��"B���Z���4^��d�$n~����'V ��w�:���V��k�+E�$ߏ��D�J��P\j��ҍ^�[w9~P�c?Tr�Vh1X�]�G0��-w"j�Cx1�B������u�xW
�0�QW�6�������D�����3��q 4�D�+���Q_�w@�'�ĳ�¨:RA��}�s�%��ȵ7r:^̼yMR*�2`j{4��Y7@3��������w��E-�yL�g��x3\!�7l�
�Z� aRj���,�s'w��>]�y\J(�x�������&y�����Ք��\�C�#G�,���w^XAߢZ݋κa	�v_u�2ӤRE_�@;t��Ϣ.u�U��[��8p-3],�Z�⫮�*j�=�\L��72���jVVK�l�c���*�I�ǯ�͗B��Wt`�~�=6��t�n�\>�M,R6�?�8�_3��0������8�K�E���DWrq�h��� ���8�7��R��z���F������/t�8I��B%����9�o�Y�(l�8�2���%�]L����`���_��Xy_�
�B��f���!iG���W��1��@�@|� 6��vGi��~��4 ��Ͼ��,�5��͞�pK�;�oG�jS�>y���Mre p�j�y;����9~�ɥ3;��?�K?�fȳ���&�q�b��~�
�fd�uVg�F�AT���?�2�P��S��:ّҥ���sb��չ3~��2�V���&g��2J0A�����f!'�#)X��Qs�ճ��Fҿ��?�<�>º�X��$���?Rh�(�QW  �~�r$G:����X�g�н�N��g�ӛS0/�Y���$ͷp]�w\>w��\I�BNYDd�w�[�-�=�9�8��T����<"S�3�3�*xXX��6�g%��o6_��+\;ãFJ�k��C���F@�%]k�}S���=�;=����`c�Th��5�O���?6��,�mKj�!�L6�_��ؤ����B��_�B��\"��>g���������,.��5�8�BJڶ�J�Ļ�����t��Ҏ(ʼS#��lR���ɓG����U1n}5�h�	�� -'���Y�!M������ �rw/��]�0�����Gi�U�V��0h.2/�]��*}���Q�xU�`i�~�&�8�����OJ�~���CE�U�h]��3�!��LYھ0�&���n���wBϜ���ڙ�Q�S�]�]�BT����N�C���؋�p/�:Z#:�S�~'����cl�0g�g5�V*�P���Iψ�\F�nԅ0+_��$�_q?�dO�D<�$�30�Z�����f6i��j@i�+7 ��p�t&9:;^/�T���qa���TIW盙�iw*����Bߛ���G0���#��> [!�Håv3gj�$�ew�	 z8f�X"�@��+��T�+i��\&�:?����O�$rj?$V�P�̈́��Y��P�_J�r���O�k����Q��Pݫ�T�BjY��F�G�۞|������ĸ�Ď!*�N0�K��	0�T�1��5�̫��g���DPj��ۯr\f���q֛���!q�P��rV�g~Ve��u7���u��~�~�fS���ƌFzWp[���d��p�����h{o���^꿆Ɗ8;m�p����ɮ��$�]yL�ق�$�����zl�\E!�;7ΓgEڝ����^�;����B¬kZ�&���d�ޜB|4�c�{�(��J���p��#<p9�k��Că�+w%�t�Phl5���[��\·i�5�k�9�_x�uC{1� ��?owb]�WS״qV1�ޛ���7��r�E3��Gv�\v1�t�+(���,�K���y�r����{ �SX����F�J�Ƣ)7��A����6<��6�F�4,p��H�l4dy��p3q[.�����sQubM��mJ����ʤ~�(�:��?�L�͢�d��iuM%)�%�<)���`�:1���#J�w-̤��/:��.ٴ�)��&
,x�4���tC�������{ ����m��m����Eo�,	����R��㸟Z�G����n�D�;�1J#st^ϭyxB�3"�
/��b`���U^ڷ����u�r������}A�oU^~�	�����t�(�	���i8�ݫa����Z�{Bu�=1��k���ˇ^�8Z����E �| x ��b��"[[(h�QG�b�%���0�eنo&��)�u/�m���T��=��f�yI�<�����w�឵�=��Y���f�4*�*�N^�4MuXZ���Y8�0�m��c�.h�.1����'�D������vI�־�	/@`����R�J:*�W�[�]x�y��0ǐ��{��KU�m�Ƥ�]`2�˺Oqu <:t�X����q7_��+���)�?�/����]Q�
�E�]�&�rXV�#�Uׇk5zRR^�pis�:+|hd|�3[{%$�����iP�2��m� �������K��O��5p-��߲�$��@U�F��d\�n���Pv
BhȊ�=��`+�F,iMal�� ����q�=C���}@��j��Ի�e�y?��>E�2�l�w�������^=F��N�k�1��
����9�ś����F��Y3��{d�����AKp������Bv�F�h͝N&�*U�쏇��O�u�Xשּׂd繩�5Q�"��CIqj�T=
-{~p��1��ǀ����^�X*�xșk�9�,m���;�"��3}4��#�d�[ �����d�J���p�~:��x�Ζ㒒`��R?�x�'�����(B'��L=y���8cW��h퇹R
&�B���+��G�́��ГxF��?��f��&�jL"�KD�_L%k��M�������3��8��v��b�;/d� �x2��ן*��h`z�;;+�mD!�ܻ�Wr��z�)�̀�`��:�];����)�0�1�鲁~�SZ�W�%o� c�_����nVP�7�4)��T.��W��f�X��v-/9s���㮨�7W"�r)��T�t�J�o��O�y�ri�ĕ��S��䘱W�.}��G�%M�K�&l�lBt̗�r�m`�Rlk��6 �>�f�J.���ٶe���,�ǝ�k�������ե''�EA�	5�R�;��ʮ:(J����@�䥫?5���A�AB�9�}-���I�����H�#yt�����9O�;vA��_%�	E�I�p$
���s��C��v!w�]ʴ�0RTC�ߩ�1�_�B��uYـ7�tHs|ʭ�ԏF��H���I{ ���P�G�e�n\��l������F�4J���I��p���^1-�P���`�^�j�n��wz֟�
��ar��u�}�9;?׷j�7
�v�xg�6z^��U��@#H
���\Xp;�/�|�"AY�T�A��.�}R�OZ;�����O����L���`���6�{��߶Q�-��@r(cC�W�̙G��oTGp��L7�oj�Ы,��?�d9T�>e�<�N��Ni�'lQ����U��>��E���g
���"�
��b��gY��ؿ�*��́�	��2`&��{7�.G9�a�»j�_��&U���R������bz���;��{%�\]鉰�jN�Yd�&w�
�g���-^1��=p�� |ܩ�����P�ƠX;���V�i����7�^�)YTZ4Ze�>-Jw+YiT��Ӹ)��kTGm_w�۹Nt���0��_��d��z�q���p���Ap��*�HT{!= *���ׅG���,���A�8g��@mK*�{q �q�Kxg8�]�bxRt�v��-�Z�Ӏ�R�쩧)���t8�c�қ�O���NS�Lc����=�4j@O:�T�;1��~<�����X�h�~oX;D����d�n��{*5�����������/��FT$u[ {�������#ʉ�Br@K#G91s.C9@CX������B&����Nd�=g�X����T�oaȎd�\l�op�ބKS�C��6^��{��B�]����?�6@��7*C��\r���=���X�['Ϩ���GTz>�p!R�L�@)�����&�.���M?�x�o��n;�۸�����x�=�-�&���}V�
yq�o-���9E��Z��ے��xo+,��e��[���l	ўF���K!��0[���s8�O����N\�at[�x�4Yt Z�&����'���
�aJqR�x���|�-"���F_;7�����ty��o!^���$�Gyy�N=ڔ���),�L�	�SB��TU+���Xq ȕ���ޏUg�������������R�zK`��S�/�� [��ZK�D��	����W��d'>�خ�\�7;ܩa�K���T���V���D�Q��q����:Ѓ��G�,�uC����R� �x�͙�cZ?y;�@"%�i{@�U���-߿"��>�)�p���p��1/L�^�4R�~�"�6�t�&$4x����9�Malwb�mmq�]��bli����1�Y���2��Ϗ���ԉ_K�
��k%��p�]c�r�2]��0H������0� �
����A뽀�I0�[��쏦��:k,�����ے�C:(�}ف;��T���34�[�#������N &;�6iϮY��.�^px�
�� ��T"&�?�E_Ũp���[��,�qO��i���]ĵ�Q�ʍ.�&��fٚ���Ba�_ߑ^-��D/s]�`ͅەZy
��ȝAΩ�פ�U�,�,�+���{|=r@�?��z�
Z@�0�1�THv�گ���FߛU\����8?~U;���ǈ� �,;�(�1[��j��%[x������b�*��9��E��HA���}W���Vy! G=�4G�(2w$rVL[R�� %��iҵ3�W�>�D��R�Y��\�P��頻��qr���2��J�"]��4�B�Z�k��?���v��I}p�q+gNǚ���v�)���l����0n]$�aF8�`����������hx,����mj����'�9�����k�2�_�"��ς>��i,8(�|2�M�&�]��O�������I����*"�*���x	93쯏1���rH]�M�nξ]�̀ǘ�n�A��eЋ�14���xo��ɛ_��s�D����o����8mNARl�(�6޾\����I��M�aQ�d�[Q�t��I�DE��x� pLn0^�,�e�Be��;���|/Z1�� �3i�C���ӿM8����G�M+�J6���ې�����P�r�5I�ʥ�#b�#����9J�SF�;aI����Oh]5]x��Sߡ{+����`���^���-C�	7(6����[��5Yz��$�nc�
~���.� "x�"�.&��u���,���-����R@�b�6^��o���m�H40V(O�ߓ��+�_s����_C	�aI���dُ>�6w�v������mP�;��&]�R�5^ث�H:���al���2]��ћ髐���������xj3�$�«L�<��k�&����-�TA��N�t�K��B��!
4O��n��_zui�yN1��2�_$�>ˢ��9�)�
���HF O�v�i�`� #<��R�y~�y��0wF٢���r&���Tb�r�4yx��`�U��[�����g`P���˺��[��w���	�YpZF7Ȏ�Rҭqx2F����f��3P"�����h��\���|�j��N��N�
<���r%U���"H~�٩i:؜��� �F�sZMd#�n�l��2CHmS$���=�p&9�dB�*�Q*'ي�L�y�1�@G����X����O��9�A��U����E���C��I��e�l9�v�$�Rw�[��e�ʨp84t:҉>ZG�b	J07��g����w~��:w�R��@��d�+x��L�
$�L̠	��;�ř��bA�Ax����~��Ӫ��=yOy���5�r!���ٽ�jK����D�Ј�0��l��nY�Sv���;qs ��ݶ�`�gNm:����Є�ET��I��z���ö��Pd��3[L# 7�g���-�J�����ގg44��<��> #+�Q��q`�pI���u�%φ�iW�89{��<�Ok�����]���&X*�c�Yo� R���Ǖ��y����B���G6�ˈ$���?���ɘV�U��f�| 7��~���|�=
����F�ۋd*�P��p�P�>��u�D��k^��f.@xQ�o�^�ZI�K�J%=B�hiO��:�Nb#�O���ϣ|����"��K�[���+0�2G�8�Ux�&!O�c]!^�[D��) �L�qe٥|r
�N]Lt�R���y� ͓�W�iv�w���;0}��X^�[]�>ʋ���wF᠉���dV�Ts7�Z�&����{ֳ"��O���f��fN��هu�m`l�6j/�1/ ��WE��oe(��90�����t#�̤�R�1V�t���?��E��[����]���=*��`�$D����]�>�н'���@�R�.5*u<&�m�����)�-��cE3ӓ<��O �^�0��6c����Q,�/�>�6�3<֙�
]GTѬ�i����uNZ�,��h� �{Q�.S�I�%�O�GSP8�,�G���x'���/�/L�S2:����9���j>�C�q[�{�n�0	�3�9_4n��,�?Lc T&O��!������*W1��K��
���b�\���6���*��B��u����ת�V7D�K�ɫd!�'*'f�z�3y^@HsRM1~>"���IcO�e�K�`���OJ�[0����4��k��jTUԭ��W���8��6L�T*1�F��}$�k���<�NpU� Y�w��e�!F��/�(�ϋ�0&�5����O�ì�R�@"u<��vHy#Yf��F<�rE��{�9�ۓ��yt���)v�.�������&�>>���[��v���#�˼ߩ9�C����?4��f\����uX�(z�8MEK��JWRr֦@���']���Q	g�J��K�S���!��\E!��I�����G�5�iV�p�S�Ŏ6ɇ�O\a���~�B;{����? '8������Y��y���ݢK���{��̛Ѹ��aC�=K���$�gm(�ݑ2獐%r(���wj@`a�#�Wfet���`��j�>9���EY[����מ���^S�>|�������������(u ;ɥ��!���5�]gO��w1J	�q��΂3x�������`���
�G�Y\MA`�.�D"5(�Hy-	C�bނU��v&�+խ�.~b�4�gMʶ�VԞ	BE��yiB DAْ#=����=�0���W�����9���_�uf e,�P��X���44\��	��︫VD�$t�J������>Ee���`+�n!�1)�BZB�I~�Rh �1 �	g=: M���U�
,ڨ(�!�W�5��[��*�x�*L�oܮB�5����N&�L��淞���Õu��=��xP���5_�J�a��0JVV���T	bY�q�;I�D�����[��j���7jH�%����siӀ&�Lmw,`?ca�\$�D��9/x�;����m��~�\ ?d'�Y�z`���6���V0�?P,L �@��D^6����f�&���~Y�B�KG�����������������t�����-����K]�q�듺ꑌ����9�F؟0,���`,?�r��s�������T�ڽ�*�t|�WE C����`ӗ�h�s�Pjpm�ؑ�J��ؔ&�c���r�b�MYI.AH���f8	z]C����H�Ǣ��4c�Ś$t�0[c��~c�t
��O��V�n����Ї�ʱ�{D����6�4����U6��&��Ȇ�Ө��ϝzH�2��틀4:j�d�5�����ul��ݧP^*PH�'��E��]�*��H�q��ˤ��+>�,	��i�(gP��u�< ����2�;�DZ۷	w�{�JO��
&��H��xd��Z�#����x�d;l[r ���NQOS�İ�g���&v��N��Pf�;	x,2�[��^���i?�^�A��)����$�>%��;���}t�%J|.|���("�S�`���վ� �!|��C�B�m���M��Fm�}S!���^?-�ܗ�Z��9�lC��>��@}�W�w���)�Ȑ�"P�|S�M���m�{���t��cRg�S��ch�bI+��#�Z�Ⳬ�>�ʟ(*��"Kx�Y��Oz9����Y���o��eJ�H�)�,=�JL�C`�(d���&{��dXb�u�FQE�����6"/�46�A�F|����h�ǽ#֦'��Y���z5�^(�9RĮ	y|�-LADb��#�N�<��S@I��'և
+ڇ�i�N3q1�0`wi���]��D�n���d�;�U�=�l�ΰ�Zm�O��7��^Q�����}�)h"�z����m��2�GV�p�RQ��9�h����ߕi�ukj<-���I�O��;�@�t��ͨf�[s2-��
�d�4ճ�獱�TZ|���]#}�XJ�f[}P��s	Õ���%��Dh;6نjݚ�{�K����w��ԫ�����\^ )���j-�|�:�.|R~-�a�w��jw!XQ�-e�Ӹ�}3L!����� ʝ[ �nN��rD
���	�h!���Z"���[;8�i�~Ar^h�U! ��t)wYߪ,�9�<$�������H��1�fz��v-.�M>� ���㳯m�^� ���8F2ȅ��K��������U��t�����e�]��V���+�J�v���������Xy!.-uˊ�!��V1�8�2�Va+� �V���0O��PA����7�ˈ��ؘ;����:g��gk���e'�Ƕ�]�X���8��S�?{�s�SyãL7�k�T$oE ���6l�q<��R�8��Jc�nuUQI(i�� �ѓ�&=ۄ��8�8�ԙ�V?	82҃��`@j�i%�M���{sA�%�E����GXR��[g�a0'mc+����š�|�uT���|%'s�Y4�Q$����Afj7��d�V���n��Mw�y����*|��x��Fxxn'K��g�y�*��Eq.�T���Hǰ5�����{ŕ�l�RZb+!��b�!rl=�p�	�������	}�󌏄���Ue�m%FAņ�W���N�} [�d0�P3</O�b�X���6��3�^3�A
���/o�+,q����������j#5��l�;�X=KX+�W���ޮ����]�^^$���_��;���M���ി��9��UX�0�^�z�-9c<�%ߙ�4����~W�c8}A��Q^�#�9�I
Dx4$��]9�4gX��k�K�lp&\{h�g�øfӺ �����J�q�Ќ� ��\�v�����K��ķ�Sp�Kd��2�>�Y�bg5�Ur��fHG8���6����/|ljWp=�Çb�<ez�W=�����ғ"�Z|��&��j������K�|ʐ/�]��tH�F��� 鯪\Č����>��߰I+#g>-d�6gLO2"�K6~�$6��ˈ��Ժ�~���?	H��?p��<r�B��k���'�T����f��f{o�ރ�G������l^�m�2/ϳ5��ו����-f�{'����[ ����H#���T.���!���E<��߳q�W�wh�0Ȳ㴠u�Z�ȇ�5/̊�;��LI�BZmv��eoj�Gɰ�e[�wѺ� ���(Ճ,
���K��^r�V��k�X�FB�
I����᳣�QXQ��r:	�K�4#�w��Wڙ�Gb䚔��~�n'p�N\�L�>�^_�7��vRK����6#n�'��1���6�(g��]�L��g-(�0���\�+4������k�JT<��A�v+hm[�,�!�h�����wi*h_u�0~��N�cyo�E����T�Wg�wʣ��2�-(ڇD娕�t�ڶam�̹�R��t��㱣v���>�J+OB�<�֢X2��{,�&��ÚfQ5�Q���*��{��6���(�R��[]G7��NHe���_W*�+o~��	4\+;�NE$�[Ք�KVT-QF��>�z8���' (��h�w	��?]X@���f߲�1x2�@��ɂ���$6J��b%Ķ�ޤ��d�m{HA^�nl��<OrX����Ǳ�[��JA3hZ� �����}P���uT���ir�5���u���mRߩ�3�`���53*DdlF�cuD��N�R���ez�O�C|h�6Z s@������};���=l��ˉ�#��O7�Nz�q������_��L2�%#��C�?f������(ʙ�1�0PY>�J�-�ۅ����$�췒��A�z��<���=�4640�P�.��j+g�t\2v�T��CS��*qY���~ܠ�aǆb0[�Cr�]fI����z��V�ъ�+Z��3$e��%>���t6u\�e��&+�4��M70R������,��?��#X���jZ
y}0|���q���Z�@��&�̦��e���P
��@7Q�W5��I��m����i�+��q�i�:�l9���]�z���S4[�TS5]DK?�e���D�~V��h� ��}8]��X�B��i&8d��l�����������W׫$��i�mUyMC!��=���S�0u��G�x�==��]8}�Ӕ���#�c���$��Q�w����������yVS ��o��6֡��<�P4ڲ��D��)-+�r@�H!%���mэ��k��ܮz�j�d��g��C@NyH� �s�῁lF�f�OSqZ~&>�4h�t�$/q>�/�V�o�t�kW��J�ص���=o�p�~�M�J��o�)b��ƭ��G���P�5�����r|�@��M��m�g,�ٚED�$�J��*>ϼ'�Z2���5H��bk��Iɲ6�1S�ՙ���´pܫ��U�Ar��&��7`Ri}�˃�ү{�>�nx��Ζ���1t=/�NC3�NT�^����X���'t �̧4 �]}����x�o��t����dm�~�^�B?���ׅ/�@��6c$N��F�4�d5S
����� �>۶Ӕ��Թ� �����56$����I\`�xf�^ѐ~�(��4� �Ii����!��&­�����m�{�����x�"��Mq"C�d�"��h_1Q%�XR��)�'_��A�����0�@8�	rW����^�P��P�i/|�}��f�I�l�t�Q�#t74��}4���]XDp�b}��[0�*�P��Z�Έ ).T�,%w;7���"�"#{�׵pMF����ZXV�YE�vO���b�&UU0W�3�������� �cP%㾈�&����O@�{p�;ɫ��͗�;*|�� B��c�
G�R���[�O��d]��}��9��	HV�b�m3�����VN�R���o��joSДve���d���0�^�!��"i��B.�(��V��$6����	��c8j��&��	ؠԫB��.�%)w���Af�˝�R�~���<��¹g%�]"��"IX�kҰR$�
E��&F�1 ���/rA}�xrk��r/��G���2�`fr��u�Ͻ��� k�T������B�+iԑ�����6����w�U��'�58(x����I�9T�ϭ\��V5$�'Y�c}'��%Sy��0m�r��T)yc�ٷ�����W��F��t���۫�u"�:��_�ˮ�h��8h��T���V���l��O���҈���Z-�f�0�JeB�2VL�G�Z@�f�?QAr�RY�I�7TNm�T��0q���Y*���z�΂F��*�m�ٷ6
�pr!��/�ڏ$����He���J"��5L���1�O�;9�a��
�_�-vn��2���_�h��@DQ�m�ۑq�ru��-����	(A8��U�
�����Ű�O[�9obv�o��t�I��Zψ)��zN��p�E�w���`t�l�=�� 
�xt�c�<i�@%�C�8X�o�jt�8i� �1�*�@�
��>�^���tž�{��m�DKG3�>���ʮN�,�2R��S����_W�8��Q���S&��J��.�!����$��U�mNd餆0��w�{g5�]�H���֦ܺ*�!�����Q�[O� �V1�oL�gW�j��(~
n7f�Q��U.�` �g���]��p�����O.m3Do��bb����]��7�9��v�e��O=�	R�h�?D��[~�ӛ�%"D��3�]y(,}|��HYN���Y�5�$̟���]?@>�<�4�6�<�Y4K����#��|�7�9�d�kz��<�L�Vs������� ٢P�S���A���z_x%kZA��G+�܈ٻF��«��uGl���j���1��c�0&�}�$t�zh$WK����t���g`U9�:8C�ɩ�LȅTA�Ulh4ocP��s[<���?��ux pJ5+��U�����mnV{�O��ٲ7��#�(��"Ü�	��E�ǳz�2��fInо{{k{Ijt�N���)7�����s�D���ը�! � ��u�.�.�����ss�@�V���:�/Ώ��n���e(ɈUT�5�SYrA��Y��v�����a����,���a�D!31���/��A텗��m�H��b����k��Dy��;5��fQ�<�t���_o��9T�D���`dW����1�LJ ��k��N�];4�q�j%�4�HǮ���0zc�ӎ<�h�����n5~�*��5&�F���Y�7ZǷj