��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T9 �0��\�0C���Ϥ���'ZYv�ґ��V<z?�xK���W�U����w��R�t�2���3|�1�ǆ��d�Ms/����g"��X��wT��G����d	v��d�g�B�Y0��g.����pP*7g���A��V�!�6��i68X��0-�^!�����{|�z!�S�w_�O��Q攘`��=���]x�j	�6�~���u^��J�7�;!m�<J���@	b������`�m&W�jNW!��p�\�.|uw
���%BP�H�5)�1#��QG��W�N4���r��M;�&�ʅp��"Sm5�]d�=���^�1.��-(�9�Jk�s�+gA���lwfH�ϸ'v!��*�& �ة�97��O÷*�"��u:�xU�) ��J)�����aPf�Ɇ$�zV軬X1����ƨ��
K -�i�?r'k��t����&���D�鬅_"�fV�5�}�M��ῤU��[�n[>��~��&��O>EL������I'B�B�fy@�bD��4������5%r^��Ur���|�:�)�����u'�$�80ZG��w�t�-o!��}��%�P�/���nG���9��:���6P�	 �䤫Hk�}}5�+��r)d�r�����z�mOs����W�C��&�^l�`���� s�3Ķ%zF�D�:02�׾�Z\�C����У��3��-{���Q�#DW=8R�Ѻ��M �{Jm�+-WՖ�A���B�E{�m§}P�m(�$����>�b�)!-�[TS���."��c,2[<�����bI?HC������[5bW����F����1$�+D�o�Y{�o�yrU�ɠPN0���\9ӹ�W�Y}��X;bv�b��чU����l�����+�!�H4v��祥X�S���Ѕ��y�~����=X�"�y�I�3���L�� ׊�D�h�0h��g��'Τ	!br�;���dM}���B`��7J��|T�m�5VY0C�P_�d�`Y�G�Vvs?���~ &� ��G�j��}M7��Q}��/@���h��\*.�Ұ�
�J�D�~V��4ii�jO�	��R��/e�y��;��Z�/�� ���i�3�e��������|ׂYU�S���<t�<E�fW4߃Zޘ=��X'�m&qf����yZ��πL#�{��C̫�
��h谥-�������R��ézHc��@�\�1yU(~5�]8����ܘ�j	�a���]�p��j�w����E=�`�����b�uR�rȎ�����H����]<+��&V��n8)V���v��ߧR?+EP��߳R����>}UN0�d�"?q��-+����1���F���p�����J�M���c�!�<�ecwt�]��&�Ψ`ٛ��	��NĆ�U�X�2�{@�m�9�,����ӥS�O��&�'�c\&|=�2��N�rz��L��7�Ր��Z��e3���}q6a�{���Qp�	9�cȢ�_O���D�r�\c8�L�D=]�x�:�V�6�X���=I�i��n��_.���0��V�Wp�ua���qUj��=}ֿC��?��`-X>����H����|=��X-�^�蛉�����8	���r��-7<���{X�CGEw�����4�i�����q��c6�#H�BR�"U� �\ ���f�Vr55kL��*U�ň	��3���0�u�B��Ј$��=.7�R�{`wI��w�J:���G�6��U7���|.����|Hqp҃�����=�
U�*/M�D�,o����l��q����P�{#�Zh2X�KK=�,�.���PU=}�0x2`Z���(�ׂ*�ڨ.���w�wƾ�O�(P����J ���:(��׭������=���������Y�����ER����ظ��:���ɇ�����Ӷ���~[�b��g�e|K��3�'B�E~&�������*��N�}��=�L'|�J0�Y�<S�e�ARe��p�I�lΐOuJ����'E�*<;3�g�(��-Ȣq��th�͢L��d�Nܐ�i=KU����V�J��	q2[�_h��]��ט����2n��u9$�U2��m�	%�8�tR
O�n5��'�A���j����vw�0Pj�'�U��?Ƞ0��4<��	B�9�p$���4�W�.k
j�5�&5<0R͇�Y��fQ����g�}��#ꓺ7��E�:�6ڕ�Ƴ����'��b�U�ٚ����.���Zѵ��z.�wH�d��SYg\L�}8�?��4��mn���n�O2�_����ϔ���s�g�U�fΏ�YC�tl�/Ro�|Ɇ�/���&F\�r�U��:�E%�(�b�U����-%P�u^��/:n�]��v��h4�^�f_�~�z&���"����I8��d�!�2�փ�O��-�n.~Jx����%'���.��Փ��1�%	�*?������7�Y3�����o�~y���`Y}6�RYV�p�,vQ(|�jT��)�t�!�$�݌���ӫ�JQ��#�V=,8ԗn7��/��?,*[lA<���K�,g�p��A�=婶pB�Cu����u�j�#�u�����ߗyNþ�y��<�
�j
;���K�p��H���`��깨�1Qz�[K&���	p�Ym����vx�q3C���ڑۢ���</�f�*�<�b��KJ�(�U��JКN%��/�=�GF2t֤��]n#�ܚ,'�����T�{�;��rR�ɉ�c�z����}��6$<��?��7]q ��*݉�8�eaxfS�6b}>�K/��hiT�ڜ���Ҟj�Y�����Cih=q�����ɫK:� ^��1�=+K0��Y#l^Ҝ2�r-؛�����!�t�w/�j�u���!� $E魐�J%(��p�Fa/Uy�yp����Jw�F��,����x�c�	H�c�ofdY]�#Z�J���XT�M\@�w<q�v��m���S[�X˽v4�8�G5���jWW��0e�W�)Cnս��I��ݙ�Itp`��rq�1r|���T�W�W�gUWr@�K�6$s% �)Uge�֧Sx�vV��/C�������s��;�l��:��	�iW�ecrW�G(y�;#��:��������A���J�{
���c�2�-~;ì����i�N��F��r\����A��D`�P[_� *�n w{}�� ���kCd�������_N��^#��N�`b�T�~�>��
݉6�� ��l$&OO�z֕��m��p��c~1_1�.-���~�%[��#!M>���Q�@(�y?���$L���c�W�>�=�
��`u�����ۘ2�y����1�خoLd���ĉ��Ǳ�T�|�덃����:�s�);鈴ml���]Z�e�uD��'^�Q;�9�{���>w/���{9jl%�.zMm֠J��-��{��n3�uB|rsZR���
�I%��D/�B[���rOx�`��w���4�F
o7D�F�`n)A�_��;7�\��a9Ŭi<���ų*կ����`�5TdNco�O���oD`�lՃ%~�e��}�?�y�y�?|,g�Q S�}WB�<6*%��j�Z�4
�p��2��$p3q�-�Ro�o�E��A�����VV����O=t�0�e0������2�%�X����(���f
�K#�a�n_����?gY�(�����<�`�r�K@�-aFI���s��6�<'����1�n�`�)���bӃ�ѥ�Q�l�x�T��Wq����s�j�e[�4�6� ���	F�̓�BP�><f����G���)������
0'����%�?��*���>5���6=�oO�YC��N!��N�
I�\�{����&IH4�L���Х�RK���G���owF�x�K!�y�qՔ@|���8ߌ#��ƅ��e9Γ5ʧ��|/�������'h����_w��{l�^��S��Xm"�l�����Mc�W��X꜁��/ы3%���v��j7'I6��fG\Q����l�n�m��a#�xt�������7�����ZBO�)��H^$a���e�^ib����� 0�����{'4c���v�͸���5�TlO=B&'�i�7�x�Z�K���}���b�}����hS��[�ۆ.�pW]ؼ�`R�]�M�v�����bo�q5ae�Bb&�L��y��Y�$��`��Q��c(����i�<^V�1C�#�����!�
��ѷg�9��=�^��"C`^��pGO� {-'*�H��(�(���f$�i%I��H�$��79�WG�qEg�`t���W�����>Rq�|�8
�Ͳp1:HϹ@jZ`&��+���UQ̮.Z�:-��.���kߋ6�}�㭴>eͨ��^`�v1V�p������6 �$@��Џ���Ȓ���q	���3�	+Η� L�'�ȇF�6jJ酫��>��O�G��jc89�����t)~�6��cJ/��Y��<���₡a��`b�l.r"�I7��LTtx�4���u:��<z�TU��K%�ڴ���U4��cx\>�-�j�?v�js%���y���{��mC��~�|T���t����c��0b������� �+}��0�G���&�lVR�Uc�<�f
����M�%DT|�Yt�cb�O���z�8��5�\H�bĆ%�;bkY��3�*9B��l~������\x��N���f�V�-))e����U��Ȉm�_�T��?e��^9�[�ؤ���J}a�ծ�V�	q�t����	y�wr�*:���h
�� u���k��V�ƾ5+�9\>����oX���O�ο�`bcTM�
�#7�N�@�x�X�'�!��Է�;,頎:V؅5�*ѕ{{�(W>d���G��r�\&���q�M.	��W ����{<2�=;7#��B�� ���ލ�{����w)�X��Y��|b���5X��y�yC泲��Ҋ�-O������d��U7b"�5�Q}[m���E�lr6n�4T͗�Bݸ����m���aY�t��L� �.�cV����!�*p�gs�j�v�9(	��_x��k���"��?�mh�_�����_��� e95�������D��*���t��{iJ%�Y3�/�MM���W���C�s�G�1L�����ͳ�YG��ʚ�8���Q���g��p�rl���wO��#4�D�,B��x͔�ϗm�����C��|jhr��ã�}��l�C`Q~&�G��:�R������x=��oZ�1�q��Fs�ΎT�{�I/�Ǘo!bj������xC��`-(j �-w#ekrѼ[����bO:�����w5�OUGk�����#������&���+y��8QI�& �|�~Y�2<Ĵ���������nxۖ^�j8���eJ��.:��-�ᬁM�{�Qa��D�h��(���΂G�rK�g�<!M�U�.�zW���_���'��'�f�J��ⅵG�Q�h���5ٮ�݆��m��㔨؄�'���}�K�U���$#�VSj��n�7�Sze�<,��"-�_���uA�-Β,E<v�,�샽8�~��қ�]�b@Q�g�dp��f��A��e�E�-�;�:^6�'�"8r����7�R&���O����B\v�=PJD�[����ӌ�<���1�m��� �w�fT�/�r*젽�J��!B�`���C"�/V񞯫�t��d�SG�- ��;�0��vM�H�3\kLK�����`&r��p�n��KA����z��Z$���:��|���%Sa�"sf��/f��AcѾ�U�+9ԢM/��J��Ľ�b�9%�H�1�=?b J�t��q�ЭTI�Nfː-DÍ#�2���b߸�Ĕ��J�-XB˂��t�T~%��Ɠ�%P�������r���Q%|�15G�Ƿ-�NMk֣y_�RM���7����|�}�Y�=	0C8�7�P\����1꺚x�ǂT�����
&��>�Ik��ͅ��R��c�f�q<� ��F�5ܤ��jbo�����CV��i8�C��u����C� �/&�R%ni#��VZv�J�(⇦�=Ȋ\�7��r�Z�@A��C
��m2D���3װ��1o�'��}�U7Q����{����6�=���1�"n4H�������X��������W�%�1�|���v��ڇ�P&՞���e����������!s�.�fE��s�����ƞs~���Au|͉/Z�F����(OL�r���&�\B$Ӯ��9�i�i���x�Xn�#�q�fxY�g�̔NO4��A��ժ[\ݴ�rT�8���V�m �]����Nѭ�h���x����Pp3C�'7b���ӭ��e����S�{�`��s�a��s��>�Z0���eS2���?����'z
Ø.3/[���c�c�v���q-|Y'=bP�]uT��m��NY���j��}x����mK&�`Ϝ�?8&D����=⾑蔎Z�?������rx\yhr�JP�@r)ܴ���K�i�=�ڨ��П��-6�z���e�%��#}Q�E.���8�W}`����|Ѳ���v�����42,�4K�:���iu7n�0��U�uؚOy˔�R�^���∢� Y�;zŲ��d�6���A�|�.��w�l�BW�p��'�~���?F��������J{��0����*�v�|��f�FC ��e2��z��z�H��Y����!U�����2����zt�����D$���5�?��y=���c�<Z	L�����Tæ]�;����>%�^�~�����Oۜ����-̺�dY|6�>���jy)�aJ�4�)����-l��+���T#4��$���R����p~��P6r&��|˓��0Q��P�T@�r�R�!�z�uL4 �P\���S�,D2��*�*�5�C9.�*>�l�I�r�n��}[�*i�,��$�*@��_@���2-Ñ�[ii�w5}t?g|�������'�b*<ˠt��0�7}�(&Et��o��Uz՗]���f�ԅY0\;�K�����������J�$�8 m��r���є�m��m�����+�=9��8�DgU�ıDR���aE�a�i��nұ:vpp�K
����W,ۍ��r�Z&�?ߤJ���K�m� ð~4_����u�_���
���8j9�9ЎH�u>��U��;���o1?�~�A�b6S��~�)�~S��s����G|�MYn�ޡݭ��4�d�o�+>F��X���
�+K`T�*>,M�����dSOGx�@LpE�v6��L�����DH0�n�+[�l���#���|�ַ����S2���o����ͧ,&+)���3ͬ�g�&�5����� 0h6��v�cq_#��r�:An�U���ޮ�y[UY�2V���i��]a��}�X���T5���.�n�����5*�SzF�M��^deW��>��W+�F�2Y�-*�c��GW>l?R�w/���.��J�����f�:�xcD�r����N <B��A/L�^�K�^A|ټ���̇�z�,�Ӈ33g/�{f�N+��Ö8�ROׁ D����� k�d^�C\�����35x
	��