��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���X���S��p��0���靻��2]��^a��C}����{�dHjq�9o����2�l���n������P�-���jOpg�k]��[�h���P�u�	ӂN{I@ :(�L^8��	S������H%�q����l�'��}� )� ��e����ũH�=��|'�n0�!�R�;Ѽ��-��*/�
' �4+a�'l5��� d]>v��so�;B@�&
�[U��F^�N�`�k�Aӵ߼M�C-����2 �8�!�����S�\W�e� )�r��u'��ߡW@�q����1>��̎S��������g4���-�g�ѱ7�Ch����-�>���$�7����8ruf�l�}��'!��5z	��= �*��Xк���`2���?�L
,v����G�~�Ҿ�-z�O�F���;����og���v�X,ͣ��r��A�M�K�l�V�f*S���H�e$n�)�r������(�Z8�����@��4�ќv������ײ�A�X�!��a�K�f�Ԁ2G'��4�>S3R܉��1�'�y�a�����o�
��� �X�P9���δ�)�����{o/w��J�-� н,�a\��~�~��C�����z�b�Z�tv��W�"꣩C6��g��k�#+�h�@������	���hTxᒟ�rQ`EO�>6i�|)#�"�a�_w�C(k�� �x���}��oT�+�omQ�� ����������Du��?ao�P�I�4\(���L�)�y��4�/�u������	���XS���2e�'z\��D��lx]�ێ��4)zim�q��
�Qxh��l[����<��xK>b;�Tu,*��I�:��0ds�E9M�-�S�P �I��V�Ѷ�nG���BF&�		�vlclS+��vL'�NڜvH>ʢ*�/(/�u���.��e=rħP�p#Y��.Ey��n�º��H9�
hM')�K��YG��y��śi���+�H������6��_B��8?6� �z�,�^�3�Z�E�{/`�{�~��cRz��)k�nO��G���P��[�[��H	7Dm#:����':��`�y�]����؏�N�#��U4K�d��S�g*��Y� y(Zi��;����_��]B#1��s~"���ۅ���R:� 3OV�͡,�j6u����:k&%um�{�6GkjbK}��DA�����]�|r�i�6�+z�X�8�*�
�b��G@�?Q~�\*�k
��m��������6�1s��S���{ݺ�[��' {��<��_���G�h���8���ϛb?7*{B���3��Yj'�5�0��kB$�v3 ToAfXn�|��X����Z�I2�PE��>�E!��V�߳B��	���J@���/a���S�0B�2����m�����Oe�9.�`m��Y�>�ˆP_{�T���`���8��@��,2kc���%}��5`ጏ$�F�3�<|�ֳi�]��q�>���N.�./���v����MKI'�qt�NS���G�GTſV����yك���a�G�D�z��I�l��UW�֮"�nd�N�9�'�3�����!IN�w�����ȧ#qM���Ž<�C<,;�j�.�>�e��^�d~�1���q�P�Qv&���u*�&
�3`+x���c<�6��񶔌м�o�8]�S�tc����_ �H�(%�N���v�5W]Ä
�e�<R�ؙ�ƚx6FCT�V:��Y�rJU��,��]�O�����_t��T֫��n�b�X=��$7������)�鏔(�]�w��W�}����_a�H���F�)%�.�x;�`buUBWM}^�GhF'�00���RfC�g��70Lr
���0��ղ������!.-�;��E|0��}r�0�0NJ-&��>���φ�B̸�p�U'RB�Mـ�C�����v��h���>������_�H����Z��i*�}��6atOgEUv`A��\-]d��6 -k@���b�!���u[������}�Į'�5t�_Ao�2�f.�\���su��圙/�K�m��	e)+UE;dє���k¦V9X���yM�2�_��U�[���2dM/][L혣rPJ����g{���aI�A��G����'J/�[�# %�pp3�!��?C�ayw����<�/4§|G��{�ʖq�'���y�ڕ�g�A�b�׭/rn��y��ŗa#C�����$�Pr��Lփ*c���/ղM��%�{c;tj�Y%��!�#L|��$ps
��N�C�߭��;�'��nz(Xm�Zn�.~����=�J�㡄!V��� �{ퟧڻ�X��`�-T���l����
�m�.U�BMq��z1e�T脖��=Z��y�n|rf`}��A�Z�穠qw��j��$.�O��d@Uf��~�O;G3��*��B?r�gp���p^�DW؎#�h�-
�;����UŪJ����O�tp9���IIc-�����T������:`��y%�g�J��p�(���,B�j��񾔁�)ҳ�����tN,�����s�U�)ĥ�4��,/��h�K���������_���<e_i&��z�ppS��e�V��9
���<I@Jⴣ�MD}�g��B3-N�%�Y���C�pL����R8�9��\3�� ���^��0�O����d���~�(�8��y;�����S��ko�S�i���q,%�E�P�f�Zxu�@����>d��^�օ�^r��c��~�>wF�������ovH�'�"�h��0b�K�1IB�����eD��ܚ5����vn��)���*3CA����~K�V��������=�Ԍ�v3��I���`�49}S<��n+�ꎩ�ģ����m��CS�`&�����&�8���M�R�?t���9��4_�� 
�k���b�� -����(8��~�k�6����_.�+�#OYM���(	�y��'	s�
q���ml_&ym
���XÜz3�vc~܃�	�� �Q�u$�������4(2�i</�U��bM�H��l�]� `����t�J	�hrl-r����,����ҟ�����1��(������7݀����S5H�����a�g�'�Ț��!a�� tW|EZ{�-E�'��S����Lsd]��?������L����Ǚ��,�X5A�b1/�^�y�늎�M]/4G��ug�x.n�+���~Y>f�Ag�ur=���O��
[�]k��ǊG���Jl��:Q|y\q
��r4O@�5ڪ��9�˥�J�p�S�]��ðJB���>���姧ȧ[�]�ϧ�y&W{����УP��ⷻ9��u#��A��;=��\�n)$G��@���_��b�&�1��S.�>�*�����Z-��=�+zJ���TF����9����5�US�A�ó5�ƒ��~��kn�jHˏ���y��hƙf�c����;�r#�"_��^E�h���]"�d�fEG�&�hDy��D�Ϣ~��\�u9��9�Q�<�X��-u��CN*�@�S���[X����e�0`j���	�xx��;�H�r�5)N��G�-���H��Y$IԀ��v)�Y���������:�����2�~�+1���5z��k�J��o���O ,]���p��\".dP㘡�C�Ӟ7<�~�]����iY��Y�耂�'� h�mN�9�.��7)ۚ �d�����*eU���莺�Ȗ�(�R[�yJ���rQ ��~&����B�Zw��	JU����A��>���. ���^�)�'`Tr�&�� x�B�q5F\ͪ�V����h[����Z*K���(��Y^o֪��	��)9�(�!�L�i����u��#Tގ�I`���Ի�:�<��4%�D���n�7NνX\8�D�?h�ގ<��cz�R����.� w1�	�Qc��B�O��y���C�4�8
@r f=���0��qnG���)t���]M�w���as(� ��$�[8e<���G[Uhw1T�O�ܽ;}���ikp�+ih%t��0mw�y�gVq�"Ą�{���J����V���l����#�������ߏF�#�Ε���R$]B%*v'��)����ёU�_���2�2��i
���9M'Nm�ݢ ԁRg�͔D}N����EB�G(%�R��Ŗ�[��V<�\s�C'g�mML'ғ�m/�ş��Z�����p�P<V�U���S��N/�(P@kh�Y~D���[�OJR�/��\ui�;�)�Y��L��f-�}J.��'�5i�ϓ�$1����Ntk-%M��]��~�WV��h|��]U�,L�`�0�6_?�0��rF�	�9e.Q�.�!� ���!^�q҆�f��I�9�/�_�R�� [�����Up�P���SV3���C{��θ��:,�'?t���#�,n�)?J�� BCE��� �*�3���Ľ�H>tŵE��0��it�D-|���2��kH�ȣ�Q��7����7n�Y�� e�U�d�>���'�^G�+nmɐaӝ���m��N=�q�/C�*���,'� ��+8��ܾꞑ�T��P�V_;�D~i�*H�J��xi�\����|)�����y����Ɂ�;�o+���w�k�Hoy�+�+�+t�����DO�(R�OA���vN�Q�V1������&�r�l��u�����T�x�|�K�w�I�x��q�Z�4�hB�\�4o@Y�9<�rW46�ow�+DF$���jabx�h6!�>7�GƔW$���i�$2;j2	����kp���w�QW;��*`}P���S�ʢ��Q���v/YN��yԒtz�z!T�hv�2�v�s{>�`�W0'�@1���B����)��Zc���^�bc>��w�fJM�����y����t�iP�C[K	B*̕brƾ<3���NSa�b���V�:�OX��N�*;�麏p� �x��Q����;�=������k�(
f1��� ��3�	x��e�as�Ud`pM�(��|
����e��c�%�����aܯ���E��v'���*��X�Q*�'^����E����a��zh�8(�	@2������y�o_r�O�qt����������y�2h�yX�<4�$��iɁ
��J��H��{��M�����O�3�$�r�y��^�,l�V�y�U�=O�æ
.�l�-s���{���YR�Ե+\�f1A\%��q���%a�1���#��¿��]�����,��Ep>���\v�� 6݇��<��MY�M/��F�p)9���~r��j9] ��e��Nm��FZXڰ̵�Q{^S7D�� .<�^d�27��`�}y�ȅ�m	�2��6�KrPg��L'=Qz$�l���z�8J�?�,�q���}��.�~������_+�
�+�����MٚU'���_VX�ox�V�V�s�h�c�=(VM�4d��KrxX�jʱ�h�I�d���kϹ�gM-��aMrrJ�s��y���ٕ�n�������@��\7���9�.�R��k}yq]�/Ǉ̋V	�zUS�ԕ?�I����կ���%�Y>ջ��(L�P5z'a�����[5���4c�9r���p�%�?�!�.���$5�#�󞦓 ��"3��Нd���I��	[W�C����\r������V��$�ŗ����]!�����˕�������s�?�#��q�����vH(�����Wi��9�i:.T�y=oއ��GZNX߽Z��=�j+�q��1��s�&�i�@Gz�b�!a*�~�i"���y"Ԛ�:Z�R�몉V|Yj�$ �OG86��.RR!�$�,���>��.�A�I4,a�޼X���A�m��J<���VϷ�k��WUDul0��~��*�규���r�+сŉ\(��2��V� �%�**�^��Ŕl�	Q�ѭ�<���z4�l�U�S��8uWρ�{AP	�o�H�us��`}`�g	;%H���tilGX��b�:wU:�Yvd0� SZ��0�\X����Қ��{�'��	D��0m}{��t�Ě��U[��N~Áv߁ȉ{.E���>���Ɍ�3�}����!�q�
!���,��ĕ?�����n�82�oG���S3��4�I�_���((_�[����!�����)�I�grAkO\P��O��S�{����H�&Nr¨���Dc����$j�>݂���r�Q9|l��Ӓ�z֢	�J�����Ο���gs����	�8�5��j��gTH2���s��%��c�*s�Z�^ї2����HO'�x�C��F�:��6��E�ژ����>�J<����'q���;si�����6L�I��]
U$�;��CSSm��X����x-�� �(��˫� ��G����`�}W�^&�ir\�,��2�
�t4*�����3Z@n�����1��QR+=��.ë�$��^#^9�:��y�q��%gTc���<���Qa���ݿ[
	G5�L��l*�]e��s���@�b�n���G�4 쌉�j̉�K��5��ޖ�gZ���B��Ti� 
�15�(Q_�g~(��jY%�姚-������s���m���H����2P�f�����^��*i�W�fGf��X�6b}3`@�7&<G
��%9�<���5@��(	�u!��&@�.��W�S�4��6��/���"����D�i�h�nq{q���~u�lTrd�cYFH�/c��#L���|����TL�����8y3Ŀ�ʬL�b�
���BKM�\H8ѝ�i�XC�S��(��|:z��΢�Q���C�3������$��=4�g��!��vV��)������%K^�'�Ǩ.5���]��E#�̀�N�m�tU}�4
��MЖ��8��o�3�<��E�{���l bF�r}D�ek��6�*,�}�y/]t��;�r!���m6��AQf�a�"�-~w��7(����G����l�DHI��i!='B}i��t�y� ���m�T��Y ��~.����u�L��,���2���_�]�5�s����޿I+ �X��F�+D�"�xhA� 8�?�3����k(������&�(��߶�D)a��on(%_��Y�7��Lh^�B�LhfH�/%Dپ^���L��2���pm�l]*�(�ؾ�FZH�[�J_/
�q�)��4Ftr^}^)2��e=���䟧]id�	",��8q�!U'� n����E5�Z��]V�{��r��0�Q�3���!���X6�1a�c���[:Y0�|C&�/������\ J<Ŷ�Z<�����(ꑃ]��U%�d���t��<˦�mX�X����G�`�.�tv@��VA �M�|������Zv�焯��+;3 t	D�����{ǋ^<�:��paC�dd�@/G#���Ǳ�e��ź�L��%9��`Cco*�e������®�����:�LF3���%���NfwP:����s*��(��A#\]��[�Z�_KUT`O�f�1���>�����q�=��PR��N��D�g��-�Ш����?M��S�N>R�C�+���hX�1LǤ.���	���GB�[��X���S���`�=��B>j4��G��H��bl���I�si�3�5?��a�Ѵ~
=�[Ke���:���J��n1��V�@�kݵ��:�``@�f��NA�H���
�dD��	��b@ma�Ť�1�c�@���T®�("+7~���n�Ό/�^�˅���$D{wa�9[l�B��C <��zb}��{�8��<P��1�Ŷ�P����G�W����v�/��ay��P��C�$���^�5�I�3�T,t\�:��mf{�%�C��E�PI{؎�G`��b�]�
���Rm>��6E*� �#�o6F~&%����we&`���>����xYv:c��o���}~��w�5��GBK��`t縤�8�d��e��Y�"ѥ�H�vc���֧�u�<��b_0<0���e��իZ�/�(�W��f�ꈾe�@�֗��K��ρ�"�'O�3�3m0����*������w�kʊ�IG���QVn$PI��EV�:<ǂ��z�T\��1���h�ɼes�8�3�Tڌ���w��έ��S�s��GT�?��d�N�U�\/�%'���PB��d�Y��oxtc���Rt�+K��Y�m�r�4����O߫g���wԝ�#O������M�(���"�q䃟u[_�p�/�>������˛�z/"m\�hU��o�J����d�r��B��O�[�=��x�s*�Tg���) V���3�(5�|ҥ��]��@���v����A	`o�>�N^���j�2[`Ï+6B�O�|4�����P*�[2�f� 2̡���b��k���{��2�#'�e��m�[<�CJ�i��p���F��1:r���#�U�[{�D�v-�����'��;��G�����Y}
�/R�H����<,��5u�'���?��H������N��+G���T=����oi	���QO��sng�	���%Ҷ�4��yf|�d�4h%uHva�IQ��f�&����k&ğ�ZU�|�3��ŧ(4���]4pJ��;���T���i�o"&��Vk��{/'*<�o<zo/����5���šZ�4dB�}�Ѝ�.=c��a{�SPW�Q���F�)�E����(�NSM���V�/��Q9t���r�͢s��|Uk�� 㪍]�V�J j�����P��N������r��tz]�`�%m�ci�J4uIל��Z�g��nM$]�xJG�j֛�G�U����[c� c\Q	�����ҸD{������d�>YP���Ұ��Dg�qD��пQF� .[7t'6���v���h�	��HQ9/����R�g|��W\�DEԗ1�*��`4nXj5V�XL��f0�M�_����"\u�)��` �Ϭ{jϮ��Y�a$���ݟ��Zt�`����qCȴ6�X�)QR�"�?��wĐ� ����r�s�D��?3t��>�4Gu�&BY�CE������Dӝ���?��_ ͸�G)��x�����m?#8�7��_.V��JY~V���|#�lE��k	���b�'���" ��t��d���pi�Җy�(0*_��p�9X�AYj�ּ�=o5\���a�� ��;\fs�΀��5!����Y Ձ�	LXT��CdVc���s��"��z��'�͢�ү��c���,+uգ�>AtYpQ����MHAP6WŹ��KuQ=ia�?�|��4&m�	x�:��^M�(-	���K{#;��=T�9�+��+j�;�q�;��N)����^h�w�cg��m�tі��~�G�*��䱫����-�|����R�[/�p��� 0�V�>V�W�GO��	����7�?���F���:�>m+�[�	g�i�-UxX���B�%$I�fhP��#$p�f�@MX�0#�ԟ�Jd�{��F���^*�j�͞�0+��zإ�؍�+�z~�̸B C�s��0}���	��ke��Z6����_��oD,��H���"햅�yh�8��PoX����^���/M`�;�sq	� ���^��G��ĦNHT�M�������/�˱L����!�7�~0��:�e����i����;��c���4�{�~Z^Z(.�<��Q����I��J��
�*\��N_q��c�hR�X��~�GNL|�&������z	�����b�"Rwp�WV��ʞ=߮>7�b�
D^{䌺���򺳋G�_p(놠��o�
�%&)�W�9��HG�'j���w�B�(-���L³˽��
�c�]�Za�����+4=�=L3��䷸�6Υ�:���6�5�aUt�R�S_^�H� � bU�쥧�Q��Vvn���^Z�����̌�
��m��􃞯�)�5�.�h<bf�̉�Ф���1�{@l~�a�}"
d@sЍ쪀s���O����@���-��[D����31�ߪ���l�L�J8���y��*�o0�j���I�u�N� 7��WA>�?�a��I�I&؏'P@ȷb7FZ���\4dj_GX^Xl��MI]�67�{��cS;$��j2�P�])�� �� H�<s�g�C�{�w��	!�pВ'���gS�/J*���;��Eq��C�q됄��X,�_eI��d{U�D"�O_�wA7��gT�2�x%�拵� �K��l� _�#@�d"��0�*f��=-�Oh�m\��1u�;K��DSk{���	�~D
-������qf��:7DK��7*K{����0SgF$�U���r��.H1��{�:��ljz�����!K�L"H��E������ýv�#���Ps��N��_5� tֹ�/������6��N|E?�!AK�u8$N�0��iqKUU�e
8��$�c�$D�h���A6�B��D��M���ׇ[��9f";�^<uBY�m)t�I��V�g��f&�o��w4֚wz�q��.����QvQ���y%��Âf}���'�<jE��sX�R��	;s�=¡��t|��E��{�}
�1/r���0�>��Y�Q4�}�B2,Uiu��9����$�w�V�eո~ƦB�QKkGD*��I@F�S�M���\G���FBݫ� Ty����?d�8�t�2m�& }t�ŏ����"+�m|k��t���kɷձ-� !49"�j���`Y���nJw�LB�z+�˭����ׂ��h���R����Ҋ-�|Kb�G�P?gX����ʇ?wA����I�]i�$�l��<t/P��s!c���f�D�t���4v��j���k��4
������>-��Yܯ#�ܪ� �ݔ��ӗ3n~O������qM3��v��ΉD�A�7;����>aA#	~ok�L�����@]f�������v&��]�'����!	N�U�˭�Ra'����ܟ�ˀ��q^��u"�U�=�w�#�� �g��������P�k��-a#IF����,����]g�F��f�����rҊ&_�s��+5�q��+���+0����r|��&�VO0tg-�F��7��m=[֜c��,�����d�sZ�4��'Ԅ�x��鞮Sx���ﺊ1�>��4�X� 2��hI�s��6F���!���}�򯈰��Q��5��+e�_�n!ķ�3^�y�����uDB�̪���v�D�jZ�d�V��n�1��a �Z���|)�lKq!�m6���~��V�B��tP-i�3D39��Ci
1�z��Y�&V��΃���h[�|j��u��}���o"���)�
�=uhp8P���綣
��)��!����1Y<��U���g���"(�,y�f�#��o[^��� ��_�f������%�d���<d�C��B��ȧ��,���UGs�8s�1�X1USx�
)������GD����?�g�r��tt�/��-8
!��S�Cp����Nm���e3��oĆ˸V�B��^�J�vy���,jb�� u�0s7�U*�oa��b�r�� 	\�]�]�������(	R��3�~����e�]یX�HZ��H��[����t��n���9Z��)� N��p4W^2<�]��h�)�r�r�$*�t��M�I�j��#3g�q&�N�
�Ml��)��ai�c4t7�f������ ��JKM��"E�l�=�+cm����A������@L�v�%ގf
	wz�Rx�z�[�,�ӂj�Q��N VҦĥ�+���ǚ0��9Y��pi�aT�[�D��5�u����!p�}��'bv�tM�S�E��uL^���=��a���.�;x2[`�[Bm�}�=�VX~/�{K<��M���������r�Yhs�4��y�k��r���g�\�B�Wa�� ��qҋD⦀�wS�� ������C�n]q�D��1��9od��#�r>�9��F�'�\�	�k&$֋�)E�gg���[�ǆ@�'�"��G�%W���w\1����[��7H�h����$���.�Sc/�r�>�p ӆ�p��k ���e��8�r��Ȟ|,������=�-IC�j���%M��������;B��Y�و��	���@fsr~Ri�8�3�'�	��X.��{����:z⼨H?����J����N�&�(N'�6� ia�z�S�;�vZ�T�8����P�Q;J���!E�	�[��4e����0Χ>/��H�!s T��B�qQס�P�%��Cx�e�0��>i����h�����]�Xz��D�'��dX�<��A��_n�*����PAw��G���$���7�3���H`�vM�0ՙ3�ŠGz¸{ON������1�p�g�n"'�E'�# ���_��1c���66�.��>� �wg�i#)���ZZw���0)Qz�(�m��aR%8��m�]!�f�V�FQ���\i>�L�����~g���Lm+����W�{Z�r�=4!!XLb�����,��)�R��eQ�*�ĵ(�҇�����>�R�<s�R�P�^�Sl��JD�%���s��E����P�U��a��
���\ P (����ɿ�ݭ8G�>6��������p�����-����h4H<��ս��ݦ��5Eq�ԵމCP$�! �wf����A��c��h�Kц��PH�����f��۫*�y5��ut�(�����,+k���MS>�j���!4\�\����r����M�>fsK�5a���*�\^4M޲� ���b�\�9�x"]�n����zY�����4YeM�C����=e�0sd� �d�+���F��-'$c޶��ّԯA/�b�䠄���*�d��>�i�U)��rZ�1������F���C��������Lj}�h7��{�����=��3�0�5x����@��%��&͇T��mk)��g�8Q����<����"�$Zn?��:1��r�[��
�����C$`����h]J?�,/<6�B_�vDi!g�,��'��L���%�}�TCIE?0����_y:9?$a��l֓>������vm�Yf���f���8��{�"�R$ny��A��Ѓ�\I��_ U��Y��2o:�A����B�\h@
�bφ;T�`��=� ��n[Mq!��.��r??�3�Xu���=׃�~(� 8d|���6������;*��.��S{uVS?l��[����f����"���$�`nh���{sܐ�t�줯��JQ
:��L�ҫ��+������,v.{Z�e?9h��>_�%9* �j�㱨m��0��x"kq۴�o�8�~�9ޏ7�B^!{�+�QAӤ!�7�ҶN��z�m����>k^/�>�I�إC�����(�s�;'�4W���<D�5x��,nm
z�P�ƪ��n��Z�ɿ�2Q�3����!���{����H��;,�.�D�"�,���z��ﲲ��h!(u���
�����Bh.�CJ�����Şֻg����?��j[/�pw�U��H=��Ǐ�膥Th�f���{�2����7����G�z��vҾ)_�~�TEr'3�+⪶W�{��r��������(1a?�Y�E�.�_�".�ߝ�jxo�V�9�<, M�޻-��JM�f�F����uNÀ�x�?�qlPSK����۹ٜ}o b����K�Z|�M{+��)�Hbʫ�+�ԯP��?����+���3+�����j06юl��¤���#	����|�٥V�� �oN��wؓ��B̍� �593q���.t��f�d<�/V��sJU���8��5�l+\��F񬇪��>ߗG_�/�1���4�n;�$</hG1�%m6��5p93	xj��kV��1v�wr�����&wn	@'Ǎ矑�[�K�T�img7��f�%V�z�-q��>uP7���D��$w.oX�7��!��*��:��X��~_f��A�U��yVY,{���,���U<�1��d�{Pvl�i6��O�j	���yt�{���D,��q,�Uװ����]��,�O�֡܇�+`���:�����{~$��e|R<�%��R��'X�C�����:�*�v|�k=x��|�n2��F���{�D t����>������$��C�=<7����q��f/6��M��C��q�/:9�����A �8� ���׃�p����S�
�@��N��c6ll�t�JQ���3��8ܵc�ȴ;,�����<Wݝ����|N��Ô�qҗ�A�5�3k��B����H1��<�U��rؽd��ÞV�5��USϰV��CD���'|l���Q����:�Db`�.o=�Fw�<���@�W6G}�!@��l[��!L�u�Ϻ��|��������٪4���ņ,�jH�Sh$ �����ؿm��+�P7��v>`�6�=��H\��i,l(�����Q�}����nN�t��P�F�� �
7�??n׿�Q��b�!��?���Y�`��%����[�M�\h�
��o��]V~�"���{S��}�/�+;�����	R]�_��u5��-^ӧ��G6�FF�ڛ�d|	�b�y~�q1����q�o �үz���1��ƞ6A'��X��e��;D���"A_�����e�&G&��q����N�o�42a���\-�BoͺT[�+�cw��X8G�˫8��8����pXw�pv��'��=U
V?:�$94��pCQ�v����hv��c���_�IH���9P��E�[�	��`��&׆�=0c�ݶ�G2�5�.����y��k�B�3Fk:�p���fj2B@����HKtߘ����6%)ť�+�e�v��k�Z�����,���4�1�