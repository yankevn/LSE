��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q�����b��� dԍ�,$���(�BO���okfY��%�O�%%&4X�_�1���� ߴ�
W	���V�]�R�(���+$�,�[��f�\�!hv4AP����qF�*qH]�������b��L���G��@n�Ǥ���V�����������F4��P�&[�`�.��[�^��}i���q��a�<��2Ҍ��c��=��hF��`o��SGz���-��U��R��m�0�9;����=��h�@\ZHLl�,3Nu>�J�r��Rk/�S�;��i'����f��$�oE�{Sz�2�2��M�=��H�T��(}��k��=�gx��5gZ��eďTU��S1b��ذ�;4�<����`d�>�[�_��(-f^/�(�EZ(��g�B�#r��>�;G��,8[U&u���c�����06?a�o�wϷ�чx3����������eN<�&�'�;��� +�o�+v�~aD����x��QiɄ�ɶ��eL-��F��ǹNǶ�sͰ_���	XbQ�a��v����Cc�"r5AX�g9vk�OްWz
rcI١2��O6!��򺳞�Z]�(y~�����M��,�[����w�"��^�#챵�5�Ah!n�z�}({����솫�W��1-/XM�&���)8h�0nP��c�PP�b����R
(��-hP�����%�;c��3����H0�D���sp��n$<�8�w��!\R�^][���и�ͤ�*a���_�3S~βO$�y��>� Q�_B���Xfȳ�c��D�ùh���
�4I�������j�'��(��ϢH-Rv�'�8��I��T>D&&v�#��-��BΆ�R		�� l�y�@}��IՖt����EO8�*�౸ඩ�y#��6����I<�H/=I�f哅+~ �c1��ھ������|�ڍK��e�f���\�������5�����jd_�!�,���j�_�`�	�����g(o���ٰ�<Rl���G$E��d�;U+9��;m,+��s��㒟%8h�N����fF�x�������t����ST��`�b(G�c:ו�<�4="x��L ��y�#��XGG��X(�mX7���Sh�f���T�3��#)Xc}�^���˰�B�(�t����a��Bz�%�},WS�Jz�E�i/�9lsS� ���̑��c︕�3�w��C� b��peK�{��Iy��M��Tl��I,I&iP�	��}v�|n݃C�A���D�%Sm�^gY����z,�W�͞��7n/��i�Ѱ�G�6�c��-�ys� ����v�q�퓮+�>1y�s�?x5����y�Z�P�����,�h�v�[T��F�������i��W�z�녯�؟�:��ަz
���R*����͍��|��i��J�P�PuoW&�J��Z�<$s�v"F܁Y-v�<"6��ۘO�Es"F@>����xTt��eҠ�:�l��H�	��O����sTD]��ޠ���Rv��(-�d���i�q�d���0ٶ*u[e�* W3��f�D�8��',w�ƺ��>��>Th	��J�E�ɤ�%	���@Y��c�O��ewz3���]�~J���@�L��Y��Ƌ�L�� ����EJE<
ȗ�U�:/�+]̮��	C�0�TW�p�_q$5���1�t�����s�Ϭ?Q�f9C��L�g(^80���T���8�"�­�f��j�F�ȉ��T�T������TK�WT}H����!�1�N�d�:���[1`�c�X��ϱ����+CK��l���U{�]/+1���C7���gq>�ܭ�@!M� n*��LqԌ�e7�S7FE�V�{�²�eCb���9-���:x{+:�{9#Zj4u�YL��	G��j�.Qf�O��-_;��Dmyₐ�
	��J��Ş�?����{�6ߛѭ=$��3r�~.�f{��2�yL�2�!�j�M�a�52E*?���b.��-כT�sR\�jK��;S������3;���U�:;�	qOZR^�:�A�o6g����G�H�`�Jc�a�y�6�B7 E�F�@�iyχ�V�m���$rjTTA]�,m�=�<�屛<��*z�L�L��њ�Ǵ��gb��t��Ԃ��I1��"�����Xui�l)v�[�ɼ��i��٧Ē�M+����f�!|&J1�N=�)�@�ܜ^�:�A��:~�2�>����w���#<����.���sQ��kS�V���1�ޖ�s��,�F������W�T2>��o��"U���Dx���1 �)��rW����<���ή����尴Gt�^Yf׸�m�Mb	Z��Jl��E�<��̅Q�����<� [�b��s"�o���G�~jK�n;Ey�����&a���^R�,[ eI�(�2���n|��%���`F+\uk��ڡ��+x�)&��샯+q�}� ќlub���O��%�w���~9�z��P���(+ס��2�����Q��[Wι��P�e R�Ή>��L<�5(�n�b~/+z�K�>�(j%���LL��ؙ=MO�n'̸����Q�5/��s�-.�[�I�ڃ���j�p8�5�D�k��͙A�$ۗf9j�ʤ�ԣ`M�$�ޢ��$V�x���'hKޓ�}e˙Vw��>�y�΍di]vь\���H�Р;�F����n�G%=xf����$:���W,hM�`Y�u�x�^���;�C��ed�h^;�6U��[4N����m�=\��Z���K��Sݐ4:^ ��rk��r���?&N�dtԣ�VB���<iM�ek3��m9ȑj�p�ܣ��nCm�LY��`iMx(�H~~����V��Az�Rɉ����&][NO������l��ר�-O�����-�V��7RRT���;}�J:;��5+~�.X��+���9M�K�d��I�O4Ie�~l�$cL,�=�����ơxV���+R_�&:n��)X��2]��[)5Hkr;���E=^��ʾ�1E~�0;j��m9���(���R;��w}תA�X�+YןnE���:Ľ�\|�I���B��k��4.����������Ky�	��^��B'���1�1b1A-z��d�ЪH�,���Ѕ�sng���iZ��:U�Mיzl�̻�i�T��y��*�_o��v�Ӄ�9��[��ۀ};:�k|g�m����5�Rpz���,���;�����`T� S�~�8J�W��jY���-=2��>��n�;�9������Q��rMq�7tΐ��.�����3v�k���˪\ۺ�j�^M�:
6o�~���8����lz��|��X��Q��ne��tY�o������X�Y}���0Q�X ��'�6x4r\�W�&���
ah�J��j��L}C���4�M0� E��E�+uP�ߞ9�>�"���� �;�H�:�1���N�CыFQ���N{模��헯
WP�ұ\?|G�ee�oa)&��L�����/a���o�0i�e��ļ�3�kZ����Kl8��5�e ���\�[���i
����\ł8�C8��,�%���%�8淽؄��:�YA���X��묣z��Vz�HaIL��w-�,� #�ޚ��8��9�#v��/��k� �؅�6]���w�ߌ�5�`>�-���dy&Z�I4v�`.�!��=���������*����t�p�27P1�j�pn�!��R��s
H������KQ��������/�{:O��L��tP�^D�������	�w"Ly��&��b�U�{�,�ٽ�ve�2O
�� ���t���]�c)1�	$�1�T1vD�^�%($�?�GL̲��j�v?'o*���n��ӳѧz[�y_�p�)�`j늦j�?�Řwн-���t��c��>v�����];$;<H�ג+Ҳv�v�<����Gh6�w`��9y�!���Ò4�I ;������Q��@����}��7�7Y�50��k.��I��6�K������$3;O|kN�_]y�
7nJB��7hUd���{���������l��uP����a钲��'��˶9�ib|K^����b�P����iOhڰM����eчR�)<�������S,�rL!F�$Qo@F�WȣX�8� .�=�^Iϥ�՘<r:ף&�H�v8	vz�`�0%Q�xk�"6�a�K�-܍3+NIT��k�Vb���~X�mQ#��#�]�,��|����]���0�R?y�EB8������H���fm�.���̈͡ȴ���E��`R���Xe8��y�k��S�=�:���vk\^�*���0�Aрr�8�Lp�Q�nN�����1Wp��-�� �\p�6\)�����r���Sڈt�et��8����+�Au�M���?�A^J99��������^Ȏ-��+��a7��OR�	�>kA��G��
i�����������/��x�<���g�eЛt��j���Yc�-Ǚ �SeNƤ���ж��&_5F��w?���g�Z@Ƈ�1����Y��٦�Ӓe�T��i,���C�
v��B����&(�3��ׁe�d�¬�`���(�]d����K���srP2 ��&򽙮Y�q�rF&��z����Z�
��
эLP��	(E�����pS�@-R�(/��d�� �|Ĳ����7�O~�����U�-&df�끥�]��ʎK�;�ߠ �UU4?m��5Wp�W�F�fO:�]r��u���Ww+�CG��a��]��9�`����Dl�z���]���s�1!��qjL�v05ۤDq�r�KlP��5x9��΢��?B��\���HH˗�yh��;?��{İ��e��܄