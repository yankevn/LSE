��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0&Y�y�OX�GK�!���%V"7O��r<"p���6����lb�E����<���x�@|���.�����R�Lu\����1�,m�K�͢���i�7ˤ��)x3G7�n��}Z	ơv�c����lG�����3�lCXZ���Y�Hh�
f7�6:�3.2j�T��8���4l[�.�޶�w���9x��|�
�;1j3��N���!����X���t ��!�,����"RfM�ɓ݂-����4�Z�'n6�,���{�N��z0�oAwuOBD�n�׎*,-Jp���꾐t��	T�M��d��2��K.�b%3�WeXn�y��%0�2��^�"G���b��KtA��1a��o����\��Qǟ!��ώ��F�*㼴H��@�&0�Y�PY{9�d��l���I�|v��пs	���Z=��nyFrd�;?n'ݤ�m����f�dT��e�~k����0t�	i�$��T���($/K�K v  W�tGJT�!��d�rIL�Fљ]5��.��s��GX�rp�)i�d��Db�=t�+���\2#���޻�s	�Y��=�-����t�A��-�)
��>X�Q �̜@�l��19�Խ�?�f���ٰ��A�a
S�e��G� ��H����
z�����8tcش�yCDXxY���R��E#2N�Z����v�	9�f���i�,O��. ��x��=��X0�.g	!y`���3d|�2����m$� ��Lʬm�`��
��T�,�9�X�\�G���,I����ӏ�A�rkY���,"�V?2�(�X)��ñ��K�y3�1g��!)��
S�;ȕxm���+DU��C��|��ӄ!�_�p
�������W����ꏆA��p0!y��c-2�_��"[�2���E�e귆7��,�PRq��������w���8�@>}��l���C~�	�>���.{�S�.�4`�v��s;Lq<쒢3�7"DP<�j��'�p&8����c��f���jh2���v�[���K�!d-a�u��<cه�=�&���<�)���s��
-�G/;��Z�ݙٵ	�z��Q�T`��������'����գ��ŕ�ס�M|螱��?��6%{�t�-)���&Й�5�c'��2�ћ4�`���_��4x�le����+��$�]����N�ʍ��/48g/dGq#iD=O�Hyz	�ղ����!�Xr���nH��G~cK�S�W$c���G`��N��'�-�F��޾��҂��[�۹V�������#���*!�d~S��2j�B$�{D���IN!*����`e��6\-V�� 7�����25a[BzM�6Y�7٨^D`�U^��b������bQ�:�H'���Wl*"��n��kF3
�UTs6��;��B��Q���*�Zv§��\��4:��6!�⪓�=��5Y, [�Fv���":�i�u��;'�t�fE�>s3VC���"��Ӱ�X�Y��D*c�$���i6�Ⴝ��D�SK$W�h��U?���ǣ{[/�2n0����$G,��A�!۞����Ǎi�������o����C����Vq���<adߐ���:B��~��͎9���+^MH��y�Og�_.��m�m�2q�۝N3u��;�_b)�Ǐ޹�@]d�f
g5���я����a��FA3`�1�q}�B�*q�S�@J冟$����_��䑐ui[�N�^�\O.D���R��`#6o�&�۹(���N��}��m3̲uDE8x�M�b�g�+�y���#���M��wڗؽ�^�É̠*(�BI�?�1�C?1��,#*E����9f��;Q����sDJ�n�u"�cۖ�Z�I��'��Z�Fr��l�!�ٮ��$A������o.��]�8~��3d���>����x
蹏$ؚuU�ܲ��￹.M��/�V��fYC�٘�_�X�$��Q^JS��<I���`J���#o�+Єi*���hp�����.�i�98�k�݆Z��`�c�N�i���ͼQ�bl`�]D�kbt�}jQ_9����Xd��ٿ�p��G��!-+�}�)tKa�\öXj����yo;�ݧ,Z�N�O�O٬���9h
sr���K�}5��j��4����I{�Cnuȋ�|0p�<x[�)Y���a.�ĴI7#�U+@ZkE"Ru^��M��'H�2�":  ��������n�?���0j�g%Uك)
�%����s���Ϩ�It{�̜mn�B�r�?-�j{1(��x�+(#����A�n�LQ������rOu�˛�/��o�V�3bAQS=ǣ��E��֎8>w�Qz�* >���C|褭�$�w֔����L}%����#NϚ ���6ͧ�Q��4Y��q�p��Ѵ\݀��BM/�ϖ$�n���/��}(o�O-�� �sq�7B������Q�wc��/�.�F5�%Ϭ^��u;�����GYa�w�O�T<�pva��Y$�,��}ΘrZ�F����:�A���E�y�y�Z��H�Jx��90�@��5n�Y2��?�<~��� �3��G=���(@Or��Z��E�4�f"�qB�?����߂qP�y��@֕H#�L�q�f8�=����%��{/9�c���(k���,Q�@��H��b%�%Op���5м��6گ��\M4ϛ��7��N#x[��1XI,[*���35�|��;S?�p��)��A,�Q���?�C�� B��M(G9�(w\翅�'��k���8�8������~���+t�̻��5�Ǉ��c��n`�
��n�Jp[ E��xJ��[�g-n�W�5�Ս9J�,EF$���G w�Ҽa��+Q��PT��lY>��|дL���k$Jl ���i Kq�m���n��G����k���c�w?+��hT<�F��/\k��J�r~Y�`���_9o���=@r>�!z�4ʝ�>�;�)�ba�?˱r=��,	��47~r�l���"a�Ut��:w���|�
�p`����)g��DRt:���۞Ԋ��\������br��H�eM���#�*����q���ii�H���#���a���gJ��N�f���������^ې[�{���6<ad�`�z�(���^�.8�<�x�uj^]�[OI Lx�2K�fط��MG��C��� s @�x�s<gu�8�zY�`Z4�5Q�nɌf������@f
�����p�>;��ᦡ�~^�(x,�Y��լ�`r�R��O4�s?��ƛ_2���$m�6	��.�NےNv&��)8��� � ��rX|��5������}ۣh��ʘ�����Xؔ��ՙ��t��P���-�&B���|[8���ډ��T��r��lR�j��ToE�2��5E��6��zXM5I���M3�����&ݘ�C#Ϩ���/e�Ń��Y����(a������v��z]CD$YK�$����԰F��>0���D���/Ei�����[��3"���󁐦Q���F�K��E�'������o�+�V�,re���l()�M.��Q�'����dz�oh���� �˓�e챪*Cm.4��n#$ƶ�O����������+C0h�1��N�˳7�ܝ=�*�����>��Bp�P7��I��?���YI9a)���(XQ������ ���Q����Iِ�K���Nҕ�Œ#������'�j��E�,��_��x�T����Lf��d�nV}�b��z@@��z�j6}  �*�xp9�=<)����H��F+�\�>���n.��'�����=����*=f�Xg� ��Y�ڂnS�|��֩C :���o�d�;4�n�(��4�]ٌ�-�)�%X�q��*�2k������a_D�h� �-�N��e�fQ�B
D��#�����|{Z��p�Z^'p���hT4hy�)]�iR��ȶ<1�x��Qv�{KN�ٟ�4���fw,)Y��?p�q�k�"��s->�����UrW�=4�?xAH�=�,����U�����؅E�	���-�"��mxn�gu@x�|q��.��]����&1_��14�!�1����-���� 
ٻY��F�� ��	����D���Fte��@�[��~�T��A�
�r�`�4���2�������!Qv�.�_��j$cg��;;,���Y=+@�����<(h�ɏ�!)�l�&��6m��߰�>��ph�2v@dU�4����%�[���|_���fxgl����<ϑE�D/ ^���[�k��?�*iCڃ�6 X=�*�.��Ι���7p����d��w"cV�4��f��"�AR^d�6�d\!3	�㥟�5&���;���f ��>{(0w��!_��"$6�|��R��VT��g��/�i�x!�Ux�����t�+�ʱ����8��_�w��Y<DL{��_���	�Yrw���l%�`����(�|���*�z���GW�g��禒�|�
�߾8�aclG9�#�v���n��xP���AEDU��(hY�]�-�ۆ.zz��l�{�7��@�*����N��fr��&jS�ZΚ &Ԏ�)n
S���.�ǜ��ݤ��鍺�t�X*��}�����?(���(+ =�[9,A�CO�����Y�3��g�:c�Y0��<�}���vXY���8����Q��}��;]��OlY�x�yI<��!Iޫ5w()[��SS�1���۪�2�Jq���C+��7�ߌPY�1��&"�X���k�Fa�i��5c��Oy���	f��gv�K�KB�D.�k�d��O���Pb�#�Db�����9_=�گ������ ��ˌ��c��X!��¦0=��bg�i�R-v�h5�������h	ώez��K��ۮ�PV?�_�6�2�����h���U|@��7���~+�f
�AB=bo���r��[�X�B[B�`�&���Ύ`d5��D�<�G,�P*d����j�I��Z�u�Tc�3����pR�A��F_<'HR��ӫ�̓;�6��|MMISά��I̲[�mI��}l�TsxX�l)g����4p�K�u�[�wv�j��F�ɨ7de��V܅��}MA��"v�0h�,��:/H�D����]*aҳq6Pv@�|K��F�y?�TK1��@8�nZ�#�v�Ax)���!ن�GVD J)�ܑ9��-�&!����cmW�QZ��Y������]�bk�v ���e��b3?�哕�����������]��y����b��H ��9��6�tJex�_>O���$:�ʫ>��o��zG��#�=�\!�1�����U9�Z�1��Ǝ��@ԋ�J����Ô�;�8ʹ��L�\�S_����Je���^ �h]gR�`/�s b��^@��>/�-S�������f���Yq%�K�fɆw�t�3B{�&1�%-j����9���aS������`8���^nEZM�MԿ���U����#�"���a����;u��=�-��ݲ�@RgL-|6��*͢OTl��-/�V�H�鞻,=���s��9�1l����݋�������5�3B����*�����3�O�XaKRT$5���Л�D�M�L�����O�[Y�5����]#vZoZ��f�=���4��4��ɼ�2�}6#��>����>f��?�8a*4��kڑ��f_�PBY���q��`�����|X���7Y=���]W���M ɦ�����;c�)^�ףc���/�Yq��M�xu��n~V_}�����i�[x'�ߚ@�6���B�N��~��o} �WP���)N7���??�$��6�.�#�W��D>��|:�8C�4�Yum�|+Y�!�,�l.�J&=.���W'�I/CC���\��~jv�'bc:�^�z�Lk��.9�I^��Y�����Zx��1�_߰�z"vf��
��yD޿��pΟ��<�j�|F-��P��cN�l���|��+�5D���~K���*sv�[�0�ܔ����6��7��:,��u�&���B��O����������jP��l��9�!5O�(����l�OœP�{�>Y�/Tjq���\$oů�����}��?�-\	�BрU'�Zj���M�?<|�z_@>D��cìv�c�t�e��7\�
4?\�;�lR��8J�~�P��
A�U켴d�@�q���PC'�a��A��
��8r[��3�0Qe6E�m��������fW�?$`ɽ	�N�+�����'�(y��E��?0<�]fAFA{�"�!�B�7��]�j����w����f�I�[_����[%3ɼ
*}�lO��Ӥ5��JZ����t�B�(Ge��_I�p����*��)�K�Nf�a[��i	�=TO.Cm�j�Q��뒆u��~�z?���ʡ�(*yA�{Ƃ~N�B�� L�� ����+����He�3���$aX���:f��QXIڝJ���K�GI>n�@������D;ݚl�[#��Q�E�I����2��Ƶ�[m"D�4��F.MseQl�M��*�9_"nq�x��������UX���oʙ�9�\g��Xӱ����d!DC�y�(4P֗��ѿ�w���4�=zt���J��k�����s��7LDo-t��ҜbS#��S��k����>!A���&s�ůvN���0o
+��*�.$��|��wO��?�Л�vw�p�nU� �>1({��F�����Ŗq�N���Lƞ��B�s4�̳C��?F�[-����d�}���vԹnj�W3�9�´(����[������و۾���cv�I�3�7rU�rq�m�ލu�V����%Ъ��A
����J��`7�+Jo�%{�E��VBe�4��N������5UD�U!�U��q�;�X�ب-j0�H�X�x�w;'w�N] �px8�P%���nd~
��C޲��6 ���VV��"���P}�	��
���{f�1t�5��������@oP/,@�agZ>XZj��,�#����7��M<w�"��`(���S�H)s$�P9X?:q�
%L��%5�u%}��l��
�J�2���[�Ʒ�F�
��(��e��N��u��Y����O/��~��,~�)%�F�����|�T2�Z0r<@�u�Fٶ�<4��⺒��)	0# tF�q��å���XtT�M殏���v��z�Kung�� ΂������Rm��s�?���=*͜��$(�#�7��C�JG��#���Y�E�FJ�
B�zp�7�6�%;Ƅ^��(��3�yn�Xk��-E�:�d^�B\���g��v�
4�pO��$:�rJ�P3ԭH���Y-P*��Rե�����C��n�qT�g=-G�g��?�LH�g�(wR�'U!�¼��+L���?�h��b/K�S��a_Q�d}?�NY��`����E�T H�:P��U������WG��-�]ܔ���::[3�Fg���?T��%)[Pւ|��JW��O���*�E���޸\9��ޓ�B���o��r��J�+�*�P�6������Ka'o��e���J�j�sA��o�0벷��A��釈�yc�p,�V�/jF�[Na���̚5 4�(��`������7��d���J1@� ��އ���#��:6sx�'둆Co�rI���	r�43@v���!�x�Q���Y�<�n����X5&CR��R�������Ml��kw�k��g��