��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~,�[�������i�g���RѮ��]���nS�ʩ��b2s�ٜ�����Å@�r�G ^���8u^I�0Zd{ߏc��s}Z�౾?�9}�)Y�����C��T�����g�x����2T}�5��P0���ɟl%3�gV#�,hJzpX���e��;Q�kt����ـ���lM�	N��:m�TS/��w2����]?v"P7�|�$׹zץ1u�"����C��oZ8QC3��F��!U<���5�`�s�Cd;ZP���rNNLfjY00Lw�y��ޗ9'Jqw�߉�v<�|]�?8�
��$fz�ڌ\�.�y
[�ҟ�u�N�{51
w�py���J
$�\u����y`^魦�� � F0�����YN��\d	J��"e������Ǻrל�#���o�����~X�����{�I@��d_�bJ�͊,�6�]�Gۀ�Svu� H�Q4��;!謱$cw�"��hp#F3�����#�F�\��[�e��a���\�BCa����_{I֏��7=�4Dŉ��y/`MY�>�}�hi��|ر�X��߉�rI�@E��n����4��y��ti�c���^����6��n?��E2�����,��"ʅ��x��`�J7 #DЈ��у�A#�ɔ���wn�	��/6:��9��mw�d��]��j���꓉&��|�'���'���� ��}�A2�qӋ3����c�r}���w��fyc2���������4n�fI�����|mM�Y�����c��!<3ou��e�0e��.\8��QI���=�a��S�|����h��4!]��(��/�D��[t��y͏ds�]IIk��]��4�����O�6��)�e������������+w�CY>Fe�cMT��&#����r�$bZK��Y�Fd�ꑡH�?Ql��B�lG
�V�b�E�4�EoL�8
\�@��d�x�+�	H�	�D�Kf&�q��eU��
B-`�.��ӉoG"�j��Y��B�B8�C���G���S̀����
��%a������K�79�-@��S�f���a���������Fg�O�1���ԋ�٣�/6C��G�1M�'�9�Ǆ��K�:i�������%�)�`]�Y��4+ŕ�U��}(���3�"�Tsȫ��{��&�Du��Ѿ9ϸ�3E��e��!ԋ�oש)l���u(� n�
�:�A+�E��>�ef��ڑ��gnC���HP�<0F��^�T��qY�N���^c�����bEӐ��ˎY��m1�����R�2���?�y��jS�Az�S��mi~�\���eGfY�����M�b��>|�*��90}�Õ�{ϥ�I���M��c�`Ĝ�@�	l���[�b�N�|jWls�p���[U��@����cBu��hfj�}}_C}0��6ݪ{^�wX5��zpdL`�n��;ZO��8���e����q�V8��T������\�?η=����U���!Fq��T9;�gxBgt����7r�R�#��t�f��n�eZ5g�(��̞rK2V����?(��t/9M���x�<��G��۸w6�X���o_��8���}�������s����@��X�9yD�WJ̹m���P(���
� �>㎒5���7*��dڤGau�&U?ӟ뗔��}�{"����O߶�W$�	v�c铇���ᐍ�7؄�]f��?a�H�����h�x�G����0+��b@gA�y`T���<=߃�@���*�"��o�邓�ac����|�A����fP�����.Y;�,w�gҗ�tO�{u�$$WD�l<��)Zo�����yW=����AR�`�Fh Ϟ̜��dְ'μX�8�!��:
+ASZJ�ԍ���Ո� �3b2|DhH*g� �����Pnn�4���3Õ �Or���fz�F�b���2�{Z�%P�(�wN�o�"J�L���E�i��&�`�OQ�]$nƱȸ��N~ԯ�r�T��% v�gE��˅�]Cu�C�6�j�A�!5�0]v�M��ߴ��ƓC�r�G��]��S�s4u2�h]�Z��S������q�&K1B�p�$�[�h�L�3m[!���=f���Yt�ԂMɄ����?j�o�a�������MW��x�O�|�D�
�����ǐ����K��?g~ȪN1}��m;V�|Or��i)	\����nR�18�D!z�Kf��RSכu�� �˕�V����&���/�ޜ��gP�yԯ�P���	®�k��$�@�O㨒�Zj�xP1c#� b�����QR�;�~��9�ѐ0��,e��.��5�)�~1���,��rQ'uy9�(нXjt��;I�vP�g�����ɬ� ����[͟cԣ��*��6l)1�WB�H���� n��4�;r?<g��h/�if�ҥI��baݴ�^�q~Kb��d�&d�xy�oO^���ʟ�5��V#�u���FC��7"�Gܓ���3qL�%����W�B� b)O�Ͱx�xq�Z^�Ma�`n�_�m�+�?n��\rL4��YG1D�Z�S^)������;e&M�j�0�4��~)�Oi�3�na
|��
��f����-�~$�4�[.�� 7�}bh|��������*o���b��t�r���-£[k2p��S81�l�(ފ����Q��~�D�sU85��aش�'"z�"��M�|Rx��ö`m�-�;��xTP�r��?3;ؗ"���=���|���-���� �\��&��VN3����� ��\�uCG�E�I8���V6>�Fly� ������,������H�\U6w#����T?��ZU;a���E�Я�gP��ߢ�c�w!N{<rԌO�ȡ������$56�����/`'�ό)(L���ˬ7.�XW�+A��;�gV����H��1̢��nvF>���m{�"�g��'�jW9 /��쟙3��%{�?Y�4��E���ґ��^A�>/����4�`�ql�܉	|�b�u��hM��g�|����Ŗ�.s�w^��p���5M���i�
�b�(!�̶&)qw������ �\��W��Ґ؏#������ّ+�j��Z,��̹ˮ3�!q�!�g��c�]ʎ�M2k�.�2���m�Yw�Y�,��)�,�M&��(5Q0'Ѹ��j�w�%��Q?cU�f�q�<���s�l����,-�����X@_�:$���T���^���XI?SI������J��d�J6��3I2��U�}��0�w��wY��������2������6u���@���[u�!29��, �S�Mm�Ȭ���c3�:���~;>~H[�u��ͺ�@����y1!�љh%��~�0C��K&�k\O��J@����s#��ݛ�����S<�E�b��(�N����ݧ]���0[cb/�\`/\��ĉ���NJ��bN[�]/�����B��͉�J���U$S��*T7���Cb8��n$t�:�Qp�G���	)t�5������LQ���_^����o ���1���1���wv���;U�Y$"��sX��[?����
3k'g���'���i���m�֮���oA�J�HA�R�qÍ�I%���^=N<Fb�V)��O���s�,�v�ۉ�v��-w2O"�r�3�&Y���Qz;y(��\�=�eh��F����F�6G��A.��.Y�&� h��>����9�7�	�pVF�}�3���E��mE��Ƒ
�z�����SP(��~����F�p>�/9���D.�>�G����� �i�6�q2_�7��T΀�pw'@Ct���<!)/�"�+���aY��5R��p+��WK߀xģHR�vU��y�K���r��s�nn|���(����"�N:c
!P	�ǵ�����Z���yk����j��� 3񞡊kQ �@�5�#:�<Pag���c���$+���H<
�����Ԭ��� X�����27H�j�2F���!'���!�¦Vɟ��β0-G�V���j@��٨������~�T)�;X|�,*]H���^�@�.&��7����p3��:���?\I�� b8 |��'fGK6xP����Pr����tH��w�.�k8G+��W����񇩷yj�힒�P$x>ַ�!Q�,��dǢ<7�yF�ck���P��z��O�aQ/�Rq���u?��n�B�X�>�xS����w�[�������I�}�ZZWO���JM\���if����w�<Ԑ�CR�"*�j#�!
�#e�
(��M���6���W���ޟ�#T������j�,�Xг�����H�����]��,T>�z����N�C� EJ��O5sII6$����h���^��!�!���L|�)'-���-B��K�7e��0E�7<��.�$��N�هѤ�
�!:N)������#,�� ��?�y؝��c/��l��(��(�ϐ�v��=n�	�	�4[Kpv�	��'���:r��HK�c����^�Bn>^ֈQ>���芔K������ a �ISj��}�I�/�(ch�$�.(�L%?~�^�2<��Ltw���TxE���Ԍ!�Y�v�/Ӧ��ʸj��꯮in?r���RȦ�4���/��h(��ө���6�����`}2��h4���'s���
�d�խ'�������ʵ�=�!.=���u��)�mV��π��������W��%�#QP& %2?>�ACA�y@o�2m!�'��g��"�q���\|�W%Qbs�m�}o jJ��2�)7NZ�Z��jwi#�J_�R����*�<��3��E�T�ud�D�3ad�x_�kq�>�&����Dӝ�a�)U��|�>Ԫn)�q�g��e�11�ս��oT�{@�
��Yg7,vw*�N[�3���E���;���)_��q���lqջ6�-�I��4�8�9[!��8��m-1 �Ew_�f4C�]G���$����)�>;�^��h�V���R� 1�3�#���P����!J*�?��M_�$$��Mz"�~�y P�;AP���B���Gvsℼf��B�}kW�z����C�[���82L��]�����=���u[Q�z/厝N1e�9�e7�z������ �*n]� ����Gģ��3�Z�8&D�ͪ�bՑ�w�o4#��_٠[q#3�+���N�E�Gì܌0��Op�_v�G&�b~���a�Cȕ	�l =P��Y��G���h��h�Z���]x��V�l9��;��d_ 3��;�)�Z�_���׉=���ۻ���~K���b��ִg����#��j��'�z�1���%��^�p}_�E.���͒��G��fy��Z&�b�eL*����8�2��iv*҆�f@�n���*� y�Ʃ��nG�F{ߞ�>�y��� �t��/\�kښW��jj*[	@4Qe�0��=R���q�Xi����n<��ah�+v�M	�Ϫ����j��������@�j�s �T��r��K��l&��3H���8M{}�R�F�gR�����ba�豴�����3P�p����o%.����(CNH/��o����v)'���0��?�N���,[��C�J�wѩKR��̐-.��t�� �h��cZ���K��m��ym��^2��*&����_G�B+ۆJ����=ᔐ97��F�#X!\(ť���@��`G63��J�1�b���⃄�g��`~��,�Z���O���-l�x�~'6��U{ݮ����F$�^�VDb�0���8@}�	q�:�(z#�������_�g���;��z�$�?���JHb��݆�[��F��2=,��Xw/�9<����3��Ǯ��*�;9��A|�\]�ԕ�� �@����6@��/ 	)�.X��C���.����fY�]��˻�;��kk�r�`P���6$ɚ��� I��?�E2�n��«��V�l���g�.�_T�n3
:�� ���L1�}�"��	in[�`JU��0]-�sU�T��R��Ȃ�����51qL���MRWҒ�:4Ok���f�.�%|�s\�@�X3��Q�=�a̖�|Q�NnW>Ѱ;�ٚn9����*mŅ�5�[�O�嚭����� e�T)rv������q2 ���l۰N	���a@ �e�%��hP��I'�<+�F�q ?�!��{��o2~/�a��h�Co?�S�r&C�w�6�}5V��H�����8���X�@Xϒ3b�U(�N$��(t�c~GK�������6�0�~�j��]\�J�Y�u�>�����A}{�n3?�s!c{���/x�Ng��Q����^Б��7(��a@��4ԉ)6������<>+YN
z�o�F���W���ze�~��o�U^C&���5t��8�wL����3R[��4�-�ki�aQ��j��%1�ś�F��Zc��.l�V;7��S��*�-Kk�Ηb��J��l�GF1v;�;a�F#`�"�"~���BJ�ѻ%��@�&����;`�R��b�+p��'&�O���-�Q�ec���a�S���࿷�5�ř��<��mcU[�jz�p@y�ƟZ� ��'(����� �"�R;����P�f��0OO��aN`�Y������G/S�H�J�1���I]�+�Щ*sf(:����ҡ����Q^xd�[hR��șɊS=�u�:�mܚY84^u��[���H��u�f;�V����a9$L��3վSԁ$l��r9eJ�r��+��)@0��#�ӟg��zP0�T�6Q��D��.��"�pT�v��q:�$b�N kх�壨"30����d��*T��j���K����.��	��D�z�L�>�9���h���? z�4�d���U@c�T��3����������T��G�\���E�O��wE]7�y�Pe}���O�J��<�lQ��83UAdSu�Qmz%��]�\��X�����ywo��-c�<�N²�B���?�ۢ,S����!5B�ȜN^e�M5�~#dPH��5=��an�]�c=����kol���1W�N(0�&��f�D���8�-����اڬ�O�_�a�7o�*�]����P���:�I�s���N���ÈQT�߾����s[�~�8�1D��Xm������h}�35�{ԑ̵]Ƿ=�P�#.�!1�����&x �ZeG:�l����sP�5��0o�e�q����$sR�M��Ӂ�\�a��0RD��E���?1h"�� +��$C���!�`g��D��
�F#����pj���s�.�_��Bm	�
��*:!�6m������+ij���s���=o�A�� �c6�1SN�޹+GNA��_�,	P�~��n�a}�M� �ц�Ȳ�:)}8VV�X���yi��lm�'� �b����4�|��؈/�}4�"8"��r�D��m�	�r���+?�:��J� p�9}�4d����*�f��r��Mݴ�H$��@�bְ�3I����nNJ����j'�'-�go�F�~Wg+�f�;��E�AX!ם�D�k�l�Г+�>��]��_��,����� �s9������2P�5/g۳�T�\|amjz@�&b��i٤�{�R)���4v7��v��~k�?G��.�=�1W�6P ���?�<'��?�_o�}�Rw�3:�B$;o`����|�C��I��6��(p	% V=d�B�-��U�^>���F��cd݁Lď= P�����	h������G 
"OJ�_�7�O���խMA���t�fI�;u��\(l���#I]L�z[*`v1������>d3^�Q:f���r`.�9hb�5������������$%"T� dqO�融����J���o�ԙ�Z"p���!�\��ԩ��O�T��<Wj����)��Aܰ��D��(T/LZJ�1
���BD�M���f43�~Nc�L����ed�7����}[�!�
o�2cPd�x��1���<�*�S���ؐj��oR��<�t�)*��T�'�=���/�m����e�xr�P��̏o�৶�e&����=,^�q�#�4e��L�Y��D�"���Bt �K�O��Mk����
L��a}k�9��dx��≒���qd�&�S��|�w�H�aig1<w/�ף��M����כ.������=�U�ND�a��'z��q:�S�@�PKWd�2�A�-�ЋU�ɂ����v��3(�1R���'��5R���$%�Kg�8T4~�H(���|����X,2P���>����>��H���&7v�^�������W
l,k��yk�`ޓ�IU�y1Ȍ_����i����In�㈼����BJ���nr�/r�2��5cG��n]Dw��$�PT%t_�mr6��K����,4j��w��j�����L�2��u�<��}�ڭ�L�9�,p�T���^_�#-�%�5G*	�E����{�C��Ն@�
B������鐸|Q}����e[>8A�e7$�9鰹}���bY��|�	��Q����%�������oB�b'͋u�+RF���m@N2f><
�<kSQ8�;�g{��H�G'�̿j���k7o�0�eݞ�{�Q��
W�X�/�2��׫�7�;?�<��W�h�C�����H�͈�C��MV��A�ǝ����}��99 �;q���z��>��Ūb�_�`���*�(ɲ����@�Z�ytq��}���%�I]�ҊK�I_����9�:���<�\��&�Dd�ZK�!���3�E�S�EI��B���T!�>�?���r�=J6˟�.��ܸ����Dwm��fO�:ʤ=�9�� J��o%��A��P�:>ˣ�A ��"���~��I���~ �N\gG��o�mf�3��fc�������fS�[S���e��� �@���<�{������#�v�7������;L�BMN�L�;3��u�0�R�`�p.�F��;Ǐ\>8)�,�I�U~�����n�)�2�*a��6��݁`��_-�W��n�A�ʄ� O玑��i���z����EK�Myc�"#���_�{LF�t�K�d�������/ٴUm戰Pk�I��`b���Cd�?��,cOӞ˖k�-�]n2�VL��l��m�͊�ww�V��-�v2�$��h�[��Gc�g���K���p��v��'H����X ��C"/Zƃ�p��'�ӌD���g�TI��I2��6�����!w����F��ks]�#�ߤ�p���=٘�$k��nЍH{4O������Ffc�Ҙ+�ơRN/��$%;�-�0���֣�=LX{�FV��DSb�r�ɉ�]�^�W����E�<�;= 4���}���x�}oYĦؼ	a|{M��@��� �0�Z^�a������<��'���/�@�0kU0�X��6��	"2Ō
ΪӇ��R+uY�<�4wL��?��b�_{z=$����լ�7�Q��۷��j�Պ.��S��/�u���3<����	�`�)�ւ��1_�c��W͞��@U=�Z��)gr;��=͊�yPW�:�_QB6�H
'~�WF�
�i�Y�|����X�SFm%�},B����z��}V�#��W��y�:w�o
/���^6�B��\>F��s-6]'߾�@��5�4�6��yy>��𣆆ʋ$�f�������F>�B��
�* 4NF���ꪊ�t�pW)B�"Yq���Sb-�Ҁ5�g�onN7ӜJ[|Rݥ�«Q�n�e�I�tL��l��n�g��EP�v��������3��$��w̛QJy�X�~�t�-#zC���S�� ue�	R�,z�9�Y�8W�`LX����V�g���ٴʹg��%���R�vH�@�)@��y�4���NY�p9�Je)8d�/8Q�}��c(�@�vr�.���������˪W�Z[��$5����؝�Û�>��n2Gh�2$c�0&KP%\Ŀ�;�y���,�����l�;����V"�e��ߙ�(ߤ�L���Cʑ����M����7Gr}�C�B2�@7��U�`S�:� .zE�9�Qڜ�4ż��SKqe4���Q��h�'M�+������N"����3o��>��Ź/(�����Q�`G�S��eXA�~Q��԰S���'^�_7�եD��~�(O2)t�:z�sH2�{mwN)X����&��M�ɸ#P��e&,�#�dX�t�YS���n�5'�\ �ŷ����m�`WE4z�)zU����/<=Bk��t\�x���^O������J`�-�3E�����|2T�2!�Hߜ�=�P��������i.�1?�ݬ��Wj���N)���i���8�5��lAǁ��b`&��R����s$/Sx�8Lf��~����+����x- =Q�}��!h��R,����'B��mhi��xf2�^�u�t���}7+Q�;k����DC�T�Pqy�/�� {����������U���yO�~o{`R�$�޳n�Y�uu䶨� ��ɼş�r
�gT�;��GI�5ֲ�(�E�Ьd�m�s��h���&��ݺ	�7}����3�h_�������ØG9�*D�/z�m�j����P��uLe�-DI�H��ؓ�-����=����,(�����([8GJk�p~v@�����Aط1F������`B�� �=1�L���
H�5���ǓK�!���Fi��J��uNj���xa��a�NH�+�z�a/��H%��60�g��+XI�E�� �"���֖�'"���������ۇ�4FO����r����^=ZhnK ��� ��h���,kԠM�}f&�|� xOi/���_a��qZYJ��'[�;MC(���������
���h�~�b���h9\w������I#��;:K��t���8����7���>0z+FBX8���?�`��bed�r�8��Э�)����0��8��@�+����3�+�[���pZc{�������}�H������y@4�*d�2� �9`��@�G�e��ձ�&�h~"��y~�f/ߔ�D���z�q� �J�����D�!��5��G.�FW�1�7�J�HCK��x�W�fJ/#�e�p�Q�w!��B�ՙH��!��,Al��
��J��wRJ�l$؊��u�d�u�'3Ǚnw6��3G?<C�Kؑf\�! ER��mpSv���l��Ҝ��<<�L �tm�(L�Z�ˬ �}����XN�nQ����P�0c�FX����X]�@�Pz�!H2`%earg`e~0[��@=.�a��,&���[6<b�2��JeG�=���jUϡ���6)��ȍ�n<.�������R�1>���C��,�Ȳ��4�m�"���P��y�Dk�_;���㳋z�("	H�W�DWş
�.=�^�]7���i�C�}c�6�,\�._Ӗ�]<���s�b�7�����N\��hР�U�'��4]) H��o���W�j_e�r����ߕ�����~ߑ9�d�۔�:�P#�O Q>�Vo�V������%4N�
�.C~�
�
U�^��lu���Z��]�ff�5D�7a��tB��~N���	Xd����]���=a� �����^��׾`���+b9o���	�ڃ%� 6# >D�}^���~(#[�HSb>}$ޛ�X��x1�y*��뙨�����W��D��dd<Y�]$�����.�k݊D�w��_}\Ȟ��ޝq�k��N&�4�0ȕH������u]��VX�aɫ�n�b�SlS������4�Մ$n>_����:B��'�I�(h=�)��T���.��Z�P�#�����Ϊ�2C���K�����8��s�յk6ʩ� ��)Dpc��pDV}�n�7B` w�df5�Q�s%�D�5O�t4�K�0�m�I0%����r��ƙ�[����9H�ǃ�Z��d}��b���<��T���r���� vr�`eF):��{���K��T�uʤ�6Zף�Y��˱���?��nv%1��*E���K��t��P�_��2bq��R��Ei؂ ���2I8�j����j�&=Na��-c����;}��j�D�:���H#�|�	Y�mM��Nݑ���d-�e5$I�����B�5��c(}��*,��ai��M��!�`(�ϨZI��s7ޜeecWT��b��TI�dG��uDW-���R���w҄���ڎ����2&���-�� �6���RT:�SS����,�4_"kfaZ(�՞-�I1�XfKC��2G���3�P��(���d�W�á7FE�:��7`L�=F�qˢ����N��RuQ(����a�� �s�֝����,�15S�rq[��o���f΄�u��l
#���mڧ�}��U�"���@0|��
=:�aH &z��X+�~"[b��]5���p�,�u�F��5�Ȝ��aM�X����U�A(��Ӗ0L�F�ၛ$E�����߈C�Ch��- ����Iij��I*���#�>P%���;�b*��P�Z���1u�A�s���i�F8��9�k!�!d�a�ў�I�攗���_~7�-+�$��>�2��p�	��q�IAA���x*S�'5����� �.I(���aC��ĕ���G?�j�m�w�ޞ�B�Άf���ޱ��������c��[���!p�+��wL��{���q�dXv�.o��w
�|��T+��~r�#[E����Z9\B�����`|�����=�ڱ.��:~nF�)Y+�/��� �9({ݧ�cc'9�[��o� �ո���C�d<>y�}WB�u6`�
���*�N���"R�J�|�C����d#I|�L�5R��F��.�t�������6m�*.�i�(��B��>p�V 7�?���yGfF���E���T�]�a�b�Rc)��𾖜��s*=�B�v�J4rm K�d���B��Ϋ_��;���|��;��S[�L���~�ڬw䡬&S}��c�$X���
}�sj9(��e�z���k0��n��Do�[�u����ub��V?@ѻ�`}a��B����]U,���j���{y��������r�����`^���EXٖh19xK��#iK`o�� �~A�蜳�b%���t+��f��p��˯N!K��p#? ~h��m�t���~�9��;4W�A�P��I�L������9 ���Y�?'q��r�t��k2���H�<��}]��}a߽o��n�T;$9�r6�Km�;#d���P���A�I�*�34d�*O}ء(W�%�L�rĵc�c? c�H�lo/ٰK��:Fu{�`���6�$^|F�+�:56�u��Jw������2f����)��<H��\���B^��ۈ���8���A��{�_�_W���ɗ`3����.d���@q1��]k�A���-,���=�hQJ-s̺�x��MBT�* ���Q�� n�v��H��K�i�%۫M�v7���`k}i'l�X�H� [�H��N����� ��%��nOWF`���}-�+#�Am���^�,��0�(���+X�Q�'���h.��B
����r�^HX�;A,5��������fBb�n����-��˿�,g��9���l��fk=}]�D=�x����2l�F(�ۓT�i�t����n�k�
�HI#�`R�v+����ٻE�j�J��g�U�7QD?3%u:p/��WN���y�����T~+>J���&:'MgS����ʈ�:6,2dO��w��<1�n�Lw�u0�&�G��.&��A�M2���N9W(�u�3�#�]͵��nrzi�}������h���ԶsFw��9(���E�3��L��'����ʸĴ�����;��چ��;�7�%����_f�m�2��q����H�"	���&��[Y��#t���IV��nne�1�\7W�q�j��sO��߳��T� �]K�."l���>�G`H�1��E4��F ��z��l�'25a^��k��lԊ�����n���d=�88�n`�\p��#w��o?CH�b��B�T�@kd�\$�N��E����G�o �A��^O��%6j�R��UТ�Ii-C3��[h��8P�'ڒ�:���./[Z3m�vi���<!41YB��
�0D&Hf��0�G|QY��H���N�\B�5REk[�h�c [q*��c��ZΣ�?p��d�:f�p�]=yT�0��纉�l�7p����<S�Zm4����C�
���|,����N_�D#���讅3|e)��YG�+�-����|�?U6ٷ�h~H��<��'�+-���m��l�(Ww�w�eK��ow�	T/0���Kt`{R�����Ϟ�����U���C�G��(�XW��p ~"/�� k�8p�iDp��̼w���XS�"P���`Y���5
h�{��~iE���˪� �]F��]T�|,�����3�B�R�r�q��U��j�:��L&�8&_x��:�*���4��W^��jVBǖՄ1���#��ol;@Q'��g���ݭ֠)뮻�g�(we�S)J5���j����{|̪��m�M��;H����B��V���Y�T��d���9�A>�w�,��@����sk ���V���e&Q��Ʊ�:A����{&�ٰ���Yi%�Q�EwXA5�� ���8�����#j��'��O���줽
���Ā/{�6�Q��r/�4 �s�i���~�n�c)�)�>5��^]Z��%q����kZ������1��u
ψ_�Xe�U�	Z����G�_���Y�m�e���^��_jQ*�?�aU��hZ�3���u �%W�0�͙��`՟��_פ�`�'�-�g~�R�҆��Iڕ��=a�h�q�6�sei��s�1?O�(>��/90��b�� &��%>�ZBx�Q����}���������SI#�+D��N��$x�������a��.���m��O�b/�Q�"H��V�{��t�s�<p��c[g�A�P�ޑ��@�$#��=���d�����x�[�� �zV�����-r��&�������i����S��loo
Hes:�J����i}"	�*����+��x�%�mQW�a���R�6*�3$�h�#�j���T���X��²N���j?���U�{jU�+���k���_8ei >�1�����U��LN�`i0N��2PliB�mu7���0��UR�w���%����Revv�%Rg���~��|}%�+���w�)�	R���'}��֬��3�q�߮k1Q+/ǼfC��}�jz%�Y�*��q}TG��I
?���	�����y�a���M� ��r��{��M��1^�uC���t+�V��8[�O6�1m�1V����KJP�!�)�XҨ�0À�He��n��.��l�N"��}�v�����<]w�҆�/r<?��1���c]��0�t~e����e�q�d:p���V}[Y���0��A���g\H8�Xc6@�R���f�H)���YZ���z��\��g-9qX�͆��u��������lS���xy/�i�U�⠣�άtJ�"U_#'C��S��'�,F��[���fSBC`<�ΰ���`��pNÖ?�� 'q�T�  �}��?
����-�Y�P�������OA��I�6)�����$��]5�����<>�GU�Pמ��m�?p�e�YQ}f� nYw��+(wp_BE�S����#8%�c��?�qI����̜ �^��a�p�����L-�u�=# ������ڎ+e~���R��&RF�k�tX|�Jb��\�o�ʝ��4�ԌH���'������h ���"a��߷��Ä�1�N�����b�&���[���i8�yE4��p�����=g4�� x�2Q�s����Ĥ�[�4%'�����"#m���;�j�Q"���t�+�#��~�s�Y�~�����L)c{�pݐ!b�[�X�D�	�w���<=Pa��í�5���� ���d�9j�χK��m�_,r�+a�2���_����ߌ3��Jo[()׾B�/[���Η�PM�xi�o,>���kyee��ץc>��MB,8ʒ*�A�ʎ"��)�&��e�&�B�^���'55���(I����?���ܺ;6j���iZ�����)%�J.�űX�����،�77�?� ��v9{45��v��Ȇf��>�(hV'��4�^n�ٮ�u�������oa�hY;OI��z!����}@���;��R\5S��ȫ��/���-�/��R@�����E�B���h꣘�[���_I���� ��=]�"5�T�U��M���$N V�F��0�~����<}'D���O�����]��4Ӧ+e��/G�A�)�Û(�GjGb�F�Ӎ{+�>Q:$� .){���\cXq>��F�v{,�k7o�Y�xT}H���թPs��k{�&�ʬ�!��4��
��`����0�	����a�$3s���
1�5��k��d��j�S�H;/�2����T*��1��귌HAY��j�~�+PXa���Fe�꙳#%�
�w096���M��C�����6��\)i�Z�:^�}�/ ��{mg�_�=��2k���\60n֖���Q�F�[��i���{ P����(F�^��@�K��k�"Z�&�-��~f]a3�Aw���|��p �}ԈY���z���[i��Њ�շAO�:���39���0e��uG����R�����^��ʯf�H������Q[��	�	�(�^�lj_�H4t�ͮ�])�m��~,����=���p&'}��:0{�������-v����r{K����R�k�eB��� n��K`��N���'�>��r�nl:o���7�3͎a��z���z2H(��T��}�±���E��;��F����>�tZ�+(�ܪ���/�zf��A
�=�p�:�
�fiH�ݷ�đ���.F�������B�w�����t�$&E<�܉��E���;z��k�v��E.�	��~,�Tm�QZͦ� dS���x�õQU�2�}w���+�X~�o˝+���/���O����b�{�;�R �Ԙ2G�(<�}�Vg��u�����C�^����m��6�w����1\��ly$���*�saq<���5Νv�� �H��P�P~�q�M����!ͯ��)��e����7�>�,A~jS��F�����k����/wb�sx����?��pO���m5qDr�r �]Q�?��@lc<��;Kg,�������ٻ���L�����EL�Ҽ���K-�����/����5�ƻ��6����-т���m`܇1`����6�`�X�5�h���=�>b���g�:��ݻ
���?�1q��/U�~�ҿ�Y�2a��\��>+l'd�G�Nn���s���~��P�B�w����Ò�lMM�Q��Ì(�-#�՚�{|q�E%�X4 2O;A���
����#��V6�a.��K�17��ei�ψ�c�*IX�L�GGeA�>���d��������!��w�M	|8G�ظ�S�����*YF=A�����Mh�|�f�F��cHX�<#�0���Q�2� 3Ӝ�+Yξ�J�?!PHWIh�ڸ?� �l^b��㴕#��6�(OV�j�BvD� W�M�V��u�/�zLU�n@5R��VW�8`��M�a<�gJ��z��gu��lЍ��s�OZ�*��_n��<�����:�\ONi�1�A��q������5�B��4�e(��i����W�o��A3�Ur�^�73?K��5J �߄&-3����t�^^�ʴ���jH45���,8ظ�K����׀��U@�h��`<�J<�F�ؑ<E(]�w�d4�bE�s�Pq�%��wJ��D���B����O�,S,���+�uS����ArtE��j�+�u��k�{A�����e���k��l�^�����
��È�q�}�7��xR��Y22�?���\*��a��c��&�j�^4�^R�&�����w�ajaMA��s��Z�~�%D�|�6�ct��ĤU ����G�8�^��^H]��lM"o�X���#]J<� ~<��?���^�vOD����}���:�q��'����9��;e�toP�#���9��l�8��)�.&ɛEOyV�s��$)�ᙾk���r·̕��I{��\`���*TO�Ӆ����.��sl�4����� �o+���>6E�x����W>�R\�;���3h���<��Eu��ݙ�L2�G\ /�� ��`w�ed��k8�@�$������R93_�6ۏ&�{�u������4�ȓ�(�Q#�<����չϝ�M�#n��[�i���x/��NN�t�7�W�)C���i�%*٢�ĒDϝ��w1�K����Vl�?�`����ov�TC��OxK�&�!�C3|mJ
(��R��:Oƀ�Mȓ*#��g�Y�]�"�fu����[zI}`O� �z5�X� /r��`���?m
K��J �Jt�Y8�g��u�e�윗��#M�1�L��X56��`�fZ�{��Lv��[5���)�d迧n���>+�٤[R8��@�c2��m��W;�qb�����4�Jĉey
S%	��p��؃T�\�]3���`pB��|J������:Xf��9�L����Th*�}�u��_����r��h��N%KzY׊�Թ纳55��o���R��M�zL�h�GH���k��t�5@�2��#~� z�/���1�3c#N�ho>c�MN���j�EG�x ���%�>�#vE�W�o�L��v��5,Q���Wy�.��-K�Ӂ`���\HҫD������ ���H4�%�Ooм`a��D�~��1���ag��C�C\9=��O+��9�`f��u����8�c�	q>��9S�d�ك V� '*e�À�W$ ��~J��	�U�^���p$}�Z }��ѝTsOukC�h�1�n.��<k���~��bt� ��<�Kq��Q�ö)�J|w�����cp�.���XM�L�*s鱯��?!��קŨ��[#� Lrq�
T�I�=f��p����:I�@�ǀ�#���H?�c�����n�HjgU���S���v��Ғ"Cs<n����|17fv��lD���TM�'W{���3���n���w���º�Odp�5l��/��iz��)��l�N�g~:84������)�'{���x��<���{�D��������isq�򌪋�Ho7�����l��n�e�9�5+D���3���*����Y����
�c�����0���|d/�� �L�xR�rUZ��t���	���7� �<9����&�؀=v55���h` �ݱ��T)��Ӳb��΂��(DA��f=�+x+|��h�~Y�D��#���U��`.�$pO��J�#�m[LP&���&����46ݬ�1��*}uV�¸����ĎxN?�ι���j�6xj�)�_��$wm(��6�bN"l,���q�.��	66�*�-R�G{ 1�(�r�j�2����U���_J髐Z(���!�1\�+�e�F?��/XR$������>�^�]�l�<�2�m���=���e���Sp0���)����}�x�8�Ή�������Ѱ3��^W��Ib����z�L��v��W�Ɯ�'e�@��t�=ŋ������ےC���В�55��7Z���������u�(�Eb��u����o�64Iw9y���U��K[���:xD�ݐ6��?:y�JXaZ��NF��\gx�R����J2�?3wwCA ��[�;����.g�DӢ�˨>�=]4{�ؼ�C,�w��
�(n�gp:����c<��vdQ�����V%�����0��j&^G�Z%��g��;�ZL- ����	�B�j� k��ӏ�O
W����׬ ��A\&�7]6��DE��z�'_�sa���*�6��_˿�t���nعA�B�c�$���Q�͊'5�ɒ���b�;��*Ҫ�BC�^7�����	�2���5��sZ.]U�X>�t�P�=4�}��n�_9�m��[g�oj�ݣ�!g��W7� L�_[O�9X�f���k.��~Wh����$����i���峐t5_�eq���*>�M�\��d��5��:<�l�?�s*���4�2\�U�u�T�zE����z"o𤄙ٻ8�=�X�&�-u�_CK/���?j���Y���G���P�Y�??X���C�S꿪tFk��~0�<�` �|��ޜja�i���=�$]]r�{�ޡ�%�2x��������n�吂�bI���WKh�D�5cr�5A�����p�2 ��_��v·+���"Kf/fZ��z�A޺ J�C�H�b��"{jd�e b;�K#��$��
�/Ø8�ԍCU]�H����l?���\��[���J@�Љ�� ���_k�6>v�Xhȶ��"X	�I�N1IX//t:H���(��<�Y=F��ߩ^"UvV���n�jN��OpF��h�tu�J��N'길o����ُ�-�4�č�SG�7��y��] ����yJ�d=��]��C����9��2Ч��r�_I���Qjb#��
��;ڕ�ʶ9붓j$�/�1I�%��Xמ@���X@6���K��ya�f1��	���r�O=	w���X`J��B�^�FA(��<��d��Ù�4�UIu"CE��A'��{
�����]'"��R���n�j4���]%�vy��2�\yi��[G�V�h�_whv�l{K�

�:��ΎU��Eq�Og`��s)�v��cv�:�w
����"'���Y"�	υJd���~/�#&e�D�7?j�ޒ��~��JE��9��ѹ!�2�CS�v� ��E�}z6 }1�B��p�;��u$f5�s���o��ZsnVֿ"}6y�S�c�~񨴹4~�3mVJ�A��U�}�s��kH���'�]���y�]���Ψ�Pb��G! H���8������ޅ��J�1FW�p7�+܀f��r!XF|���wM#�²�܁�+GS�iS�w��ғ���S�P���훒��WVq���S���A�o]@�����V���T���̑Fh��A��I�,Y`lz�1n!j?z�%�5m�����k>�,�E�[�jMk�bZgo�5/�;=�����i�}�ӱ4Ҡ�ͣ;���׻���i�%�4��ak��\9`k�@c�Ԅ�
j01�K�C��ݤ\�����YC�Ő`S���om��iJ�&(0q0^����n��f�R�G�~A/Zו6Ӳ-;.�6iBo��No� ���͓�ǈ�-떬@��]Og>����P�]3ݪ]u%��zI���>����d6m)e������]x�z_{a�S��Br�bWuoZ����;j-$�.W��9��ո��r��@`��v�@��dACL���a������ �$��"Z�ئ@8pd0Q��a0T���:8��~���P���,�v����(�Ĩ��gjNs����w���� ��	��뾼��!�ǂ�^�[*��x5���s2_h��b�fT_������:i۠Tq�\�������+�tuup�I���mI��z���%����L^�+���:s$>���F��m���7l�k̚:�T�˝�BOQªx/o�]n����q4���6�1��ZDx�P�I�4=wc<��R�o߅;ĸPG�Nݐ�(��g��Dh���$~
��E�$ �)l�u9��k����^��v{p;����QC�
��!/�'����:0��3t9�W4'}N�~��\lx~�G��m�����#'���&���1_y��)�*X���j�2x�0�PT(f��t���:��
ϳ��r�t�5�F ��y�_m��k&�`���;PhLc��_��W���s�πы���Fc�5#���J161u�=BM�@.��Ai����&�`�C��E�$.�j[S ����cQ���[��oi����/�4�0��jYd-/?���*餄!�S�:'��We�x�E����30�E�L�*�8ڍ�a�"́��JA%�@�!#u�ϱ/X�x.h�L�@�`���  �l���>R`<c�X����ã�5���7�/�+��O ���.n��ү¶	V^��{�b'{����|����qLK����m�(a������4��i�֋`���G~�P��b�~ �1u��"�6�0�x�+a�V��1��6�5�J"T����T=��Iq栭�;`�D���b{�׈�eL7�P�����:bљ��Xb����\d����h�;�S�S�9V8����������&T�J(�X̷�>�_�z����s�X��-�m�6�S?�"	MhG��io^8��3�«��������Gk%nRj\�� ���:������y}��{̌��;����R��
Ι,�4f��)�V�[�!����~�+B��RT22�)�ҿ�)��N�O1\Q�]�[�é7̟�X�Z��x�� qi�{�>o`=X�L�p�̅!�!�����lu�ԉ��'��Z6ｙ���9�G�K)��_�)�I���_�q��U��dN���ZGx.M2�Z�k�q(dN1 �P��S6H����Ɠ,�ƒj���X����d7&R�Qt(!%F���[%Ri������X���u������0�oe��� �u���Š?���㑅b��l[s�<^GL�ߙ�c�di��[�=�-f�#0�G�>-��*�J�|�X�xy*b��׎��l���%8���VY��u]F���杅����pV��&�a��Ẻ(Vqv��.��b�|�H��x��a�4 ����a�r����4��?��Y�o�1�5UղK��@E�)-5�M���82e���O��=]n�^����e���i�A����
o�>ɧ�!���m�k���rQ��=�n��"�\��L�*t
��6x�*�]n����X�(�1�<�W25�����yx���d�G;j��^���lS�? ���V�w��2��I��/��Ͳ�=�SS��bl�b��T)Nh_O\��	W6/�u�*���J��%�}��מ�W��ǉj�G�I� G�ι���gч��&t_g}�՜h��@QH#�
�C�ej��c21H�ӓ0���"O�\G떌	��l���}Ԣ�C����i{�f��}�,��p��g]�>��-�P�Y�氍V����m�o�.��۩0�֑*qOu�����J�C7���|�ߞ���V�Ol��QDuvӨ��:��I髳�~�����㡤�f���\��z�՞���i,E_}�j,��������}��a2O�O�Zy�j�j~*3�~~v��2�{�P5��b7���L�kͭ��㽍�!D.�Nr���#���,ر��y�aO�Y��Pu�yG1�핡b\���v��0aY�S"(��9V�>�Fs�HΆd��oGTo��`�z�P�����,�f>8Rm,�Ќ����Ҕ��2����O�a�(s��k�P�f�568��A�f��v�%Z�5�w�,����z�ع&=Q��}�/���X�Q)r�z+�M�e�-7<�����L�ז�F�nK����E��o�^�-9(��ۚ�BF1��� 7w�ْ}�!1Kar�Q��{�G1@DX�K�&���Jl+,�{Eb�J�$�l�5���^�ڽfo#Q��?1m��T���ĕ@�8��t��#���������̶�ߖx��v}��![M��:3Et=�Q!�G�H�)���c���J2ఊ6oG|?�:ra&�^��-m��
ء���h�n��>��c���Q�D���0�)�;躈\}#V�@�(�'�}�B�-#N��	�-vb$��դH��]�E�k+zJƔqw�M5l��$F}$Yd�&��JrJ�2������PlmW@i�N�_����f?�AJ�ɕ �~�Y���|_W��&@j�%�	&З�_���.���w���B�����I)B��%Q
�ɏ�M'm���/o>�Q��8o��OW��ʁa0�32�<v[��s��-�$��nMdg����j�f2�z��0��ZHЩl�ۿ-G�g�7��I2y���+0&Aj4R��[75��n��*�k�nO�mq�[k��B,GPn�Pt(yH[Î�C��R���;�F'�$��������[��D )1%�Ro���~�E�8�&�,���]�,e.�l1>R]����+�.خ�z�r��,�\����D��\qR���a�doXqN�mU$`2��BR�3�,��#��؇�L��*ˋ�0�e��9��Og`Ple@Q����f�(����C��:οgQsC:�E':��:,�@���M�Be��$�94P
�r�����>�&��$�nQ6	��M4�� ['���\h\�w��s��ig�� %O2�zrhɔ��=Ka�J��d�wp6wf����,~>`eX�o{���]�#�L����t�4�ɫ�ZQlQMBń�ټ�n��H�)���r����u�� F���2Mw�x��1p�3��4)N��=ZR1uGJ� ��j�4�*i{��$=�&�*&��=�]�[ZF��#7��#�T=Q�Q��W�����#�M���䢊���b�*Å��Z=�:Hhw��O@"�D;Sn��m�_�11_�p	��VIN#=�w��?�fWa�v�rE.T%Tŵ�V��DƎJ���F�p$�tZ �o��O��	�B��ljR}��)8qG�H�M��b��5PY&�f_:0疿.&�i�Yk/��U�'_V{n��oٝ�����(���E��S�H
�f�d�@Z���|���O���^`���7�P�2�0��p���4[.�J�K��w%s�gID�"`��J��/���� sȱu�"xg� [j���X�(t����㤠���0���PSS�b��(�>s?}���c:��p�U���j-��\�_e"gJ�`I^���/�K��M�4�&�#��l�����A/[��(B6���`��j��I�\P�Z���(BaC�.jzo����wt�j��))ż����l�R����@J]�V[!U-3g��IX��V>�A��ۙ`����+���m���4��G�"�趂[J����O�2���~C�m���>����i����0��,��ݑ	�&�2�!�2��X�Q���e.������4ءd^�4L�/c����=���y%⋁.�J a�4d@��u!��ׂv�|���R�i	[K��'6�7�o?�A��=sh�ˊ'Hn��-fK]�����d��(l&�?��a��%�����KW!_����@OT���ꅘ�b<Z�9�p�4
ݢ�($w]�"BP���KCY̹
Dۧ�Δ��!/	CӇ����_�nf'�����ʬ����Q�5}��;�3	�-��WU�[�)��g�8�M���w�n6��7I9X��`�6 �H��-�ar��Z��\Q�9�4˱8S�d�';\����f9�[��u\qל�BB a����<���+��FCr�'��^q�zp�7be��.�y�G��(?p����#�x�� иmf0O\���kEh�X���	�Ԛ,yXp��3 �{z#;V�/�\#Ҹyes?C�� \ͳC�$:����g�TNy�v��d�3��'|�yL�P�a�V?���:����Yd"������V��ВBA�u����s��c�ҍ~����Mh��$)��/�����P�d��z~W�$�͂�|>	�]n�x�l[���ȚP2�u�æj�#�T:�y�5ߙ��.��������x �&�l�N��"���L?��4X��pe=��[�&Z͍iN���Hoj\h���<T�{S˦��J��i*�����o���r�I��ن5��<! �S
k���M��Aw�9u�lJ���U��ܗ�<����t�wKn�)T!�j9"��@&+�"����(��K�)����l�7*���e�l}!��$�1�,j���=��]C���Ƌ2`V:h��)�3T��MP���u�m�)`�<<;{]�M����L���0�p�T�tAn��ӯ�9��BD�B.{�^]�er�2p�Zng�a%X�z��6��y&����|CIė��s����OؐX���rt��]8��Oĺr�(���9��D�%� ���L�]~�#{�{H�*�z:z����1���ZL�~�D���a�k[��:�ў�͋��K���t��H��h⻞�b���b���&�/����S��p'�5�x1ɱ��oօ�,P�k�y2�ɲ<6t�[���.[7J�k����,^�X?���:�W�TL��T}���i.q�sr�ٓ}1_?��g����>w0/�	5�,���b3�vdy���2 F��9��P��z��&���bI
 �&���ƚ�E�	U:�A��v�o�D�[ ^�S��Jw�go��&�8�-~����N\L�!Y��q]x�p�ܲ�W35}o@�LM�x�m�@�s�^N'�^!C��}zC��#T��5��A'���y.��e2ņ�[��p��S�	����Ԅ�c��ӵ�%�C�[�e�k�饪qn̋��7�ǻ�ñtz�#NRX�-�s��9�m~�0�R���H�F����S�#�I�C��/a��?�Z�!���U�jF�d8sV��kU�[�ض�U��>�ʴ����dpG�NT\�����X��(6��!{��x���Qy2;v�t�b�Ed/��3k�M���{���[�,�ەN�R�HB�F0�/F�+���@ЈQ����=�Bk<�
�[�{��]�����7�ޕ~@J~c5Q.�?X��Ey%�^�Og�LL�bG'��(���1�4�?�;zN{>�3k��]�5��C��$L8#�{_�&�������~>(�&��!��<��J�7�"m�h�H,+�G�ڻH�RbS[��h]� �bJ4��_Tu-��@@���b]�x�g�j�W��i����ٖ����Ħ�������*��^����*�I=hH.�@����W�@{��{^��m�;D{�*Pγ;��Kd�nck����Ekg%[�D�� -����^�NV�ѳ����~*����(㝵�}�̔��i��E �v}'�>y���R��y6��۠����q,�r����:��9�L�bB���*�J�c��S���4�k��2c�QMX���e�����[I�*0ڬK�rc �%�b�P3�s�f�.9�ٴ�BB�?�U1C9���ƾq*;S�J�e�ҝIZ�
�1��p%2R�jh�䍝������J��9q��]_��]E?�&!n����3![�qLUץ�WZ��+�FM'����ۍ�
����?[�0]ԑ�@��)�?f�7�	�`�v���j,�u���_�M=�A��3_ZA\��H�{�q�)�ڬ�XD+y�� _5�̡�o\�<fw��sj%m�� ��+<u,�)��,(�V�a2�^ڢ8%�)
����?+UW�{$.R�������v%����(Z'��-*�0J�j"nU;p(U(���ph6�*��e�zKm;�ƭ�B&lz�t><�Gr�{����/Ci��y[�����^튑�٦)M�ߩH�L�D�x�֝O�w�t���;+��[�7�Dȉ��t;���b򗄭VH�0�p6���+����lO�[m�y�3���#�	d���>���Z�v.zEzJ&V�ۧF�ڀ��� հ֜Ct�����C4�2�n�Y�%�3�x?��}o�:�.���O�U͌d�~ޜ2I*��a�g�и�؀�3 �5���J�{2
d��=Ņ��
b��,�����'�"�(Yɑ.�f�Gw�Hb���X�B<�h��������Jm�86׎S-��)h^O�ZY�=+��w�NS��p^���f��:�0�t��xXW(W@�l35V4@F��$�)頞`/�c�wv�2���=�3��_��'
>����������̬�4�����ȿ�_�
s�V�iN���09�R�)
� U�}�uf��`8�X�x6)1&��f�*�ΖXI��u�,��˚k&%��6D9�)�t�_�o�����eW�Z�~<w3_P�^�?��|�DA�<����.�qe�b�V} ���l¬a����X���J<��eWD\)��Sn����:#]r�F��U
�7��B��؜UJ7��S��J�3�}��&����R�+�!����1^,�Sz�D�!y�Z�W޼+�_n8UR������qW�T��Z�07y���\?Y�d�n���3�<��>1B8��U������#�iyY	DJ�E�����;I�<!;�?5����Ey�ݞ�xH:�ā���h.˘[�6�$\ ��,�q�iK��n!&㲜�Z�^#����ܬ�>���^J �����-v*t��g��'�<�h]P��.�;A	]���,���wZ(����Kx?��ni�&��|�jA���EK���x����Á�A
�]�ȝ*���=tKa��l(N�i
C����%k� ���47ḻN�
��*o�!0��!K�K��o׿�l#���z%w]W�c�@%�˺y�!���ώ�ͼ*ߩ�3�P���P�9!�p؇��j���k��-,3˕���d�5۾�̠/���|�}�g,]h�H2b�ύ}6�+T�JF�-������K���h1��5Z���>(����-2�$m'���� Z'Z�y�+��4D8θ" 4�"H�Hv�I���F���+ �͑-cz����RC��x|��c���+Ĕ\�vd�w]K�)����q`���ʏWTlU �(���<U`��b�n�@���նrɸMiZh&>|�,���6��7�+I)�����>��7s�'�!�;K>�~\ t�H����6�\��P�O|�����\�Ud��y���/�[��iۯ{��|v��rN9�i&|�0 ��h����?0�臘�}�����g���c뽿�p��b"^�t�R>P����� �ѥV&���Y;��q�4��lh����Ў�n��>�$E�e�ҿ �0��d���lʢ��8��Q]�!��n���#���C�
i&��8"ZP�J(�N(�ڇ��k��k��C���:,��.�w�ލ�o-�n|�_�vM�%���Vg����?�-Y��B�P�G�|D>1ˋ4X����cO'�Ҙ�g�_�9�wm�x����V]��3c�>C9RR��h}zJz	��EkѪʔ��{��ʌ���\ܸ�p��{1TRp/6��nXU־�E�C_�c�;N���R*�2�>�;-���<��何+߮�=S����eP<�!��>Us��1�<'"6�͈����=�|�w�N� ��&�DX���~soy;"�����P ��r	k�O<dNJp8�M7Y�aS�!.퀴�5���*�Z���J|�a!� 4�_	��V�[Hv���B���l���sG�� �� �`���aug��!k�*^H}�YO�j}�0!��^F�b'w���o�߄\|�q��� �DY%[䙟G4��'ZE�/��)�;h�˘�L����Ȱ�j����ms �>�=ʞ��Y}y�6ʏ�i� �2�Y�$^>�g�U�b��7��$'�H���%�!]!��l�j(7��&��8�C��1�lQ�ՠ��)F��_)��{1�v�Y���ǡ�J��s�����9��ُtAH7�]�!ub+v�y�1����rx*ˠ�+�'(���Pu�Jw�!VZ�}��0�' ��	�'ӨZ�T�pk��������L�_��=,�7��*[h����L�)L���[(3�9ͺ�,mE3o���+=W����� ��.N$�<C3"�=i^N����_��E�Q6Ab���lU\��+'�h��C�ϖƦ5i��CrG�֖�0�M�A�a~+|�:��ۤUZvB�=�D�i���R��\~V���/��ʣK��Q�`��[�1T�L"�,�L��P�?��eo����W��i�W�/l���n��3>X�&Cd\1tm����l�+o��\�Țo�n�q@%�"���?Q^�ѰM�nv$���#��R��Y=}���#�i¬�!q{>�����������yDY�H�=Q)�eE,���_ࡾ���mKƪ����`��b��oR�BU���>#��~�����Id2[qET�AJ��SmQm<�����~$�a��*���՝1��|�	V��1�C܇����%��6]�\��%i����nxR�&�75��S�^���;V���ic�~��*� zҝ����F�V�b��k�c�����{`�0���N`���Q��q�U���փV�ߝ�����*kŎ�8y���_1 �E]�ZV��E�!�փ�D��dqe�x��_#EM�A|Jok#�UA�-�Kq�|a��dx�Q�q�;���[�P_m�0w:���x҉c˲��Y�)��[�|����Icˈ�m:���P9��Ue4J���NdK��V�QD�0�f�@M�b 	���]tp�p����þޠ��|��I�*���Y�3Y/��. ���P#��A2e6�R9g9�K���N�K�T�6#{W�����������c����"��C��,!29m�� lW�&���I��Ou��	~����x��0��w�5h1�B���l׬�ʧ�5��%�ͦP�@ϕ��&���Xr^�^�0��x-�9Ilʡ#��=d6zZ�j��ʕay��"�N�	F��(j~��&%��P;�ҡy��4	���F��E�W{Y�e.�5��n���ϖ��#z��l�o�~��]pd�ӈ��鋀�^G�Z��x,��D�o�o5�C���u8�!�;2�";�,U;sV��3��fՇM�m���d�'�?	��O|gn�<DD���O�6*ķ[�`7A�G���т�2�N��T�\%��� �k�P�B\S��I��|�-w�j��!��߬2�!T��r|_֮�Y��~����b�co�=��{vV�ސw(K�gzx�;�J�p��ƃa��=���m�Hы}����Ⱥ��L�[}�U*�%�d?b�H��ظ&T��)q½�O�J���G(�[����:�ʹdU�ɀw3MR�j̄�с��#Omp������3;(��
������[�/�=K�i��V�F�5�jt��S~7H�gy�P�5��;��`x���:�P���ns؈mLL*B��
*����ɶ�ۻ�:���dz�U�Z?���m���]������Ia�*
�Ji~}j8�|K��E4�o�y�VA9������u��)�e��]Ԁ�O��Zy�W�e'�P����*|[.��j}m~K�gT6��u�	S%���{�M�@Bu}��f���'ɏhy�VH����L`V{�@���}�j�Z!�������j���f�߬�l[!ʩ�]m۠�2i�a��Z#�M��Gd�IOL���I;�C��2+�j2��,Y��E�Ak�`�Cat�/i�k"�t���� ��\�����Ek��˟��=��T�<ꅊ<M ��
��)�J1xE75�^�1Ih�!?�<�'�sK=�bg����6�<��w�H/;Ef�J�a��\ە�4͝�b��Z<	L�:�P��+�3+$dD�[�Xf��ک#Fw�hC��α��M#�@�m���Xd��F�4A��JV��,�輇uS����ۋ� ��2.s��s�w)��y_Le�Sj#�����)l=^}�Z�2�uvZ��`|�v�0��3�Mhk�$)��a���1�.�$�=��`���Ҭ�{�2�m?�ج�^<_!op�
�$#k��M�-NO������y�2or����_}ļ@�=f*�&�Bo
�w;�i��8��R݂P�˪ΰ���F{�Mp�u�;N?����P/˹B��xS�Y�R�ڣ��7;Ͳ,�Q����\Y�*a'�EH��Ʒ�دO�W�V��J��LkD|��.Y�s �`9�����A��@�4k<�`���	���>Z:8lQb��E.@��c�Z�>�D�-��3l�����@��_q�,)U��m����1�`:]�K�c����8����Q*��4� �$j��<�s/�c]ps��4�\��#]�A:�O1	��œ����~��k}9�K�Fڲ8c�s�L��׎;;D��L9�~�偶�l��H;�sv�l��QK.��ӯe������g�ũ����z�oԺ�ˡ�i�nFkV��<V����ˠۇ#��I��0��dEg�*5������,���y����Xs���@�O �wh77���ƪ����X�u�4���Y��E����wv��a��J+[\���`�����)i����p���7�&��o�� �`FAF(;�x������<�x~9����5e�ekM#@�W	댫��,r�R��3�ִ�'~����y{j�@i<��������3��I��v���4㼎��8��
�zp|?�t߿�:ٺ��	!�d�s�3�U�#�EA^?��΀O�8��i�g�����@p�� �y��I&�'^.f
}�r���N�	�%�=I��E�F7��V*�̮��M��e��2��UT�:����34tX��y��h^U�v�������l�52XG�|Iܓ��z].�+)w�ي���We�ڰ������7�����YO�Q9}�[�yXN�@����`,�+j1��-}L��(	M,�W,�s���p��Y��]�T��WT��	[ �)�� [��xm�އk+}����!U*7lHk��Eƚɂ�sn�1����/�
��o�f����M�B��2� �:�㤙���R��{�8#�Y?렺�A�;��D=�~�XS���jفFO�򠄡�(G��&��5����w�~8�.������$�tڏ���hE��j鱇Bu�Ox!Rc���n&�O����3�E_�rx�[~ި}�fE�)�Y~}�֚��LH��S����O����pK�/4I����/i�~	-��K**�� ��r��^��ےVYr���&b�j��$��X������q�FT��w�泬�⾯҆�t����|�G�c֜��0P��Bŗ���Y�9�oT�/����鰳���)��cy���w�K�"㧙1
<"���㹢��tN�c:U���tDa��L�3����N��1����&Xr�({d8+��,1	�����LKbAFƑ��p4�x�b������p?..\�!��]+D�:aq����f�nB�M�5c7-� �+��L�����4T��+��&`�/�m<��yB����d�|��Z�Y�O5�K݇L���Yc��O�^�����thB��sk�#A�Dx~<	���9S!^HBr����z��]�E_jK`�ڐ��P�M'��+��x��?t�cP���t;���z�������8$0&���)V�x2�6��ɩ>X��I��af
�:��z� ^5�s_�Rwv�z2��n�򓎼�w6%�H�3ҵ�����O��o�<0�q؀�"�T;y�68^mF�DotC��g(����^A�������P�7P��b����O����,%�#�(Ro�SNd�q�ł�W���d�߃|��ngSc(��M}W�C����d��+��g�D���/���e��v���G��5�?�M����=�јL��zxw�bZW;X�|�coO�2�V���*B�H�H�#��S�@Q]yc�F^r�Xs�9=� 'M��QBfe|3�?p�1᪢�~�΂S�~�8R6ɣ	4G���*K�b�s���U �l�H
�=_��H��Y�[^,~DL��^E��;�R�d%�������8�T�%$��=+�aF����ڗ��i�k7G�2�]�V�G,��.���3f$������� �>��UT:2[j�m�u�23c�
�ǡ��c`./�j��@���ct�S��H��)��4�o�M���1k�{9�C)�m��k
�<�Ȳ�(�U �ʕ�;L�Hעt@�n���aԖ^����Q�c*%(��� u0}` �&3|v�}��=�<'3J���NO�����q��F�]#���!)SXu]M@�'P�F��/6�u�-1g�'�B�f)Q�Y���Z��*KS'�r�3�.��;.~I~�|e1�명�f�v���䏐<X � WE7���,�8M�鶻c;:n�CQ5�ua��f.�zǔ��M���Mg�-Ռ���{�\�!�-�y3���@-��pO5
��ϕKϲEpǍщX��O�.=Cx!6��ә䘃���=%K7���|2uzW������d/b߬�������c�UU҂�ow`��[r���ĥ����(S}�����8Щ�LП�u���r���A�]�@Njm�>x箅s���7Q�R��$����G��+���qC�/.���-��M�U ��9��^���2�Q�<�ω�V|���as9�qT�L6���l~|�͉�6z����7���M��᫁�؈;�8��%�����>��+I�H��I�����ωΥ"�~�Qn�>��w/g�΀�Df�}}�;3�P����RaZh/�D������{��s-u���T=��-��"�D�:{���{I�Ĕ>I|R��x]*�'��ވ�c��Z�}����[>��nޖF�#����Rs��=ֈ��rr�����X!������apQ�m*R��Vk�=#e��+��5~�r@��y���κ���/*���4��)�"�2�S _a�2?<w�@�$�y����k��L�Ɍ��`����0�v� ^�N=M�N�\�P+����;i���6���F�V�@����+���}�I���+�g������ȉ8��mO:��:nσd̘A�w^c�`?�XK��������M�J!��ړx+Ni;���#%�U���{�T�"z8W����ԯ3��7��q[����u�rY-�@�5�:��r6S�r��3������f_��c��?��E�YLW�L(	)ڱ\�0���|9w�7�>Ml�7�u��8[���xN�aRs���-����!h��d�����2Mb+�4'�"7+9�N���SXx�_���,��"CsZ=���9���ֈ�J�l@�q3P���ƕ��6=����K��y�/p�!�A̻@�r��9��2�\�^�ͼ�`g4�+�|���A��V�iU�}�ֹ47Y�'�_ι����D����r���f�UUfw���r�ʠ�톻�Zޢ`�Ke
�
O�'Vy0�v�I��B�U�� 9M�&!É���?i�R_��A?��~�X�M&	�~� Vq�ۼe� }P�{}З:�¿R	2��}�� �"9��g���Кy�8��T�ON��e�J��M�&9(����{�ctv��,;S�J8xhDd��G��`�=T-=i���|翦/R�|�k�����@@�>����v3�����b)�7��}Nܚ�HG`�|
����J�����:���$S�	��c��Py���	�)�)�n�%�_&pS��+���XU��W��AUR^@�m��w�ӄ��6O�_ʊ
gcx� �ڗ2���KZ�E�/2��qO����/��	Urw��@����sv	\]i,�TjHb�Ѐ5�dS�R���v��$зA��Z���w�9�鉌�pP/��U�HH�o􇗉Ռ��r�HI�E8a����9ҒhN|h@��v�ʸ�7r�|2��$n �'(�g���Sh>��.���|a��0��X[�$���y��R@�&z	�za����.�
B��[����V�K�u�B��P�������3�.�y�R��#Oh�][�~V�3LR+k6p��܃��u��Z>9g����nm�v���Á�[�Z		\z,��s��\�����C�Yc�_o�w�"u^�p�1��{Z��s�s�����S\2ͣk$�Cg�\�0�-���h!���w�'3��'��[\r��"~��r��h�����R���QI�gM |��CZ�|c���̨��~g�S�����:�|G�1B�A�`\��ު���!pk퐨�����m��GU-�޿���H��y��}�g{z �~gg�Ҵ��p�&�yV��֋h���	i0N4��֠nBh�۴]�����/�S=��"X�Ԋ|���
���Zw�a�/>sY��7��C�~��w��5��1�
F�oZ��m쵟�ܧ|fs������z_�h<�؊���l:��J����yZ������-qb]'@nx�:��ո�$��\�R��`��#������&��t���Nx��s����2�Z�O\.�C|X�l��R�6���Ya�����k�������;������� ����4N/|NA�Y�y�K�|�ռ�T�u���]�<Yd��ӊ{.N�M�1{@8�Y���bJ�W`x�)���L�ۚ1�9��#�߁d4ڕ�+0}r�����z�.��4�P�A�Bϲ�EU�:���X7܉��NΈM�#,���6��ǆ���t�ds��5t��t��	��#b�+�U�bڻ����m�'>�7=Hr5�f����w��`�xcY�p�*z8z��4��krGE��	`ڀQ��%�&�
n<�Ye�a�����swӘ4�/���Z��R��uS#���Si���c'�:���t5�@�Фm�ڏe��=?��߇`Nq�V��Z�U^ %G�n�{�1��v���盵�/�Vl{�Y
%i�nZ'�h7,j_�3m(E��P�UB�¬E��D�r6l񖨛�H#���q�_��nXC�)��/l#q�cz{�̽Y)xw,�Z�T2�dM!���rԾ���3�Y/�zn-i��_g�p\�
~��3��+����i������}L�����ҩg��%>#�^�A�E�Q���d�텩)�C���&��#E-'5���]�뷙jA9�������]ǸV���EV�}.�$�^Y!#�j�����Q��9��Y���I˘�Q���Z�u �����{XwM�)��O���m,�I�W�o^y� ��|h+� \�}Du���,��A�;!@�u)�G!���2�(Ԙ���}��^���
�#R��#����h�ꞂzN���nH����2�Hs�H���AeG��t��?\��ٔߡ�h�8D��u�_;��l��! P.~�rm��J�t��P��v���l�Cz���iʫ.�4%���@���"�8��B�z(�ƚ	@F	&.���I̍Ԫ٥������A�إM�8�Q�t�ր��V�z�m��^G0��o�Uj/FG���gK�=V�e'�#���TV���.�oYi,'8t���8u�ě7�<�Х�tF܆<'��@Z�i�����v^^;�aJJ�}=�Qw?BF��y��(�(�>�iiƉ��� ��S��O@Ə�I�c��gV�th�'�B����OsVZ�d��!̍��x�����I�h���ܛ�^<?�)71�;�0,�GP��$&�W�XCt����-��>��ˀx����@5��k|�JF�>�U+���2I�yV͓�] �	!XX k�:h���B6)6rY�~�	�V^vU�2R��O2�`+e5���
����dR8`)��h�g���>g�7>2K(b^e�Ҳu�|n{t�e��_���|�"9�#\ ���c���;�~!�l��>7������:�v�����t0��n���bXy�������y	���hܕ2ʕ�"�y�9�5����+q����Q�]K��烂<
Mx���P+��d�Y:_w�i]w=X��<u�������# �0"������Ue�fJA�������bJ�J��-䢮h�\��U�ꩆ0����FȜ�O)�3�x�3�JU��>1���k萲.�����ǻ|�:#X���З��Uo�HO�H��ðn9Ȁ�B�Ղ� �0��Ҋ�ݚ��7��ۀ�h�#�v��u\~%�YpZ�SMI�
��j��y1��Q���P�?4$�.�C��14ܥz
��Yߝ<�P�!������/u��B��u��?���"��%8�齞fŚe঵��A�(�9�N}��"w�!�sDT�j�6�E��YdD9Jq�Ly3�;��\A�2,�3�]�Slw���E���u�>'ٙ���=�ѩQU��<�Yۥ(%�%]���-�(�v��&t$�~��9u�A�Ώy�3.lB�1K����<��@�]d.]��t=�1��F��`Q	�X��-)cu���*��I���37�~��a�g�Wސ84��NqS����]��� ��$�ҵd�0��m��ߓ�u.fj���H}&/���K���y���3���O
~G�E�byCݮ~��J#ڮ�h�+꬛�|���@�v��_K�����ϣ*8*.�`aV��V�m ����@�TS�Oz��p���~�ʒ&�BhH�>�X����d7����F,��u�d��(V��a�6����6+a�O��=�"#��BB"<��X�&_J�^ۧ��v����u�����Z8����yI26��jI����r����3��j�{Q�m�K^2��@��Ar0 pVl�SˮC�>�~��s����b"�&բ���Po�͜2�Ȭi	oʜ%�,a��VS] �+AV6�����Ϊ��Д�bɂu��c�t%R<��X��E��΋ݼ�y��C��iD?˩��X$��B���6G��f��� �Ƿ�6�2������$	%uQ��iJG6�!N�?�Q�I�i�)M����J%^�s�%�T3��RGу2���@��V�`�Sָ�Ef���?��mM;�س���6wN6@�I�&����Ɍ E	Y!�g��(G�v+#��MH%M�C$�R�cL[:O-�`f��W��vP]��2������1g��@yu7�;������yy��5Uj#����%���N�&KF�9$�!�B�%�0� �p������}e�`��>�M��ӹF���%o�~Vr��0�c��]�?�?�{��OJ�TOU�
��Q��@��G�]�0R]�������5��Gq�nz Sk��~5:/�X�臬e3�ĖD� w�6������&����-��ջ�W��d�����~����|�<F|_{[���p8rr�jef���G�덻؀�k�/��p��3�$|�al��7�OЛ�Ύ@����)�ɹ��
@v"��������X�dhέ�N��'3���o�}~�ح��{F��q̉-<�\�2v�$9
`��Z�?�@Q��q`�:��b[�����)D� ?УdQ;w�[��Y����b�J��1��ŠF�I��p�$v�Vs��b ��@a����B<R4�Z�ף���`܊/��L�qȍ�)�������6��y�KC�-\Kĥv� "���<Q��﷜$[���{9��׆�Š��r��?����W����'ϻ��m�>үvq�R�YXI���]Ԏ�|T~����k�݁&� >rs��&�ċ"�&��^��<71��c���i�uO�^e�4�H#������>��9�V��=�_�Ƕ 3��!��&�z�����ߣ�2��V�!>������a>��g0�ɰ:I����h �ϖ��'�\��a�1a�]��_ +�E_���a/�䰌���?X��x��8t@�B�)s���}��`�����P9{��s]Y��f�.��%�0.�ٳz^cO-'��q�]31����lv^V斌�k�B�$�0�(�v���ν�@�����i�te��0x�UK��=�B,����f��L�=�*m<</0+�0��T��Y��Bj�r3a�Kvt�y��p}���Ej��������9Q4���(�8�Gbv������&�̾��-v}�
�"��r�wB��&����z�{�&f�N ��e�0O�h}g�����᭖$��	8=f�:��^RU�!�I�f�kq|�	!0pj�A�[d]�!�ְ�K���.���"i���)=�|���$K&k�J�(2��pM�y+ѯ#�!�����+���o[Kj�eC���IyY!�@���I�����|���39�O&7���8J*���M�����|.�;,0��"��B�{�`�k~�[Bgd?�����tl�}��P�1U���$�Y�f�5���\8tct�'K'>�m���G-X	6p��X������?�n?BO�O|2w
<C��h�Ĵ�"��u��)Z�<���Ro��p� �z���y6~X���7}?3�IccҒSx��C9��5z���>��0�νY\A-� "�����|�e����r~c��P��`�X�i�P�22@��*�q����Nv��i�}15�[ �i���������������D���h{���I�Ty���twJ�|�t�#��V�[�~�BL�	"(	ץ�(�L��L%���=7w�&�_86�2"tX	V�ac��2�!�H�Ƀ\�h <��.D�MW,�ڼ:_=���3�&3/�B�n\��E11��מ�'�HG8�9i����.���l��WK�ֈ�ה9��.Z2���]������I�}G����'#���CBfG��B�(F����zu���t�tx�if����#�A�D5�Q��@պI�)�D7�}��`�u��@�h�������T\R�?!F��rzi�"��&�V�ý� ݙ�{��Q ܔ
�ЙcHP/�M�k��R�L�[j&��v)�HS�����^�yO76Y�z��q��C�'����F���S�N��xQ*ؾ%�T�DN����K��E$3t��1;�nN�p�L�k��g����K�c�D��=�M�;f��;�Φ������8�@�g���"Q�[v����-�-�HV�U}��D�Vc�8�pxi������QN�Y����K���W� ���sC/����/m���?>M���/Ĝ�(M�lX��I�c��D�(�G5,7�{ϊ3jy��fDx�V4Ӟ�WG��'���|J"f�!WȞԴ�wc
���ě]�b��z����N����!|'K����?q�j���J��2�m+�!|�_]3;i[����S���E]��mb��}�1�a��cY��	%\���\�j�}LK��!�)��8�N��w2�B�w��vښL�I��h��^d���N��%M��.���AǔOTl�!��#���J2�q�l0�y\��EGd06w�U�����h�
�|=�tӭ���K��֝"�c�Q�2�� �"�������
?(��(�ߥ}@3��;�PG�2\�2.�Sr���� g*��L+�����\mTN!�G���p��kȎ��w��_��Y}8��aݴYC! e5I7&IP�\���ÝQ!3}>�F�9���.8{�	��}���&���Ugs��+BJ��N����{|/�=��6�#�H, �2ea�K ���xX[��E^Ēg{5�'����Gh�(�"8�,���mR1ݻp��]cw��co�Z�e�<f�Sxn� ��Z�%��뵀XG���,� *
/�t�3.�b�r�ͦ�������^ܛo-��?R�]��b����IM�}|V�O��s�q9�bRۄib�L���{��GF�ɤ�%�H%�s!ƶ#�r�Q�{�a��2`����lm9l�\�������t��dŇ�4�-��%,T)�J�>�>@���`����>�~�}�4�E��������_lT�������f��c���T����P4E�����a8ez��-W|y<�ˮ-Y"sq�,�M����||�緺�7��+4a7��˻�;]��4{4�bzV�um��0;hXŗа�0�^���+���x��I�DY3��p�_{�wK��aH�k��)�!�'e�ȣ��b�g�|-��G�|��󽾭��r�H�M{��� z��;q�r{��峽���!&��N�����첟s�*9����\
�� �NlA��4��Elڟ;>�=P�'rl]8�6��R��ʝ)��F7U7]��|0N,���֛�GG��:��)�k"��Pyu�
�1�J�_K��<\)������7���A��I�-0�1�T�?e;��i�H�ɷd�
�: �0�	����x��/�\�^�r�ҡ1�.�àI[���c*1��q�w���Q�������J\i+�� J+*�	X��9��sr��KVI:t�����^^Gn�ZZ�N&G ����8]�D!���5W��J��A���g7 ��9iM�s�1�[o�W����YjK�ʿ��j~������
>�e�E.��U�~}�Q�i�k�J��fś�0���<�߭�K����ܓ���37����|�s9qz�����Tq�r�����q�^��)wҦ���!M)�E�X��z껋��o#o�;j��s���I�2��P3�hhwxw������XM���^��+J���V�G�|�G������Aw��0g �]))<!z}�1t��H�N�H����|��燆{CaoԻ�_����.Z���m���oQE\2S��������%
A����v��uL~�D���ݘU�*�EہØ�!���;�{��Q���8"�C2�$dK�Íj�AG�����0kx�Ah,M�rٍt�_A�f��c߉�$�N�GQ�7��7�0�Q����?�?� �[�2������a!qWoW������%8�7��-�� ������7����sl5��LVXhk�%��;5-'��)��3$i�F����
�S6-*�6��Y�7����n�Al�A�[C5"0�
�_��B8*q�V+1�hsw�g�%f� !�Oq� <�)dʘԖgZҊJ�h��i�):��<dtEz�G&�J,��s�-6�����e{ú��L)F�(��;��`x5"�ZF��z�K�<�˒�zm�{���*;�t�kv���}d��ڋ��0��$dqr6A���Хd�S�B�
:2A����N{��/d���S��S�:���X㯛�2�SRPL9����?LE_q��^�\�桎p���J|����1)�����ι'kMK�J��.��>�t�Sʔf�=46�L�9UTa(�e��+�nP@�t:_a��랳nm��|����`.{�5��x��~�-�+5�}J+�ZϠ�`�['��4���)2�|H�A���pܷj�1n$�'��N2�N�C'&���~�mt���J,��3�l'ZՇ��pRl�+AO���6�mdz�1o��,��|n��Y�>.R3�v��.�U�+�˾rN��*5��%j��+��J-��RS��"e�v��$y���$��`,Z3#ˡ�Zp��b7
���sF��� !G��͙+`I)�N"�i�B{������k�"����5�B=g�p�Q��}΁�c������3�9�3H��:nr`JLDE�U��#�rv���$˱��t�e�k�aA�ʭ�;��s T��嚶z{��������B�����b\���[�#��$��(!����2��r6f�Cۦ;���	��?�}����
���M�kl��f��"{���~!if{��voGz���/�Ɲ���:�c�r�%�f	�'�&����ۤ�;6	l�
A�k��hj?��$�2d}f�ݽM���+��ʒ�E��ĭX������SOL���O|"�ac��Lʖ�dn���~8�P��L�D�ĲF�Iȅ��R����+�y�Fr(��AH(�G�V+��>��$��2TV����Qd�嗩�5�Q� �Jp��ʒ�F�Ԉ���)h����l�3���8�Ɗ X�cc-�E����
*�_ȏH�?�f�:,��^�ѡ��u?���"��$���I��j�a�'m![�?.�I�0�XA���~��%r#���۴�(�q5�2�?��ă�u�@H��!n�G!������aB��|
C��Z(��;ϯ���㛲��	�x��Ոd;
^�����Ϗ�#j����bC�ŉ���3@n��ZC0�~��c�0[�/,��G�1�M�;�]�ŵ��KF'N*�L�B`�����8���ʅ��\V�$F�АA�>�b`�#�͵S'�D���ߗԱ�WL�sD��<#��j����<�xa��	��7��K:+�6�uF��0���pr��W��tǅ�iU�EI+��o��B;}�`�y[�j��H�\��O�d($�n`�l6���&:��@sa��*�ν{]	F=Z��NBY���Jg��!��Z�7&8r�&.H�1`}B 1�����I���>=7c�Tj!^�]����e҆���7���i�eQ��Ziߦm"�:��|�%��ؾ�����ٴ3A��<������@(ؾY��[��=J��
lU
83{��E�jԡ�a"��nw�/�dg�g�ӾfZŢg�N�`^�Z,��M�f�o�q(z<tcR�d]3�U}ab�ά\=�j�[�ҳ����ZDS���(A
�wG�HL]x\l�A�PW�wyXr=�.F=�;犇[��i��K��(~7K��	)=!�) ����+�ӈ��Z'O���h�lF���i3$��8n\=��7J��ck�g`�l�66����s���:��Ⱦ1�D[��麏�j���~�'���/�
/��_j����Ѯ3����F���ٸ͎+��*�2�Ee�n��W^��	�l�-���b�b|�)x�.[�ד	���ܘ��,�y�,��3�V#�/�d�s�S䄯��-�ܮt�J��,��&ܦ�s&(����RF��6P����"��߰��Ӑ�����(�Z[���`i������
9�Slæ��մ�W���S��M�R�R"�wP3^PM�ܬ|�U��y�#(�yAuԾʤ�D��BC����R��,�|�+�ɥ�x�$i�%�[+kB7����g���OYp����/�����:]�A[�7b�Y����-a�J�o>��<}�2�ܹmR��H��m�b����Ȳt��|�o�U�������4lӪ����f����� �F��s$�{1�K2�^��Ŋp������g��gk��]:���2�X�>؁�]%h�>���@�4,�K��!���v��cyOh�����RTv��8��M`�U��*[
�yw�
�i�Vh: ��5|.�BmҀ�����?�V�u=�u��nc��zu�ʟ9��PK$?�sݛl��!p��څ"�vi6��E<[&@�����i�L�� �,ݐ�����T8¥���5�Ս�����c4d_��R�b�R"$�Jp��x�����,�\s�T�o�[�|����N����ޒ�S���HoG�%���T��F����*e#\o�!?�l�V�]>�G�����X�����<�M]��p�d(Ǩތ�F�A�`\{[�����Mt�Uy�A���yD��G7�*=�H?�a�oΟo����8�PDmK#����&;���t`�N�G�.i�����8�I��B�U������[���z��ᾮ́X�@�$N���3����F��nI��4��ڃ��	����*W�!;.itS�e2ur���n�C����p	i����;�� �t��'M S��Z�<��R�/����C��jڙہţ���k%�4�C�@����~3  ;�Sm��1p>�E{��T�LD�_�����l.��[��U:)���ؾT�.��,9�� $�Y�<$7��BL�׹��gW�l��YtTȏ(4~T?�F���R��K�d�qW��GJ��T�k�B���~�:���$E�2V>՜�Z4P66 �Ѳ1�[u%��Q��y'w+�����{�2���e<�]��pNL��0F������� �����\��i��=��j��v���Fƺ	�F׺<l�����tj�V8�\���~|@1�P��뚿pVi��]ksT_�O�����K.7�h���{�8I��d�����5��OzRI2�2��c�@�Q(�0m-^U���p�K�O�� y��-Lp���n�������o߁�Z����!�_��;�* Cz� [Y�����˽�h0z�n�F�"�!�L�6`N(�VH�-�G	]���gI�۰$�#nZu�ѷچA�����f̖],E��A���wI���pSU��̱�[T�B�J��=`Y��� ��D:��H�Cw��<T��#+IW\�2�%"���>)m|W4,����xCuk~�t���{]t1l�����X֫�R�C����#!D��ď_�L�F@,����O���9 �7
Y��Cz4�*Fe�m-kh�5����.�́� ��>
�	��	o�����LS&x����\��fw���Z�˶�ډ�P���EN�Q�K.�h��&(z6�Ȝ�t%��\��EK_�&�8Ǔ뻖]�(��:x�ҽUO��;�&Z��.��KF^zˢ���+D�tA6^
���6ݳfYBU�Sp��nae:6:'��&�����2F�4��D���B�������ޚ2xpߣ�<G�����\���1J>�S�U�T~�E�i���.v�Jl�8G&;�:��ghr�B��$F�����_yhΆ���T������m+v��v	ے�Ɂ�ȕdXd�I]�D=
��J�$Gv\jF�<��[��@���P�N�o��Xe��R�%�&��@�*4��u>�4Y4I��?��g/�BE�[ZD�����l����H��/�N?�26|�����[�!Ú�[ r0���(�-�)�)}l�lu�;{^  ��u?�p(�w�c��m ��Ƅ�*]f��.Ʌ���-4���'д�!��p!'����1C�J�Ni�_-��J����^��v���暓�+�E3�@P z���`��j+8�YLZ	�aS�޻Q�j��hD�=�4�4U�/vσ\Lm���)R��/�D� �)�юxe�7��|�{q��p�����1o^#ᄜ�3;��W�\f?����4�F��������{��[���L(�pt�$�+c_]Cq�0�
�L�X�"���0�&AM�\��O�����ftZ{\ԃ�<o�л,)����]ΟݤݸZjKT@=�*Ѧ������jN4.�C��pk�?f:j���T`����V��Q�@��9=Ba�����?8�2\e����"ʩ٭+t� +��s�/ң
���R���]���.�/Ή|O�U�������=��J݊�*%��K�=�X�ʬf1��tyb(�,��L7@�[�q_�#l`�̍$+Rw��,�k NrYV]�z��~��N���}�U[5F�D ��:����H�^M{;[�JDe�A����| 6)�'��f
�wh�:5aҊ�q�6}h_�8�:����;�6s�*,��B��X�hB� Z��.�}ݗɢ� ���s6�!�*A��Х���jg!���i���J�-�q�3�J���t��/���)'���GH�D'��.����]��N%�0���&��9��I5�������K��bt*Gѽ.�/G7^��\����Og#ۅu-�<�%�#9���~�3��*��uL!���Ɛ_�yAq����$02ٴ9u o�2�!.�4�f�Q�~���}l��0�7�{�^�H��P���,�2B��:�QD���a�����-���>���A>���Ի��&��,�_�k�ހ<�b�����Ik9����}����wG��1^���Ǡ�V���w5
{F�x���H�
���s��e�D����-Ƚ�G���Y�Ko�/�����|�?�װ=SH��C_
��L�w
ų��NP�B��·��. #C5mϊQ\��V\�jy@�A���,r���*����Ɋ�;o�<�����za d����Z�oG;��x�Uc�˄�A�Dm�h�u���xHH�VQ�Ȗҁ3o�$pÏ��a�a�xNp�"����f)@�A��o�̶v=��(dKº9��0aZ'���X��J-R)(!4��T�q�PP!���<�$��YuR��F����m�8ĥ�}逃p���yP�1H����b��D4�o���m��W�ٵ8a;��/ ��!���̪������bq*pV��Ļ�A��j`�Y�QGv�0z�|����.e��"�S�tc|���ˠ��`}�4�r����3�lzk6Q1�)�ΈNSR�|�56gǘ�U�>�YG��6��9���U�{� X�ө�&��{�QJZ<v�_r�F7B�4�^~��c��#�GU! ��x[�.|�o��	�ljMr
�WHN�Y�\@N6֣T#��P�j�P�o9}t8N���u�H���)ڃ������f)�1�^"8R�H���r�U~5(`�;;9Ѓ�� �ƹN[���1�t�2��"I�˦B��)�Y�%�N^r��V^|!�ۨ�ʹs���Z�Stʁ�kC��K��|'�G62�vA��1��Z���B����C`����$6�0z��%�6�>���@G���{��?
�>���fr�V�nP���Hh)7�o&���SKY5��:�u�����}ŜH5��Z #{�� 5�.�����IӳY��3�,�F��s?�&ĝ�B'6�h�"�~Џ��oa/�-��@�s�?�� �"��p����Ӣ�s���?� ��C;��(���yql<�3D��-xPm���ny�=OS��[��)�+����I7ƌ�R4(`��J��P��P���KЋ�6�V� �4eR+�7h%uz�u9������gJ�`�)�� |t��� N�<&@���cv�_ʴZ^�gr�a�D�6��f�-\f։��^F�K��zX+����Ft�n��{��>(��	\��U 3v��u��^:ޞn��Y���9*����/(��@�a�ҍ>㛾�[�O�.%��Nj�K��n��C����{/�e�!RN�����9r�� ��B�7�n���	���"�W�$7������|�9>\��R>+rcݰL���qe�Tّ���T���$��X�4C��f�!hL'=6�03��)�PC"�`�
'�(���8?������A�� ���@̟T���Y�����|F$ݮC.;4��n~*{��i��=K���Gӆ;�Y����`h�~�ZX���&P���m]� ����>W�g���#���x�H�;+��a �����C\�uO}L�t�.�⪀Y�%v���::�亩C�R�ܓ�n���M�}Q��|�FA��@/L?�*��u@��$Ei$�G4�ňgSXt��H~�\s����� �3��ؔ�CJ`A�c�-4�(T��yg35�ʼXC�Dn�m�P�㜭ˤ��&p
w���\d���sr�z짳d�/z22��H�vD:��n*_=� ���.�2u���*�����n�����0�
Њ,���ɱ73�0L�.�ݓ�����#�e_$��Ŧl�V������?`�Ƙ�p���ٚ���s�$�lw�Ck/��7�s��;o}�rl���ra��識k��}�w�����<X���������@�(B�#=O�v]�� ��W�>���@��>� "��Hpu�2r���8$�D��#�?��"U�2o����eܘM���W!c/��[�E��)4a��ʲ";~KA�@�s��g~U��ߨ$��7�G)�,� �x��-�d��0&���쭾���/΀Y�%�}&����(�WL��a����N��U#��]t���D��,�D[E�CQ�3���f�0���pa-��f8��1�5nh�ؙ���ښ�W\�[[�Ɯ h��Ta�^��g�=��sψ���?R�]��d!it�et�l��b�ʓa��.�/�����	�����m�P��=/8y?�g�sm�ɗ���0�F'�X\�춿��U75�n�'�4�Kʦk���8���s����%��yɛ��7?Ia+��x[[��i�#i@4K�W�V��RvUvV�a .�]�ތ��ܡAs\��t������ ����9�����<:�v==d�ܵ�fe��uV܍4�[s~sJ�,8�3N�-ֻ5F��:-V�M�D��cpdς;y��9+��v�S�C1J��&Z0��@���U�����] ~M�7�uN!Q��聹E5���,����.̃w��C��k�	�ᗚr������FPj��H3frm���y���|��Ts�[�dg!ד6�"��t9���]��%D�)���)�ni���8�BX 糡�R/�#򡱸g����FN��rq���u��V�n��qR�N�AI[�d��d�.5���j	ބ�Uy)Mc�S��u�P��&�'����'J�=-�@�e����:����a GA@��_W���z]e��W\`���������r�F Tx����Ø��	�J�6+�Eob���� 6��q6�ض��I�k`a�����ǈ����dc��z��+r�߂�M)f�̹���T���J��zxr�=Bm̺Y=����.�}iE�^������q%�A��襍U�j��`K��& `�\Uƪ�p�*hC4�y� �<R4|�X IϬ�NO�?���C��"�Оw�bc�����:�i�*¨�;���7�8�!����'�P��c������S��[P����dD��ְ��i�R�T�� ��m�\_C5ȅ�G~�"�0�+�/��(���m8�;5h�أ�E_[�r��_dO&7�<�C%�AV��L:� ��g8�k��#�b�}_���Z�J��z�0 �0T��F�8�ᶓoPM��C[8?��|�T(f(���
��]<�v�C�lb�]�Ms�Ӡp�
��������n��'9�1�Qc�8+L�NG�ּ�P�[�k�2v�� ����^d��Ԧ.�Upe|`��9�8���-�~�~��7�&�W�i�����v3/q�����]�;u��F�H7���&F�}g�[�שc[n.�g�o }�iQ׮�3_�tKKd�8i$=�)#����wY����:���'�p�v�G���t&H�� cv�îGu�����;1��%s�b���dut��V-��G���ׂ<��{I�-�?���ȉ��p'��c�c��}��Mb��<UL��Y^̉ :�WPC0�r՞o��O���*�a<��$H(��k:Ć|R�j� ������s���线�����F��"�`�#z��1�[~ɔ�l�<E쳖e���W�̎pLFz��7~�u�=��ݴ�+���u���h��l�"C����x�� �Aל~Ñ�3�5�&����&���[�ē��~�;b�ى��'�a ���0�;f�]���8�-XcQV�k��)�J���hN���	3g����i���ٓ�M��ƦTyho�g82ŋ/��c�OM4�k7��:�k�I�I�T�(!�+3��W<�9-�ea�f�1��Mƛ�$��m�f�W�����n�5<�4�&�[��p
�6��L���Z{�[l���j�^#j����p�2,�"��W�� ���8���j\)��V	�=�D������#/dQ���������4A]�����ZFN8�#)G��+��)j�	o`[�0��xΰU9��ع���j4��SS���)�8-S�n`<ܫ��<~X�h�3U-b�vK����@&�52��&����N� ц�p��h0[��_,6���zw���`��5@��@qd���v�7cqI�佱V9�˄Z�)� 6`�`��.�}����A٥��7�'bVMmܯ��IFM����D��"ԭ ;�q�P<������鿽�%vՔE��-��N-v5����m�?$@�P��dt�]w��j�r�;"-��Vo&��H�g�v#n���$��K�:�V�0#�,���#>�Ҵ$���ג���5"�K��{�8h�2���f����m�ŏ\ło������=	�ȶLc؛%���1�%���UG�e��(�kC�=>>��;��?�O=��v�=捻b�j�;��Tg�\��!�S��;�)��)��O�g-ۭ��N���N���ןr���M�A�u&�����31�+�B����;.à|���n&�|����i��n�j@�d`V��0IH\����kH���vp���'/��k��(C$�a��N�dc/vN1fZ���-�)m+�LJ�pΣ> �I�Zq-H4�5����=x|�Fe��%�x�o������[�=`���O��.�����y�d;w>>}��Aϣ�3[$�+ls�؟z}K�����:��3�y�R�&oS��
g2rA'�(nH�mF#z5΀U/���r�8�>
�
�˚�&R=�*7��t�Gݟ�l��*��WC+G�Γ�j=�]7�}#�8��~ܹ�[�S���iTg�����aߗ&����1��1F�}+{�m$���$��q�i	N�Vpmxe>��~�&cp�U�ʩ�8��JW56�U��;TƳ��2T=C����m�V���瑭���"1�n�^��}&�N����R�%�b�;[�~L�&7K��^w��vӺ�[���(mٜ<W��Q�~1n; )N�8�+`��\���_�$<�b<��1'7ѽkP���L�k��`�
"�k����N&,-��Tb0���"#/�B��*������c�x��:�ۨ��,d��O2I��w���L���&�()���n�'��@�d�{��@����(V���� ����EBd"���b)�����΅b���c�qE =D�>�٬Ro CX�iar�G�?"+�*i4X�0e+�΢����t���[��w�c
��$1�3!��l�� M2�����p)�����␆̤��I���;	~x��O�\W�t�����k���������;�$٤�:+EWwM��N?�~js�#�"�</�p_�QK'�@&�4�u�3�4�F��$q�k0E1��ֶs�^�T��k{R��^�Vͧ%/C�\����ۂK��x��#o<po�tV�wl�@<JW�u��ҫ�����xN���avi����S���}@*��t����C�6{e;wjX���4�1߾<GK,�ܰ�D�����7O��.��\�3T�~��zi���P�-3��c
ߥnJ_�����xMY��(xFX�g��Uf�kbSB�����b��^���Ǝ�t�2��@�r���f�G��Ѕ�jo�g�)y}�VQ�~���.�0�����m�N��\�N�0�Ә�ZX`�ߎޤa���=%4d�D��Ԗ�ɚ����u[���%��qh��'_�{�Z�����9)^���u����>���z@W�a�B
��#�t����\�n�t^[�8���R��	ƲrO�f_��gOٔ�U�L`4�?0���)Q�%s�k�x�#�_
S����!K|��1��ԝ�23AG�8˜����
�E�BZY1]��Q:h�$�E�A��G�1�Z 썻#��s�xn�<�!��gIKT�,���}ZB�F�1�2F���>��["Λ/fg��EC��=�*0R�ڗ���L�d�$����U+�1<���8�U,�l��4�}�- ����Z�]�2_v�M'��!X:��Q^���>�{<
^���)?< 9���^�2}� 5b�Ǹ��P�!o}xC-���liy�=��V<�5bp�<b�c]�=��^D�}�J�Y�dl��&��h$���P�?���mA�R92K6U�;Po��4�� ��"����
m��a6�0`v]V}ܕf�/�kc�k]�%V��&y)s�5�':��D��d(C��X�]\>Q��c^�&�
ܶ�M�0LC2ҷ�F�|_����;`Ľ�[��1]R������_I�΋8i��u���[����૨�H-�H�u�5��!�)����2C��8Ao�4$$���u�a� T{��L Dj��9R|;vۀ<G��tZĹ��^-�\���s�nL��n��7�U` �t���H���L;�>�+1Eb��� &TȺ^���v.s׈�pN.�,D��>�q.Y�o�p�3#����"�Yݜ�]�hhj��V�aGJ��Ͼ���*�UI'��L��\@m'&�B��dP���N��;��xTߺ6=](P@��a�g��� ���XHR6�j�h��� ��*�S�"$M:�8;��݉�f�|��@5hES�2eg.��RU��GM=��](͠+HP���&����ೌ������Unl�額PIj�7�H�mp�Q&?���L]�:GX�I��Y���I	���QMp�m׈��b9��DŁ�FB�����do��A�a�a8�v��z��`��Yx���f�uL�$V��6���N˄X�%A��B�)�\�טgs�!��F�5���^C�������/���	����RT�\pA2�(�C��̽����~�V��{ȷ�V����@#���^�-���F�;�MȺ쌩5v���8ú	����2.������:�H:Q�1�����@��ܡ�:\�_ߊ�m����r�(�V�>7vS|0�#�����&L��9N{���ժKǕt��w��%�������m���^��
�.�����)!�F�\�I*�Q�L�&�v�1Xk���F�?17J�n8�zG	o�`e�2J�����\Q��E茢GV�6v���Ş�0&��ۺ/%E�n���3-�$H��������b�t��ī�uikT-D�E�e���Q��V��kMXq�R���RoY��CN`r�&$E����4�R�}��J�8ts-�k�!^�+������0��Wf���莾�v��˨#���J�$?A�Ѓ���gYu�w����.P!޽̉˗�.���Vx5�婽��?]f���&��a�O�J�ǡ��32��i�w��W�R��.�jEĕ�d}?�ђ&�h����s`�^�)&V4t���Џ�o��"�s)�z�.V�^�V���9��zr	��je�s��e��ı��R�KHjCl��'��ߕ`J܆qj��_`��^����q�|�ʣ���!;��Gu��A����y�Cw�9]�����ZY�L�\�%��i��f���	N��qRA��ﯥP}2��"=������5�2<��v����k2�y�H�Hh�vWs��ѷ�<3�(����Q���M��9�x���.���K��z�s�Ӏ�nq�-�5�[	u r�N׾.�)���C� �^�§����u���F��B3N#i �_��&�c=���2U-O�C�t� �F���|�^l�I��i+6�&�K�P�CK���r�g�Ũ@�ǽn9�x4�`͹�#�"F����Ũڊ�5l�ֳ0��\R_����@@�9"B�F-#vS��pu���1M̠���f�.���v~>�>�8��:�&\��dW5�$Yj8��' oH
ɨ1à���\�R07g��!�E�uZ��V�s�b<߁P���p���`f	u�L�i���_��a@�M���V�b�'`���3�'4O���_�9�ß��,-�yˎ��KQ���#�`EvH��#VbO	��Lb� ��N�
f\�e�L�Z��M�\���
iq������*0�/5�-�4��W`t�Z�=/j|gzwޅ�k>��d�#��.��[/�h.��꣎������
'�dh:m�v@������l���w砙����1JQ���u�.��o?����R��QG�Ɵ�}>u���ō��v��b����:[S:��G�O���0bҢp���4������Fnl����O�g�B��,G���;*�畆��W�T���ȟ`J�T9�5���c�s����#6�L$.�Gm<�U��[��
���h^O�o��'�W�����)F����lG��Rƭ��3nd1��Ȭ�B�Z���Q-�n�Ї��q��r4�ʣͤqpțҹ�j�j��Z��,� �mҋ�����:+2P$��bU��M��RB������7��7����9,ӏG��}T�t}k/���y�܋�#]�cnL�yNy>�W�}	��ߵ@ϲ,�7�hX����ܹ��a��c����.����cR��zC��_� �����0�k���Q���T}�:�Y)0"�Ge�`�XMB��I�z�
��`6�n	mR��2�)m��iX��B��փ�b�g��N���D򟀽�I�Y(	�	d��L�Ҫ\#�V�����g8,뢏����1�B�L1V�G(�h����`��j� Ε�������0x�N��9��C>{���)G5K�o�p�6k�'8����B{�S� �UC�D�� �=��uEpcI8�����}	>����+�XXX��d穊�rS���'Hp��7��!J�!Z���H��ɿ�)��̝�ǉ��lL"f^�Y�Ɗ_q��K�'�����	ta�W�ԥꙣ�qcpg�!ր���g��0m�� �!���'�,��å�A)���;��y��4�Y����E��6/�|�k���2�
���(X4]V�E�,V5Ex e�����l���'�!�N5(�Z�Lzr�Kq���8�
F�)�yaB�N��[ό�Ֆt���M\@8�`�H��`;��r���N �_,�^���Kx��_��e��Q/�,=���B����U�D�*���l���82,'�y�3_M
�S����_FL�����:��Z�`?繱-�?� U�nZ�>�!$�rz����
h'��eW�?S'�B2�#����N�Xp���y�c.��N�v!��ܧ(U� 0ȣ鍕_/���Kӡ�Y	�@0��NEV�d�/k�=�y=�MÊN�fd�h��bt�bcj/7m�����͕g,b��itpĊg�I�)��Hb����XH&�r�c��7Uđp�բ04>~e��	 ��aӋB��>: ��B�
����pM/�X�xߍc��~9s�j°�gcba�ύ�LHy59&���d5p�NR��r��IX}nf٥Cz��V�6T'z�6?�4Chu�x��'���8����5I�T^"�OG�{�$S��҅f7��-��J��t�zܚ��+�/�5��@SROMh�	I����hݲ{���2�4�P�1i�o'��}����y�RQd%~^sd�]#�VK�iGn���~����
f�;ϻ����ZU����i:R4{3�m`�Z�&�zN��H�\o�[P��>V)���5�)�������i���2�@;>���!or�
�M�l2�93�a��}+]5+��J~o�t`5r�M0LN�E���xF�K��|��'X������	��p���� ��"'�>�vbs��^ ��S��bz�S�#���%g�qa;���z��N� �e��G���ϰB:�� �2�=3(�R���{mV'���R�0��=�_�(��K5��*8>諮��!��d�����ā�R�q�l��� �&�;���K��	���>�w�9L���uZ�����BWO���zo�{p��Yʊő �%_0ID�B���d1_x�!�f���	���v�y��v¡�$PK .%+�Ȯi�$C?��mu������~e���bS���H;�t@\)	�m�ګ�I�U`��r(q��R�-\z�t$1m-�XN�.\ր�̦�!���X~}����GB{����L��Y@���]����bj����[b�A��[�w�V��:%]OE�}=z����dŐ��D�`�$�,+�ɂ)J�)R&X"^ʓ�)� h����0@<���2o$���D=���o�$�&6k�uih�zm�������k������a�]���/�(| f�%�D�?����������A��;⧷4�{���jQn�H�w�c�R��� X�@U[��0:�u��@s2m�ͨ�)=���t��C(	�S�Z���n�F�0,�N�c�h�ţ�G`_�#�1�m��yOg�R���o�d���ر���G����-S>f	���:u�NP����-��2�W�C�IG��@���e��A����ar2G���qR�3�H*�e��)�Z��:+_��Z"A`�{	V�O*몡�`�H����������>�K��6u���]��>ʹY��V���k�Y"o��i�	�vs�!�ߢT�֋h٥}�T�uJ�[�lrCA��H/��8>��>tcM���B�q;��DV6�֩��9 ������F�K��^��G@�HM��Y��t$/�=4�z����X~���ƍ�
��ÙbL�[��g>uCM�d>K��d�/��� ���4�Iv5�~���߃�	 ��:��\�I���u��h��QN���t8z�ȿ��B�gĻ���?j��G��p�����9�]������kAC���N\�T��Z����%Lb����-������2C�!܎en-�cygP��-lk�p`ȋ�>�h#�A�&��qT���Y�K�QǼc�4m.����X3� g'�:?�e���Ou�&��S�_;(b�B���¿�H���x?�I��}0솴��kI�l~�ׄ��q�2��'�6X8�Ҹ_���a�tj��&�X�P����|��<�ҺT/��l���2��*�[���<����l�bŪ�����.��ln���PWu�K�]�dn����pXF�{��e�z�L�S�����Z���*�f����A�0�@�`xy������Zs�N�6��Y��&R ����oK�6��!�*��@�D��t<ҥ�1/P�,K�w׍*;���]Jmk����m�5�Oj�O;�����Уq��l���=O~ӟ.`����P:4K�]����n�?@���C��Icg�k�e딭�2 ������N���dڛ‐�
�7##�I���K@��rK-sSyy�B����4y:�+��J֠���<�?l��!�߁˕�3sJ��P?J>I����o +��Y�N��k���`L+|��͝�T��3����J�s���m_���g�SEu{ O�.%dB?��T5"S��˷�湒�8g�� �4�	��J���!�\������IcL�H[ͷ*��g�`�c�u{�K(q�ӈ�xZX�[3�u��\y~8'	�Vq���|�.)AW��R�D��ؙ7@�e'�([M����PXqi�2�}�4���m�I�W(�"���΂Idu�1���y���u����<G1�pǢ���Z=s�1��D
ln��-9��� �A����L_cʦvSk�2&3S0 ��%��f��o��{��~�8��r�����X���5};��Y�L�8ea��ɴf"�&f��p��#k4#a� t0ح����9�V�B�`�Mv�����6؈��\�Y����-ｩ�#v�,ҹʸ/�N�D��Ő�<h�wF��Fj"��0�(����֬������R��b���{��X�H����Hk���7�TM���1�!��K�s�VfU�Yj�e�-�=�v: H%�G���U�B.��elQ�H'Y���`w��炐]�W����`Tol�H���nBtz?�@uv�^[���Iq��B�U�[vkh���h�c	I�د��5~�3pN��*�ң���.
�'KT.6��:u2E9d8B�՜�%C�w'�PT%��>��<q)���A!����%���b�(d�I�[}<075�T�(�x���I	?�R���/�[ۗ��3Y�&Q��>��m[��o}�c��>����b[�(�pc�4�#^�𭓰�͉@�Wb8�5�u{!�̅��Ԉ�Č	����̀��d�0)��/ 4�@�n�ک��/��M��>I �j� �=�т�>�*U@v�g؊N]�#��{-W��V^HEt�U�P(3�J]�~y��_^=w�$L<�k����Սꗛ(D󀠑����bZ|�[b�7��.U��2��f���
��x�&b ��;F���z��R�bl^���`n��/�H�s8��L)�%�Q������:���F���9K���-��кNW'3R�A�͔��)s�<�7�r�s}��!c y����W�|1��a6���GN��A��_��^ks��zm�eKeyH���f4��D���\��`e��wÌ�����-��~�����r�?��s�m9|��#6�����W��WfQ�p�lX� �G~�ѵ����^��x[�|-��XkC��!�M�=j��*��A~�|Q?3�����'�B��^�����&���ג��PT��и�޳�~�*�X�aǼ�G@[=��^�H����1Y|8���- ���W�ӛ۩�g��#��6��o�g�3��S�'�W�+�|��K}��Q+��RI�n=L�\'1���G�V��}�_�$� A;pV��
���ɂ=k��7�.��x��4����o]���H7�������F%�2�"�J�������Ɂ����7�W1��,�Pl����H����t�=uW^-���{E�Ft���[�#�gU���o|u�͓(�w4T@��r ����<���;����_�\���x/�tf
Ez �� �
�г�MD���e5�-7 K��4��%�O��4l�4ۉ��sI:�(߁^��?@�$h�~=��6�]G?��î���+��b!�QHi�6�Z�ȅP�a5����\G�Q�/�����{Y�G�8��5va]�
��9��}�إ�jr�@/��ҧ�ڐ����r��[E��ƈ&�/��О����Y.�'�n��3U��V!Y�&��n����{�h�X�(�����i�� ��&�|�f�}�Y>7�mn,p�N����3�K~��rj�x_�BvB���3���,疖�PXe0�9/���ٮ�/��������Y'����oa~frM�#�����M?��=�v��̦���Q�Uz�W���O��ī��q{� ���|���>#P�y�0�茳�oa��JM�C���Iw$w�#�*֡�)�N�v ���0b�{A�����~#��+\����Oo���8�+�Y�pU�*(]�����f���N�R��3k��e�Q�Q�[��[!��^��CT��yǦk*ط�z5��˴����A�z|/J;�gG��r��h�#p}R,ˇ?]�l��f
�8`A��vz�\�0'#�_�@�H���`AG�@��� Qb�3������.�266ڻ��N�<��V͕R��2r�i Z.��؂��`3���;1�d7���;�
I�⏒�Q�Z�	�>�#�/%1�
�#CC�$ׅ�__'z�0��Ӝi+5P������uf����&�݆�V�}Gr�ZOF
��dR�3�
ƚa����<�U����Ȗg&[L��gF��M�p;Qs@p�w�o	-��L�b�^K��ٰ#��A"�[�����$��*�����6l!�yA.�l+�MfLf�gT4{t�M.�ueO�(2�4��j��I虜���&�9�d��<��RJ��S`��cJN���Þ��4P�^�&��sG����Ou��H��z�[��y�KMVo��TPD7�b�I�y��X9]"e�J�(1��mB퇑��Fz=�'��I] '�|��D=m�2�6��}G���b�l��ۯ�@���[��'3� Vwd�?����
CKT�����Rx��<�Yu= *@s9�����l�-��q�o-�Y�f�z��QN�����n�>�ۚA���ǋ���-�M��~h�FE�0#{h��3л�l�d�K�pc1��`��n��)��{T��sOҭ��c?�؉��|(�`�e�|Dk'|�,Ù$��CTh?⨑�h���?�,h$�?�Ө��"m %������%����a�W�̩ZH�9�,X]ʘ�v���D=��.�?�Ж1BA��'�.�7���j��Z���wϑG�u�YK�V�B�ϳ�p�T����Yޮa����<,e�e��*��A�F��.�mp�M�C2-9^�wR�Eǳ+J%,k?��F���y��q���mϵ���6�jS��>K~��2/`��ޓ��5h��+��{Z�e<Y &)��0',�6 ��v��XB&�瞱L���+�v����ÂY��D� ���直�������wbuTj� 4�(�6f�sYJ�r0�N*n-�=��u��Ôg��5��#�T'����m�[%B��6a*G
�s�,�H�����o����Q�v���UO�ֵ�����!Uͱ�q�	���冘�S?[��ǈנ�ѿ��o�X�����aU,Q�{z�X�u���U-��H{$��%�3[�!�0��t���n�s�'��K�A���3���6�mmR�6��H�D��'�7J�Ǌ�&<~eB�����Q=�w�u���i���n�Z��p�B�#Z�B������{�V:����R-Y�}(��l٦XX�U=�]��hv�r��7��a���b�H�LE�=�+\��Ɫ!��dwj���7)3L=U���;�:���B�ܞ�-Y�~�f%�LAe�^^�B���NDk�'�LuLb�����3B����Z�E��<V�B���I�Μd�7Uv�d����4�G	¡���LDx�)��I��=�L���ۭq~�tۡ0$�f�N1|��#i�'
y,�*y����w�EV�)*��aq���S�G#fm�,�Z�_GF��<x��=K���k�`��<�,��ҥv��6�}yo���X�gʚKQ-~��fT�vYcd̩��Z����K����Uxz|֏����y���З[��8,��6��-�N��9�A��}F㘲ef%V&�+�.�՘����,){h4<��jô���w/�Qw���P��u)XA��+���*x�7��,u�h�`��oנ����q/DAц��
n��Z�V��ɪ�lq���	���Jߡ��흳������bz����e��G�$3��}3d�o/L')�n�C�)�60�S.E����C�3�k�"�CA��r���p�["@�x�,�^mA��!��ieL [0wZL(�n�rp�{B9.v{^�k�W'�� ��q"#/B~|!M{{�����ob]yM��ykw��6u(u8�(��þ�"�q#�wR칊�,?�Ư7��cNa#�I6�)�>vJ�wYP�*xZ���tj���X���y���:��vbD�D��R�IQJ	Z����.�%�2�~���1����k)�� a���9⮈b���	]ܴ�.�p�^ze��3�֤�I2�nt�~C)D�V�5�ݏ�y�����-\X�H��	/?s\0��4�Q�r1�k����8�jN�����r�O�?�(z��`��9��;������(x�SNm�;Kk�b#�zM<����b>���0Xl�P� �b�V5C��o|Xw:�J�ㅷ�m�iČ�Lu��1n�W�lucms��6(�
��.��d(�A
����n`S~ ���»7p�ʧ
����y��/�F��.A���2ZB�!��(`*_ӵ�a�g¾�p���թ1��I��4�#_v(����(�7��=��祔L%�1)<I2�G�i�{4�[JЖG�쟘��:+f>�p�]s�*e��˶������߻�����]�]�'/�&2]�j�m1Ih@��%)�]�ի�-��=�G2Hk�H)P�㊏�v^����P�Z/1d�2���V��̵�5F������:�F��tF�c�bfC�Rn�3u.�SY�k.ZZ�i�_�tC�dtO7�����C�qbr�h�"�ꜫ:����:��)W�H�� �O�(�ȟ�����+�'ȈZ.m���@6�����Ĩ�r���9�����W�b�Z��������n�'}��aQ��ss���UF���oa�X)� ��:��r�RF��v�n�ǟ����u�o�8�8U�u�14ve��_�;�P��7G*�(�J"W�����rGtk���휞h�{>
�=�qD7�+�pz�
t@h;��l�j��]�_���m�>͵�R��<:�9���kI��xP����º��ή��?T������*(���Rih��V�5�����
�nc9������p���"n���t��������@����c���|<b��f-ۉzou(�V(̗)iF�T�I�+܅d���-G	�V���=�0Mt�/&s�6
��B�%�kmR� e��RR�� �l�Q���Ȋ+t~���X�Z�y%�Fa��a�I}M-�pf���/$p%�����3%�c.��Ȩ�M*ݣ*u�zy���~:[����7zz3��f�/
�?2�:�;]B�k�3+_#8�s�@��g��*dO3qɿ3��'���Tstn�t�fX�kPȓ��a�[��>�,͍d~�񂵋O�U0�i�1s{��x!�i�ų^���3,�\�^ :I��Q?\�k�����U3�@�īq��uXz�*f�ԋ�v>!RJ�>�KBT͛�Ӷ���w��Z�	Upd��֫�_?���KI`AhPO�j|�;�p�2&Y�>J��0OÐK
�b���+�s������r�dhe؊��59ݖR7�j%䚪F"�u�c�'T����������(ۺ�V�cʁ��3������WkW^u��X�����V��ꧯ���=,_�"=��>���ю4"&C~F������S�.P-ƚu����v{�mqwΒ�{=4{y�}!��}�Am����:m+GB�B�C�PuJ[=u+Kq@�G 1���0u����V��,�,r7[�iK��3h��6.*�o����7��1��h<'�����
�4��6Y����K�AO`qP'wg�JǊ�b_������W����Cv>`urJ�QNwz`�ygZf�??J�4�x;Hd�YGU��������Ó��9��zܠ�_Gpi b/͑��/��"��f6�������)V����dm��� �K�4ѵ��_]9Y!'��X�409hl�R�tQG�S^Hy���כl���ϱ,O�>�p�^� ���Z�a�֠_֒s�8$tr���(.	k3�.wh0Q.��kZ��u��KBPi���Ug�FSVXcy�KQiǍ�ֽ�`vpӞ�c�ߐ� ���_�QE�[�#t�/��zZ��S�O�e}Fm�g-�3, K��]+$3$���_zJ�|���g�\^��M�U�	^��{h�f�ٴ�������Cd�w�q�?�V�������[_ ���&�t��%��s�@{R?�v�m�&��M��`�����1
�d]��t@n%���s	&�������t��.Ȱ��%�q�K"�i�ǜP=g�u�9����7��Ȥ� @�&�}ylpp�T%v>F#ǔp���<ݕ�ft�}UM���d~�094G�Bq߳9�r�\�V����۶!�Q/���H��#�n��V���_`,�`���y����u��)<�����Dr\�3�m�M(ؙK�`�p
���AZ5�]ũRP��BE�����`�v�Bi�˸B{%�P�>�H�Ԡ�{�dM)��d�|a1|��!�Qu!Q�k'�V�a��~��*Q��b��?.�͞�jZ�݂�
F*�6t%N���8���I�GY�-f'�	VH�g)���Jͬ�{ҲǍɿ+�#%ø"Q�T�v�۵Ѷ<q��lk��uc
I���sXa�#s|_���� ��P� 3���~��}L�n��iS`.=����5����j�]�ÈZ���}��U��r�$�h�����vp��\4�P{�V��XG��<دO�D#�룱����Qg�_�C �a�7���f+�1���@ۤ3&�z�D��/qw�Z5i��p�(WQ⁑������kώL0 �h�/$�Y�(}��4]�����@������K�P�FT0Qґ�B�f��5�#yQ�i�L�b��4Z�*��Un��?2����Us�� �9��b d%�B_��&\�H�vÏ�����ff�k�إJ_{@T���χ���Yd���7�<�h�_�g��b}>iZ��3M��	��&|�0,�̜��Z��P�1��|D�h3x��m�$��Ff�S�}���p���@��|~ ��z�\�#|~�7`s�r���K۽�miI��*�ڿ�g�~��~�M�f�y�:A�tt|�ڎ��ee�f��b�]0x;:з�,�F�vŅZ�r���+�: @jS�Z+���o����*}�L�9�)8�3�^kI��{zR�`ݾ� AL(������x��_vf	-Gd\���L�!Z�
d[dg�s��^j�_J]�#`N�������y�ċ�jƨ���}!��,=��u[4s���YY�pV�
��'Z
v��
ZEm�������ْ=���z�N����Q�$��"̨�����U��P�� �t�Z�*|a��A�����Q[*�'x�[�V��3@XurJ{v���D��d��DN�F60vLH �|⬮�h�3AE���B;ϙ#n�nr\6c��'�;vK��W<M�	�X��a|Т�bV�+F	�ɡ�;�TSV�'m���XHlN��V����W�q-��n�%��q]gC�!w��]`7�A�[x��;�~%�a�0�#�N��F]�$�M [�x��g	Xuo�]��5�W�(+�W4�j�=�����6,��)��̧/"ݩCQ��Q�3�sy��~�5��4�D��J�t"�ah�Th$�vR��L]r"�0&�ηa"��3��M��e£��~������-�*C\́?���T�I�H��8o1�0.�I?�DE���4K�8�SɉS���Md0𴃦6i���"_fG��u���i-�ӆfIRu�*�e�Yu��s'�����.YX;��L��*�K7J-�QE�n��I����9���p -�P��{�v�E����S%��vz�������)�0�_�� VQ�B��0��9��C�
��J��(.V_|B"�G3v��N��Z����o0�Rp��p̈́N�K�v4d���
��W�����_#&N;�j�H R"����c��	�U�=,*�"�$�w��\囦���5� 
Xq�jɟ!��	v���v4����Y. ��\LC�9�NO���8gd�����c#D�12x�z'�Cd��X�g>X�FJ��4�jS��┢if��!>�w	�ɽ�^y�:*��4������?>vz&b�v3�J}%����a��8*DՃ����蜬�!�Q+F q#�˕%=lo�{��@'p�{�X�O��|0�ݦ�笡��{�~�8Qd�<�a��� B+���H���2�
�5���	��|.{�*G�m�;4�������ee:u�}=˦�3`�n�Fś�ZCJP�;���:�I����"��4*�%ȫj��Q��q9Ў�C]`:�ʝ��
�M��[	��5�+ �b��"��6�:�]��Ne����gkT������d�}K�����`�	��(׌�U��l}p�|il<�@�9T�ڹB����4,+��ʸቚC*66:�	�&���wާ.�0o�)�O�Na�m�J�'s�;�
C�Z6��U�������"���V=j@#�*��krH�Ѩ�BK>x�r���)���"��	�c�tC?�Z{]h~��ڳ5@\��C�t
��eQD��*�����y�ғ-ϸ}:��d�V�F{���L"b�|5PX����ְ����i�����5lC�>i�&٢�~�T�����
R;�t�ӯͷ�"�Us�(S��������47L���X��q��0��x�����US��67yb�����u���8Ѩ�O��r�eP'<�k��ǚ��zZhF5�$�(r+�=���z���uj�9�C4��PӰhpް�!H�{��ݟ�J��4�O�RV<�xҴM)�W�9���%��oU��cf�GN�<qv(/�y6�i�9V�"�:�n�y�V��$j�gVH+b\N�u��r���ߗS*�l�R�>	e�Y�"F���9��dˏ�u�C�]��ms7�^�I��$$ �;�;�i�p �z����=�eL��c��R��z�t��dQ��O�(�|F���R�^�+g��Q��
�dK;��\�C�a�ń(*��%ζ	� �-�9ݏ�M3P�q��;��-q:��k?�*���a�t����e�22�@.ʒ��oV�/π��k���
nȜ��̭TU<��@�����2�N!�r��8��0
Fi��$�)��-O����v�anVp&���0iP�r����٣�E�'q�^�ӧ���I��>��nQM�/;ϥXV��Q��C�� V�5~Q�T��$���8�N� ���i�����l��2�؆m��;.!��}����&��Z�x��IA��͐�؂�sf&����(�Kv�����VF�71�v��*.�`�.*2�Sq�i�y`�}ۮ�+�Iro���FJ<w���,[4�2�8�@aÅ5��N3P�H=��v�f��L��Z�)@�D�Q���ߘ����%�-*6ˡ&�(�^�����'_Me�@1���h��F���0�%R�|��T�(�a��B�5*#�4�����rK68r�D]�AKD�>��q�}�uh+3H����a�ǯT废5���r��!y��IF'آD�B�ҩڽ
�;u�ARA���t�N;��{@�fw��:�)���,k�Uߛ0�Nrܙ@��e��lKǮ������fP�ւ�[Rh��H���F��{n��ؙ��f( �·��R",���q.�.'>nx������o.��R�Zû��*0,��c	)��.Y%�p&G7���"ô����ec�[� 3����)	���H����&��z�f�ˬ�� Že�y ��~���/�Џs��~sv��|	~{p��~7�16G���{4�j� �'Q��<x� 9��)L*b˙_qw��!Yc�px�hLʢ�e,�k%ߎd���"�ѝO����C��<�G�O���2��H���_��=�*@��#$��7EM�?�����%4���kkê�*��V(x]��7������_����Ј�2 ���7$������"�q�;|�Wp��%rֆ-%E��`YA��[���+�E*0�,��qR��>Q��լ��|�L�O�cͪ�F���Y�3Az�IF?h߰����:����������v���sv���;l셁ޙ��U���i9N����l`����{��mx�,�f��#p�`�c)r����u��&*��II��)����Tk����oH�hHVMe�rD�T2���B����蚙�>��7��r���DBD�YB(���{�F�/H���p�R��J�+�V
�[��O�ן��#����0ֈ�FؤU$_���spgJ��^���
��֡9�*�U_{�s*<���:�1�1����P~G��Z7��W�2m���M�"c�q��8��u�;3f�]�U��e0ĕg�� ��6�X��ޓ�ǳ��O�vz��EZ�)K�E����V8*µ�;ed�s��������ʒ>}ð"�&�w�g|M9�-�x.���?�I�j�*�.�t��-[�$���nJ
��·�\5f�U
2T�c郧i�M��/`�B`�*�~ߐ�P~�[���p���f�i�T&)>4w0��}#V���4̒�lMY�*!+�<�c?T�x����6u��ظg5��w���&y�1��γL{�����"���|����B.0�BْTSA(��jԻ�yB:myށ��Y�D��ŔE�Vw���56����@�z�/8J9�
�5��8:�p+�-r�f��?�@PȢfk�S�(����a�
D�ӷ�y ��\m�����+^(�m�y6'ڏc��X�#��XLL��Qe����Zb
8\#B|{)�xq��}�Б:!��pۑ >��ڸR|�3ض|QSZH�j� L
?�jzbO:3q�>Wd�7�hTԳ�ڡH�v����рO���q���'1�]�q��R��O4J-��.Dm�� ,��s��#�Tݐ��;�,S�]��V�n�w�_e~0�����>��`��fJ}���W�h�������J�����}r{1f���5!��� �B�Ng�"�G×�܇c.-1�+�'���j��^]K�j�������ݾ�G��]����߰(�%��u�pEh�����Wb���H*����^�8S.�j�T2�+�Ŝ�{fywإf@��H��ý+��|ۀ��
k��B�?�@��}WX�qa0r7U)O�B��!P�y�z�])�8�N��ʿ[E}h[@\й9.tmx���9(D9�?W(Yw�֋v�D�:x.҅ 
%�������Z�8��<޵2O'������t��U%ci)�{|�� �ĵ��������=X���j��[l�Ʈ��Z�٤�p��_�'S�n-��t*�TQ�����Ί�K�J�uF��<qT��{��s�S�eZv7�QT�^ϻW^y�&(S����D���=�Wd�ﱴ>�?�E��<a�Zm�_JB-��I�R�E����2z�P41Q��0�_��-I��N� s��IE��&����U�� 6�OK{_&�"���x�87\��87w��c�|F��3�:�������d��QPS��N�����vk>�8<k $0Wy"f�� M�	��V#/Vo�|�s)!uC��;,�5DL�o��r���Lķ��h�*��MHõ@q(�9)x�l߷��g!�T�����%����IE���'Iԥ[H�"�Jc�++���/8�cȮe�P����Y惏�Ю\�I�Ey��ԯ1��;MѮz��Wdf�v4~!������ҲPqW�׏���Rp�48*�*g�}��`�?-�@-����ׄa�YP6O{6_��烻!�����k<>&�=CS�iw���Z�=z��%���*x:�jvFjW�=�D��x����:}Y�:�(}��R���c�(&<Ά��<Ϋ�nY���{B;�L��K�xy�3|��֕L�=���K�5�'�6�3����Lw��%�80��4:�;m���{-�4��jU�۫�[D����/��O�(�+X�d�g��x[�N�"i��Q�WL����2������3'���e2Xbp��>�!l����z� ���V'b &����}��WF2�G�U�?����N���V/%D1���O�[��{��*�LU�b�E�p��~&�m���Q���0�#p��_�f��摻T�{�N�����!����[Q�)c���L�o�����`ꊣSڠ�ϲ�%-9j�'EPp�o�<ea��+v�3�xaM����F;��u\6ҥe�ן��"�S�b-�����5i��nW:�S�i�64��d!����f"�-������鰄�H�^=��T֡��㰲��E{t�VX���]$�iľ�@$�.{eH��'�$���@e)�v����h5BǇZ�v�y�v7�H�mK*��Yic��v,�m<ڈ����̅t���.�A�t�������Ov���#������nm�Aχ;3KtT*�3~eC#ع��������8�
*����
.k�.���P�;�lF���O��XQ<%e%�l�.C�p �_��u��\��Z�b�ɑXm�=��K�&
f���(�,X	IdM�M���I+p������^�z��tJ�s�0���|����������	,_т/`�z*`�p�hP����c`d��3oF��I��L ��<�\��X�9�ݨ��Dw�,�u�����?�Z���u�ph�T3h�%�p���Uy��Fh�WثpB�U����i���3oV�'�9���\�H��FrS��u�[%�D*�Z���jM��绊��o��Մ#�#��O�
�ؚ���Je{����F����C����}�c_�z���������?�pL\��x��j����8���:��J�8���?5H-�%y��v~d�G:5��-��~^oj]�a��(})u~����+��(&N����2z�v� �2!i�Z�ĳ+w��o�>^��5���Ї�>��o��̂��H��A�#����ϮH��Z|��w������]�Lk<�a3���������ޤm��pKی��M[/��W��wRe�� ���M ,>ɜ�ep�uo'���Ea�CG�w�f�Ũr�==z`��Ԧe{����h�G^*/9��xα80n$e�4�NN�o_����p%���f��_
 ��Ƕp�f��#���u���M�bf�� ㇣���C0t0U}Ԕ�������u@��1BU�)�$�����&4-AR�-���|u��:��x[�n˱��|�9Oi���p�1c�:5�=� `E.���A� ���p�rl�e�[�	��5H���&f�+�����[�\�$H|�4���;2n�l`b�D�[9�u�+��TǺ�%gqRS˖�90v���K���>#&��X��Ǐ�Ǥ����Ev�C�e������5aM*��	~˖�i�	6�O*�;��@^�DA�c�	$�t�~���� �����W%OX��t�3���V�m5-FsZ�^_8i4��6Z]�5V�K�xT�� �VV���;g_�#`S�Xc�ߦ�zV�,W���Ntd����KK^��;��t
 �����.�^j�����9�hA���ٱ�����j�P
m�H�
x �w`��q���F�Cay$No�+4���m9f&�jGmW(X$	���F��a$�w�̫˫̪\��>t��1-�2�kM�G#X��[��Eo��AL�6t�\	�S3p�㜥�Q� t�����x�ZL�O,v�+HP�Ve�]sO��K�lr��"[��yu� 솃�+��;\K8� �(��HZb峻}I�Ӡp�{��dm��n
�3R��5��f��z.���G�T3�������E���m7U��@�4t�Ω���d�h�id��,��݀������5`G V�
F���y�l��%(|b��W� �C���0��9V/�̀��$1f�=
��MܤP���Ƒ8[��d2�-�uϲuga�x�A;����Ǡ���y�8���)@�$�Þ���&V"�:�Q�]�4�&4�`v���Ydةb��a EJپ�,��1��.%IQ.�Ͼ�~���-�csjĺq�x8�Z�"�s]�]0�C���]@� g�|BI-���e��׮_���|������1��_v3S�S�-Q�:���.\�'c[ü��Ha+�/���o� "��.��&(��@zU�;���gh���.�_`�6C����voݷ����=������ w��4�Ȓ��du��	~����䂝sG'u7���m�9�A��Ez8 ���쒯f�����S������\uD��60���r���3��q�B<����F�|��䄳G�x��#����*$ajN������Xw�F�'�[��+1��>��)D�	~�%5O��.x5��L��[���W���Y����oU�$�m�b�F�"&�{�R�=��q/A��9�v@t�m��R̰��Uj���O�~>��b���Xh��4Lo#�ИD�>�z]��]6{3���n1���DW����!N���:�y���=ݘ+x���QF��\~�PzL&�|;�p(�=�&nHbO�Oa��h|�.'����1@�=ənH�I�F�U����ϙ��M�Za$n����8�U&p��G�i���|���2��6'�!��b�iS֛��;�M��PH8�(�yeF��]�}�������פ0ݯ(�v%2�ڽ̅{�c%p�*S��N�(	b�<Џ�Z(F�r��_�sP*o<���P��g���`����?�8�Xzh��� ������Ҋ�x��A'L�K�37ʘ�(���i�qd"�Vd"-D֎ʓ��)�m��H���`8�q5���1t���X���S��<���~Q�o���W}Ѭ*��9�<
�@%�� l�r�O~�����%�����p� m�x�{z��݊^���2�V�kA�H���_���W nj���̽�e�}��?v^�_]c��"*��b�\� 	�-LŰ��J�_���
9����*ʪ�w���o��W-'mp�0FƇ��`��QT� �,DO_b�@�yA�|+�f��#GWk����]��2S�d=��3WS葄�o!33̚�M�����~�_IKF��w˪CT�dN��S��^��FfOyMيl�6��Ez��c<�Ө���RS���L�����U��xbzk�2�ސ�����v4Vځ�tD���j��q �Y��+Kf���ǻ��,�rC`�	Pz�~>�0���j������^��d���������W�.F�Z���(�֖�+6������)r�3`V�<��UHzMYX��|�u��\�j �thc@����,$-]����c�?��Ib ْ��r�u�q�枂�)���6�{������z�E�n�x�mpD�f<J��6��f�u{�.���5���h�k��	}ub���jk���n�9�E�����F��w{kr9R��M	;h�'̺|"�"��Ǽҏ�#� �& ��wp�W�g�Ѥ��C;��)-�V�
я��88���� ��@�vC���w.�\����ڭ���Z�;@�j[9&�']7�-�:�}4~洼�`�~�
��Bp�(�W��u�-�����TY#�ٹ&��O�=�c���.��	k�.�Ő8H�
ee�z����ǁ`Z��t�Ce��S��M�_�E����E�5W�c��y"WIz(�؞ѝ�#�����.]�Q_O��{@����k��3��b1�?��փ��he�6�a��UhdU"F26�-r�d�u$�e�to��1�Il�ʴ��1��&JmG*�`]NEM�r��)�ش�F�\L�]�oX�v�䮙���.�X�*���ei1t��Y�>?=�N�*9�����V���+����k�=j�%��;��(�ڄ�p� ��e��+�`��|7S���nt��>w�$qT���vUo��|؜7�O��	�<ͨ��"��+tQO �"�;�Ȥe����a�A���3Q]�6T�n����x��a�}")�%�j���^#S��=�D��	k��1T��N9t�@;裸�����٦�>i�|��)��d�y�G9{'3�Q`1���#�|� B�[�Q���n��f�&YF�#�W�~� �Nz}w��jB��;��%�l�u��mW�ئ�M{��Le���S��L'j.#Ӈ�J�jk���X[��BÞ�9DȬ��$CN���K�W�.4^;*��}�����Չs�}ds��!�ͫ~�<QӿI�{�>#��2w" �:z4L1�IX��� �I-Fsl.({bU'%�56�W���T�Y����>*3���{-H�g���%!�T�|">/5�/o'�t���:�����f-6�F=�v�[f�����	�%Y���Y�8���m?�R��?��؎�J��JJB�N	յb=Q��.��h���f�_Ɇ%8��.0*qG�~�z�A�v����v^I�^��G?.G^A�#<��-|�|��q%1�#�K�j�x'���1t�d>�Ӱ�ҝ^Ç�bS��-��
�^��c����$�JzArL�w#��)��ɺqăk�T6ߡ[�ZҲ#sC�X�$>����X�����:��7��|�B7��~�h�N?5�X�J	��b���$QB�}m��#%(���"W��3�&���
׾���,h�!�C��VR�����v雬��z����(�Ԛ�������7v�"��)�MQ���
Q�t_����4Y�q'I'u��wYI�xá~��I��t�TM��!�Y[7����i�(d���ti�ܞ��<�4���/DՕ�h!��0���P��yB��|���}Nn��}޹ɕ~R�Q���~�0i�G@��WS�Q߇欴�{}������m��ĉ�7��}"�,�fI���M���~ک3����D1�ew�	����򌺡	��8¹�c�`9<�a���v��N3���hjj#�"�D>����Ӟ����.�p�Q�pQ���r%\.r��^�e=E��´S��c�r��>猸8�2�G�1<SKα���Ʒ���Ų�mZ+ʙ�q�pM���XU5 ?Kn~�6*��ת�������t/�UJ��?q�H=< ����~�î�1t{U�?�%����'[��'4���3�QV)�nq)i;�5C�ա���2[�f|��n�Sh���Z,h �`ߛH���5w��Q��)qrI"��c�{����ux�����)Uʳu��2���o��hI�l(fۜ����Eſ��B���&�X⛔AJ]���)_r�T٢L�x���z�v�YF��LE7��].��UHt�S=܅D~LH���Ύgy��E��v�^�[[<�@<�����)���O���ҩ<��60v㭠j��YqUQ�R���~�_G��\E�c@�7��H��'�DGp|U��u��O4?^HѺ�m�"�GnZa��M��g��;��AY���z�iɧ��-�^�>�Yyi�i��Y�
!�˺P"��g���Ȭ MW�@p�Ky}�n+���P"_��{�XX��Z�����(Ac�t_f����k�H5�>f�qOa-t�1Hg�Wb w\�-m8�\O<ٔ)���������3�\K��2��f{�6�91��Bpzo.�H����o�P��a���2^�`�F�A�5zޤ����5�ǥe�ȉ�]8��oӴ�I��g�$)!�=k�6�X�;� P��0�)-+�9n���9S9,AJ��F=�s��>�,Κ	���E}f.w���P,|T��0F�AC5�� ��81d���+�Х<���Z��L?K�9"�Y?�,�\���&��3���~�]$����쉑03:hJ��U�+��e#�*� ����������&�h�3������r�2k@Z2k���
u,`���� \�&�A�mf�:l
�^Jah���s��Yk>O2I�~U�*%�A�g����?��0�,OC�E��x�[��m��s�A��4	]V<e0dcP�T����F!K�0��0,o���E�{�Dc�P2��j�C#�+����"4[�
u����qD��~.M2Г��-y*&�|��(.Q��Ҩ��߷߰���εU�zM-�|t�\s�ث�1�1Ar��`�M@4˔��٬�6����h���P��ʰ!�5���~� UE�Uɩ��3	�����dMںcmy!=����ae���7���Lly����Z&�vi��d���G��]ͦ�����j%L �Ip�춉2�r�4�ŝ���Tw)"����Y4>4�@6<��j�����ef�c0>t��(�f#�ў����%�0L�Ⱥk���������W��L�¨N��+��"���~�[�ݙ)�nx�<>��Sh�̌�����(���4�V��� ��@�C��Gp�|�V0	<+���g�I��������n���QXq��xT���P?��s�ܗƝ����'Y�q��q��uFt������ �e¥w@�2f�}�k� �՟[h��P�QkŤ��\=I��"�bI$��@_&�O������:�qǾ�؛P�~:е�ej1����(��2_�����.j���('���M��p{��{���ѥ�����7�(�A�;`� ���ތ���jig9̢0g�Q6 �t��ᔩ�
^©���;�����>HTC�,�P?"��{�����w���#�1tF��;)k�h��!u��{Z�$Y]`�)m{������fr�O��V{f?�u�Jk�N1<i��\s��E#�V��Â��~͉������/X�]�_��i�2����&��K���j�u�0���Tc�#��E�&=���7 ���A�O���H'/ɓ���k)� ����lVjx��a_^�諈��R��/ Z��$?Ĺ�.u
�� K<N �R����j���K���a�pᖲS]�q|\2���s:qu��q�Y�z�Zv%s�cN�Ɗ�5���w}�����6-�(��(��/Q�2(I;b�ߔXu���nU9"���1}>!��������t�ڙ$�2�ˀʎ��[,#>w���n|�o��9 ����ok�upI���C�6�Z��bl���iߧ�! a��ŕ&[^sTh��k��e�hAhA3���H�� 
$Ѽ�޾����;�9)1�������w)(rӸQ-'V�7�/7J�v@Ӓ��٦�v&��.�\u���W>�~Ȋ���!e�k�®�Ry��Cc;`fZ�j�����X,���_��V-�81�W?�ˡ"��tk�t8�~#ܼ�aMj.��*��68��f��ߧ-������GM|��$y�]vB�­�B�h{N=��?eP��AQ�Ѧ#�Q��� b'Wd���Q���߈��ô��)L����o�I.�_7vƻ#�On$А�K�� K� �@{�z�����<��{�����[X��v��4nsEt
�C]��6&"�/���i��2�ѣ��{+���/}U(�KJ����%%����G9���1�Z�郎9_�`{�}C�bg��֌���-q&_$�z���8��V%\�34#���vf��I>�Yy�eH$���
!=3�v8g}����_V����+c�[Pa~8��>�ED��p����O�H�;���X0��b|亮�'Cfb�����P���y�HT,�����@a�wű=6�ҩla���O��j[��x�����Le�;�@p�J�s *W��QjD�NZ��չ?���mS����t\w�5^y�f1s���6��_��&���×5����I�bRN-����I`r|��V3Gy�U�Kw�0�q�T�)x��Nc8�-O��7ޯWl�[���h ���n�:����~z��d��['���B*�O�H-�6���������z�Vf�T6�	D���.��sP��� "�j�fC�����D��8��F]݌@���-��g�y�"�e؏R�v�cYB:�|θ��V�<" �qԯLB�g��������B�OL/�VJ�)U���+� F��� D�V�*sA��3+��=7�D
N�j����.;��}�/�W�ǅ������B�9S��4� �[F6��qxK/�i&��N���1%�#��M�%x���;��ny��m�Qr�'@@<i)�b��}b�b↥�W��
%��)`p����/cqB^���KD���D�W�I�+�Z��?��8�`�(�P�.|����ȁx��8ɾ�5��I�U���b��,$W�fP{jx��2�����q�,����^�����ϫ"���o�t��1��� ��玘P�Wv�ASMӗ�j��}�^l��7���̆s�k��
X<���{#�z����P�9��?�)�E �=/cX�7��ܤ2��c��#̡�"=��C�zE��<��C	X��^�o[[���&������S�'�ݨ'�p�[�E��LMT'�����ӂ�^�YȬӋ�1$�3��@U�L�y��-N�`5!4

/���6$��v��(��nl��h�5��2�:��,3[� �Oz$5�`N��t�~��;����{�$:�H��6~��0�H���rq�i`����iD5��a&��g�S��4*�P1���H;4��\xk�O��K8X����%��7��5u�h�'�1CI
4t믭m*��yu��}�U���0=ɹ fM��̅}�pRS�¦���	:t\$&7pd�t:>쉧�_���Z���Z̷i*�ӽ4lj�iX=DYs�!)Չ��烉9���7~l����I���(YA�h ���fqq�c�g����W�ù�35<��9�ry44�����	Q��[$(%�[q@���c�"h�/�2s��֥G�w�lV�Kфk��X�6#:�����2���-�e�2��0��������~h�}�&˥���B�.Ov)����% ��_�1����c��\������jke[?�j(r��^�7���r-5�Loҕ��Ώ�\�!Kɽ�㓨xZ�b6�Zcz����F�Jg���q����&w52��5�"�-@���7��e�l|�1zJY6^��85���ش�礬'Y)?\Sm�/��H�/��̫i-�?��WY޾�� ̞:��r]2O��/O*��9'09<f�2I�	-?�ȿ�E���H���b4-?�M���Ru@��u���K�����X�d�'�z��Xjr5�%���B*��?)H�~3�~���85Hz]���БM?�}Z�	��RH���/S�~,.!��R"M�2�*Q
]�� ђ����7U�<���]���
��S�B�#�ǔ���J�����z�LnCN��j����b�Wʠ��$=C��N��>�X�{u�؀-��d<�%�aF�
���[Iꈧ�L�2y�qXTĈRw�45����z 5m�)�����f�ڡ��H���W�T�����ae�I�γD܇�Y���m}�Y�\�7O�7��������"b�B���~���,L��[�&����� �������aҽ1�ze#����`����9�H��)��/��a�>��m���t�цuzDbT���E���`7��?	�{>]���nB��Z��h�{��'!�EIZ;�`�jy�K���H%�z���Zظ���	Z��{�,,���p���K�lAt����5��_p���Y��^ȃA�ʰ0�mc������Z��h�4J���=9d+��1����=����V��7IfwGBʰ���><�}�١��]��N���5YT����5V�"~�jֿ��P��8�1��̹�=���`�E��pqf���tPg�����-Hb~j��SD*l�\�ؚB�Fe�nƺcB��#:��I�x�	���9�,�m�����h(����~�|ini�IwM[`\v�>�'���2������+��BpCzcX1P��w���}%�Ιc�P�Q��X���J����M,`���>l��ɚ�B�)�T8<����;%�I���ߚ
o瀐oՒ��OLa��T��Դ*[P|.��|-`T�W�f�r����E�ss�:��8!q���;	o@Wv������l�R1H����
��n橑35s��b���^�h��{�������j�z��@�3�a�`-3$��4S��$7[#qs�wKO{�(hE�]+�Tp�Y�-��KJ���7lB��
p���)�,1��L�}<�Nvd��&����诮��ja� "OT�'-��b�Qv��w�R3ТƓN�Ut�u0z{;��zTǆsj��'�G�(NN]{�������?�~c�V��4��K��4����Lك͘Ew��>�p�?B�.�X8����繊��bq���U=��~�@�[	�==Di��|���q���qi^��C�!~gI��3�O�\�PN�9l≁�d�V$��ݣ;ߦK@	dO�("�V9�²�!��J�[@^'-�`�	����,�|�0��i��P��w#`�آK����.P��/y?���@���z�#�`�l� LM�=��r��4挧�� ��Ƕbd�-/����{"%�P�ʣϞg�� .AU�˷&�FIj�ȹ���F��{�5mI�	��/~2r���x)3N�Y;��7 �J�͊�ڿ�'@lz)�Ԉl�K�*1���^U�X8C�f���;'�6�xm)���c���{��K�d�W�E^�1�G5���������K �&�"*W��6�z�jL<����R��J�x�>sq���f=�p�vgL��ǖ7��o����G8׹A���Ohn�T|H�+��qa��4���E !x5Vvns j����W9�L�u�I�woR������E�d���U��4R�DH�/W@\�=I�fqi�G�^�j�Nlc�?}�w�$��y�Z[MԎ%FB����Z�(袎;�놬�U����*�G�ݗJ��0פ��D[�FZ6��ѥ�����݁hj0��ٴR�Alcq�}����ͮs�S"� k��`#w��hb�����N^!p!N٘%���U.X��Aڤ��X��:� �\p D���u7��G�=I��� �L!�Y((��U�Y��U-�D"�14��P���BS��z�#akL������[칮�ZJHD�(�G�� �W}2�ސb� ;Q���ԇ��d>��1s��:�W�������E�����Z^�<P�$w����fU$fp�dѲ���R�?�HtS�u�-q��b��;y_��	���)V��9A�²7�QU��j�-�<�{�X@J�{��u�1�\^u�l�#��:�f���@&J�<&��Q\�T�[Wz�iL�
j�|�K=�E*\�ܵ2�EeuyM����H5�m�c�s Ex؋s<0/�=��]�<D`(CC���/�AA}V}���s|������6��+R�ҳ�Lz�8��#�%Aq�����:�#��re��y�
O
�������V=HDӂSjX�\�k]�����Kn�O���;���v��(��[:�N�L(C/� 2b���&8;�J)�����W���={
��3�6CE�X����T�&~`R��!���]���N��� ��)?g�u��wE�tD�Ϳ~͈�Z�I��,���f��R��D��K|�f�/#����*3��c�j�Q����`�e�Y�.�)V���| ��q�@���J��⾲�l�wSt���!j���g��ۄn�����3��!��\H�@�$j��V[�W�3�����1��wzӉQ�����5�a=��~���6AΘ�˳��-�rx)���+�V֧��nvTA�WP�u�$8�>��#x�h��Yx>��[�U�	8����t*�;��p=l�����m��Vf���������L�N��v����w:�vӸ�B���ⴶ��҈�E�-����`l�q�(�ߙ3�XЕ6���/��[3ʿ���M���ŏm<�r�_����>k���f�@�e�K���-�K�i��$2tj����݅�Ia�+	��ҳ$Α�8%���Mf�ɽo���)I�H�����7=�]��吖�m-]�"벉zs��ݮ�p����fGY.������۵]Q�nV{N��A��w��3g�t;aG��k�'����� �C�O8�]�|�8r̭�%��+��&	����Mu�>�;�(�QOL�V"O3���5������!�m�t��1�� z�����5c���[��F�n9�pD�9e�Z"Z?��	�@�{�NԺX4/I����F��KgX�.���E)'oB&��QMx��^��nxa�tF�X鑑B�����N%�3��Vq��2�)�{4`����,$���9��Av9��F�� ��%b߲�c6�F	�`�E�$����&��܏�-G����-L ��0q\;ۋ���lap7�R�ϫ~|fDVJ�v��u�%���>�:�����uRt��-pO���� �Y�+f��N@�0�7�Ab����mQ��9e��h�b�rK[�'L�.+��0<o�x�v�1:���(�5�f��V��&̊ϒ����ö�YǾg�1píi��nqA-���x�)&zbD�M���8Щ�D@�/��ⷫva�g��pZ�c�����Q�@^v�
�M.�bF�|?��w~Q���)�,lA1a1d
Z�D!#ʔҜ����F� L������bd���(���H�,�;�GTh�$ӡVA8�M�M����̍8�\�IGp���d�=M\�u(����ZH�0Ydxe�
,��v����(z��=q ^sە�}[3s�2��C���UX�[ƌ!���j �]�Q�J)=/��j���Y�]�I��Pͯo��[&5_�SZWtD��c3�,�Z*'QG=z��\p���%����+�*�c}��DɌ[s��i=q]v�[��@o�z��7n��Al�kPgL#:i$Wȉf�i��s.w.��޶³���S�L�I��ǳ%A���:}��z%	}���*a���)�ޑ���P��:� \!6Uֈ[�Nb9��{�l_��%�L��:TM4o0I�:��@/C�.@͉w������!�s�0��AA�W�[lZ��1�O���:�I��}-Z�<�#F��{uaHs$������k����צK{�K\҉�p�J�H'��E.�s��
�Id��x ƨœ���a����}�W���e3�+��¾�:��mї0qh9QM�9�"rJ/.[J�k��'��U8��;�ÉG_�؈�X�S��zyA�Hބv��κ��'=�r��iq��q?/�����$�|�y*<gWe�饸a�ɓ�nJ3��K��B3�|Ȁ���zX�7 �zPh�anQ���o�����������NR��ϯ8��g���mQG�_^�P�{�]
���A�K5RQ�����@��q���3���i0���*�!��ʱ~�}#}T���O�(d��wۛEGq����uq�I�ˏ��E�]�+��MJ�ReEڣ�ɴ�;��������G�Asܡ�
ݡst������1��<.����������A<?�!�x�t֐l���v�'D�́�`�U�P`i������&�~2����L���Pޥb��ַ3Q�S,V	f֞�K�̨�b�0ϴܤ개^�8�R�"�M�î�t򜣍��P�,릁P@�b�U?��ㅁ�/�7�Ь�0�n��Pv���]8��gԣ�ʵ�+n�g�?��S�o��d�8��%���r@G�����S�tSwFs�L�r�`*g�B�����a���>߁Z��A��p��jFz���!�W��������e���Cq�κU����M�S`s�C�=��q,�>�G���=�Pρ� �ЕF��ʭ1+ه��d/���ـ�!r�t� =���ﾾ;�Ng�C�v7��^~+�c�ϰ���ܢP�z4k���e��&���x��S\+1h�m��f9x@�(ߞ���FK�Ӎ�-H+ʍ�;�8lmhp�7����*[ȫ�h�]�|��C�Iu�K;�=,wA����e"= {w����-���#���V_Z�O�3TQc\$�'@ؙ[q���x����@Q�S�l]�֥�.��^4���5��H��K
���Q���y9�r|���vw�8zn�e���D?���))�c�N�W�(�n�w�Fh���\a��>p5�U/�Q����T튝nѠMz�����f�}��o�o��� $���{.?Nr�f��]�(��2�����ȏ�I������_eKr�9�[d�5	��mz�Nə�6�&����Y/=���z#�����tZ�����bGi�����3�-�����j��L����V�wY�)=qֶ�(sX�/�n�g�=��>�Ej�C�UX�c�;2�N�ؑ��<�p�ӹ�8��k��x����A�!���u{�p1�/�5�,!�ɔ��³��8,�/�D!o�^�8e���i�l���aF��p��%fڨ;.~�Y��Ҧt�#����Hqظ��b��k�	��¡�X�i�$���I���vÍ4����v�$i�%�2�L�
μ+��X##�B�Kقj�O�_{�{���R�
8:^���-#>~2�2I\��vD���1@�tӞ0�e�=���Y��g�Ӡ�CSk�?�_��IHzͨ��E��t�n��Sw4�;�}(�y�fMe��}6�P�W�k@7���Y.��P\��l"�q��LU��X�2H^��s��v�iY��� �}�j�A6j�z��K݀.&��c}�I�t��H�\<������G�e������4��,��F���M�W&ЉT[���~$#��7sBi�������[q�H3����N�K�ǉ�H�C�f:P�P1��)y��OiJ���:�+C+�i��-�����nLU�Q�N��%��L���� E6�Y��������"�Sv.P	���*�H>�P�EQ=?�?!�7�^Wh��+�G���:%)�k<�gI�<��j�O� �%���ܻ~�y�����e��$�dQ����Y4z�e@?c�tM����s���dh��Ѓy�1K� �!ma�� ����F��@&B� 8,�j���%����i_ e�
r.og��4i^tS���@�����4p��u��O�P�\⴦�~1�`�<ޖ�5m��RSw��P��b�U�,�/�Eyi�yf�8��ҥ��h4#����EA0��C؀��w��o�/���AIg >�W�)��C��؉9��c-�}bj˔���r^�*���w�Yr�J�l%��> N낦�(Y��󐐅�겮b�?���!�4���*�z��җG��02��+�t����fˎ,�w��8�b��c		r.װB
�J�/�-�2b�~U���
d�V�ї�~�U*T"g�Q�p.dTY����ε��]ߝ��*�D�8�:�`^QcQκC׍]W�u$aU���G�I6�g�m޵��Ҝ	�o֤�w]Q(1�y�Y��S��)�`8��A}���鞵��FC��� 1�e�{����Ф�,�و�Б2 �&x�����jw ����3��yw�.��q�{.�Ԣv�ǧIƎ������@��� ���09u~q��F�c��)Z"�[4�	?xB�l�g���,d�W}
�@M2���!!G�H�ua�ۋ��8����ɷi�3��ɐ�v��r���n�U7����kV���F��,0��D�j܊�[��d��I\�aq���)�V:á�v0���M��h	�s]�6q�E�j�i6��e��h2�:����T.���
kV�#�ݷ�,Nx�g��P��n�e/��@1���0�h�kS��ڝ-I��L� ��XPH��[�,��.r=���+�蛓��;Q�ˉ\H�&,g�!By��
���� c_�k�-t���kT2���w駢Wh��[{���LׅeJ�m��B�c���$�[��y����9�����0o���H��
�B��f<���u�%M�֍�NA�+T��-3��J�S @R��"�,Ƕ��������ZN��;Pv0�\�S�Lp���F�i�-?���B�b�'O�F�|,�R	`9�t[R)�v�Q����8!R/�1�����n�?�`��K���[B>_XC}Ɨ�,������Y�'(]���^fI��g\ɺɠ�3B�� <�s�u��[y���(,F�S���SU�(��!�Ur"�~�NUJ��[��,�?���G"b�a�HPc>Mm`�Y��,�m���7�54N��%Ѵg�|*A���c��Gw�5��q�	ܬJ�`F�a�Ī�Ly��|r�O��1�����-��I+�C}�b��R<�ɝrBϫ�H۔k���~��	��8�3De��kJ�e&2�ӞV�`�ȗKs�]��&��x,������H{�#�5"���"�����h��<���ͬ{�w��ө����>�ac�:/ͬWN���oճ�/�%�����K��,�Q<����	t]a>,T��r�^'��c��Z�-�P7rv�H:�ݍ����"�&���M�̨�J��^�j���A�<X��3�I��zuգ�¹�|mO�οL7��>�^���� E����?��#uj85�o��1-h�~����d��c#@�Mq: ���S~�`��#��`�n-Ac�X9���a�@�;������Ly��P��ε���ϥ>��wQ��ӻ����<%��2 ���꟧��1 ubR��@��]gs8�"՞��n�F,��S*Mn��q�3��#���u}�9�BJ�j\�����+"U���/˸��J�c|��u�% u��:m��?�*շԾb��L*'��E^�X�㏾�����+���X+b\�As���>�Λ�	g��l<v�%x#�t�@rMY�̧U���q�������~��;�����˵��m?�fl�����8N�Fh�����ʇ��j��x�7q~�l�n�_s>o�a3p�n䚮8���?�a�hd���m-�N�V�}�̎�|�=�<j~�V1�l'+E Fi){~�����;��}�kUK�bi���lOE���L��uw�j�&8�n/+��t00)z���^VC�+�-V������+����OԿH=���|J"���)$�3���
72�/���V�oGR����B�u��Էw�}94�Ã��Z A�c����	Ƴp���o͒��^����kG�&&S�tj�s5�h���P��Ԃ�������Xzm�eʋvZ���ؓ"'��vt]0�[䀉���#��k�G���0>��\�9omw���13u6FW����2���*Rr�󉇸���r�\���Y>�t��J��BX���*t����(�q�pB΁m��p[|��1���.gң�i/zŘ���yR�"Q��+�V���1�!#W踀��� ����
��x�$֠c��s���?�{�A��:jȍ�h?�?��,J�[i�LǶ[8��Gd��Y0���Ci!X*=�"���ʼf��$�\���1^{?ܷ�4zW�R�{��fQo��i�C�@���$��CK�oq(����Ѻ�v#+���Ȃ��2��~��bxc�i�W����B����Ã�k��h>�>���^�Kw�����r�Z�2��}؍AɜKe��ĭ����3n����o��n_0�()-���Ϗ�����0�v�M`ņ��`���J�6�6e��8�yᮀvyh5¯f�K�j]	�����[����5�u�;8�Y)�)9�-\z z����c�J�͟S(����\��5J��Mh�w�>���}��@1��iMV@�y�_�"�<łb��ļ@Ii<��<ϒ"� 晖��ٜ)��1�
)��� ͹+w������n��W�.�5,�Co��f�v0<ƈy�#� OY���HW���O�j��1�����`��8.�E��b�z(uc@9#�:7��k|���l/1
��x���1��?�`
mw�2곪�]>/{�����<�Z�֣�p��_t� �W�Ůuk`����˙� �Fu&F�|ڎ�?4°pO���}��5	G�\15DaN�9�Cɽ߀jc�R&� g�G�i��
sj��w=���5��p��j<9�	}m�.P����П�ll��5crӒ�%m��x@�"���y����@	�%5����Y�]�TC��*Wᨙm�F���<UTI$rL®I����F�a:s�N��.��9<�*vAٟ�wi�2�sKi6A<1�!���B�Ri3�=w���	T�[y���doqvBG�����4l� �W�%mH�)=N�T�;�d�(0�n��q��)���]v�[�H�iz���G��,.�D��8ܘ0�3{���S���-q�;�����b����D��D���� 5�2%�̛��g����9�d���T\���m������M'!�LIQ'U��Y��k;(��"˔6ζaEC�+	Lp_�	2YmM=q��͍oF�F)W�A����y�V�׿fH�����o��z�p�.i���������O��lև4��7�N>ġ@`�#;@G�P厁��Tl�&�8�l��F�����I4�*���ƈF��a��uEQ��m(���e-��,��q
6W�۬+X�H��h\�W�����虺K���M��9�J�൞��R�O:^��+�Ԍ�@����t���	R��>�e�F�\Ѩ$�p�,f
��4ޗ������_�F��٠�%�K!nʙiBa2R�/]������ >}����})���36Q9���MM.<'�s��q;^��4�g��_��2�鎟�sBY�>�9�����F����+�������Z�`�Д���h(�S��U�;��N����K��kM��m�=4��ob"�?:S�X.�;=z	�*$��X�7�B�4�`NP ��cOX�LZH�/�ް���G0?�����(	�D�"��h8٪����>�)�3���AKa�n����8'�f4Ϭ�5�v>�F�I�j�����Uv�����^�����¬�*Xz�^7X�F��2������/������1�P�8��M3u}k��ק)���=���<klF�W��1?At��j����%3s��+�Iy~y��z�X$���%}T��c"KT�� JwD��|
��%-�⿦.'
�4p���eQ�Ъ���v��P�ta��Eu�.h~ �����O�?�,��g���&��XUF��"0�8��A*�@�A�'%���AJA� υ[W[�cd��R�@s���҇h�w���=V|f~-Z�$���.k����\���Ԛ��x]��.,x}k~|�.�[��gO�Ԉ�=��ݲW��p�K�Y(OEH�r|j�c	�pO����=�h��ۜc���l�
ǮВ�, bY�O� ��>k����8+T��60��3P)D=#d"�w�NI4S1�z6�f����ԕw�<�,vp6$���)��f�}�w�]����s��纶ڀcp�{a�	q�$�Z���ެ��DF�)Ww3�(�*f����$*U��z{vx1������1��y��+���73Md& ��q�؆��9�%Qjo����i4Qm�|�N�@,s�|�Pڧ�q��s��6��)��Ƨ��bޘ�a�ޒ_(C'�8rg"ϗ_Sد&޽�U@@r������l�?'�^�¾�z���vl�H�Ɩʓ�U6�_��I��ڙ��h��Y����*rL�b	B�� �cņѿД"]y/~��S�c�b�d59Ֆ�Sc�4�N!��k#nӁh��Ƒ��Oc]Pp��<dY��_�ā�TK�wZ@8�����	V-a��]~��uoܪ�v<_4����,�Z�^��%+P��&jy���4)s�\}2Tn���Hw�����<�h�j�헲[C�Lĉ�ׯ��tt��P�S��ОZ���8�%�^n@fG-�lH9R3Z�,,��ﵱ)^k�)X�r
N�ܖ�����$h�E�n�дf�@@����NKE��!a)�P�^{kH���p8<~|Zo&���9\h�
�AM�ɘ�'�����:E��&�x��o��xB�=�qi���Y��A��)))P�0ҁ�'�)��.NFxQ�D��@j�:˼gP�p���=�ǽ��i��˗���a�"r�q�&��K��<�0/�v�s�ӽ����]T��B9g�����G����ć��Q��{�]�F.�kqk@�ɴ�>��W����[���N(0YBy*��'�GAVT������|��)�y*k�Z����
ӝ��gӳ����/�:���񸁉s`/�a��#h�����z���{��)��%�{;2^�W{������:����	d捥���q���Қ�c��ye�?���k7�,��ٺ"SN=�N��b�d���!
 F���Z|\:R�[�b�u�?�S��C֢��$��_}�]jA5˛� ��_~��@��}�]�6�E�Β����@y���"DbV���B+L֖ Mp��a���8n�?�V�n�Jǲw@���Uar��{�+�:T}C5z���ϖb����&��BJ�X��3���|d��x�v�;X":�)�T�|��T�JV˓�Q�K�Hl�\�O \y�>]Z�	�,>�yv4T=���]�� ��9�We$7b�:�F��b�ˣ��B�޷�n��������ء��>���a9&-A�˹N�Q�5���ႅ"�\s?�d%��v8!k���!�j�}]���ʼdT�{I�I�C�u�(!<
h���,È��-j�5�8�A�|Cl�>�9���
����H�xz��qB��R��.
HB>�V�U�:�@�b���:�{���Qd��$�1��4dE�鱔����x_�~�I�6��L�Jjjq���k���\W� 5#y���-��_p��h0�%�_�|�t�n`��|�NU ���j��B�V9������9����p��"2�@�Nkۊ���p�Ҽz�ɗE���o,�ʥ��BT8E��׾2'��@ī��Q��V��;W�����Hs]�X�%�k6���:X���%^���F�X�d3H̢[)鋘�ؠٸ�����Z�je]�{��K.�/�w{Y8�w,"�{iK5���P�@��Swld��X���5&��!&F2	a�3��	3�R���8����������e��~j7V/�c��_1�
%K�0�}�82(]��uN��#�N��a���y��Ś|�!"�j��
���x��VS�^\��߬�� s����!0
6	�|{9�\h�wi-�C�h��a~2�$TmC�����:����z��Rd��.���d��ʇ��@?L�/�;k�y+�7��M�K�K$"P4HiVM���/�+�Ũe���F�~�!,R�0�jGg$T	�\Bo(��ը3І��w�m��e��[1�o�l9�iC���� DC�MS�ֺ2���,�0���.~�G�G�B������j��2�������k�Oj���J�2�w�C�Ҹc�zN6TV�|�j��rm�͹"�EA�rj���
i� B�g}�Q1Hw��Y*�(�{�6*Yh��rK�Z|��-�$(�k�O�; ns)��r:��������J�Ū��5B�Wxh��;'и���T�]��JV�1S��Mw�6P�Tx��#8�*��rS.��#+ꎶY��\?�{�F�o��a= ՘�����MU\�.9��W�<|�~�z7�B��ovh2���~�%��V̓���'ٓd e����J��7IOن ^%X�F`v�Xn|7�7V�w���^���4au��D���1�����m���1����[Ӭ$���`��1�m�L���nu��M���l�o��lYۘ���J�4��h͐ r+bh}L=�s�"����	�߷HIӿ���7���y�PLb'e������E?�1L����LOa��x�I9w-�\cJ�L$I�¼�^5�Hu�|C2�6ɮ?y 
H�N�Ooe�$]�G��c��W�'��Յ�d������\����R����8�N����MFP���`�0�u`ڼ4@����3e���d� �b	� ܢ��?$��!"ۻ3Fx�M�>�p���4��H�`dY�������1^z��-޸�K�5@�����!�����a�4�kl烧����δ戺m�D�`�����i9�Y������R����s�5`\���]�3d<B�����W��1��� �̎8�c���Z`%i��M�i�����IQo���C*T$
���Qq��1�g��M� ��Yr�����S�-;��f#!�����Bc�25Chb	���--/�U��\�����RWH銼���b{f 8���]��ُo�Ex��ϋ୽��l^�&bY6!��r<��pX:��k�pl�x��X ��<�]`@��oo+OO�Tia�鋋��̹�E��,(�p��h�&��=d���������h>̵B�c��7D��o���<��uC0�g�Hn���,�X���&��륯u�[���M��>t,��kqGćkO2ޡO3�F�$��vK�T���<EY�`A�Y~�}I�����1�*�TXb����oч��'d�� �
��E�2�I�cq5�Av�{7(!c�+�ׂ>�~�h�0�YgU�sk;O;��{�D$4��ke��i�?{�^G-	����é�e�I�!�w��wQ&�3��V=�oLfg���f��� �ZG~<6:9ȇ!s[��}:��啁�t�� ��Ge�''���;m�+[������RA@�Xa�G� 	��8�@���( ���F����c����	p	(r��$����6؁����V��lg;qP^�ҧ��b��+�-�w�y="�XV���	Nѥ$���!S�6�KAp>6P�+�ɽ�w΂L g�}U_(�<X�R:�4=�榍�IN���H�O71�b��R�~�M�r̟ΣD��ل�)������%�g�V�)$����ĤЙ�3�&�t���c\9��`��3�[�;TEr#�e�R
�WU�`�r��w.
D����ݾ2�Lw�4q���5P�F����'�ͬ�[hS��Lr��G�>��,)az�Y"���Ry�| �L���ѱ�ݨ�hCm'�#޼F�=��|�YZ@l%����[�ؕ%;�܁���]�"�Ho�Es�ġ>G�@�c����E����=��a��Ck�Hۋ	K
@�f���o}ޗU��mV�D�usa��	+��^wR�z��$o􀙅�Ln(����*�/ת���*�F�{����'�w���N�=�a�������9K5�?�F��L�Ϸ�Q@�0��jR7e������R��ɺ�N����)MQ�,���v��J�Ny��+��i`�����"��L������q3�����a ��sHdk�ऽ�PҠe��R��)p܏���	DB�N�Ģn����:U�&�e�~>4V�,��f�(�c�B'a	�1��a��� �AE<|��ޑƇëN���4���� � �Xc^�]H8 ��.��#���e4���|4��?=�1��5-Ⴔ4겪"
2�e����T~���>���(��)��J�$Ul��:w���& h+��ע��^#w�.� �R�,��M��eh���G����{��w�1�<k��f�ĺs��O ]�ЈXNCW���O������|���L���'V��Hԝ�̖ �3��^�]�e��0�87�+hN3�b8C�$$n��֌�p��Z�U�@uF�g�lw���)_����_�z�t���)��U
���.��$ߋ]�� �JIr٨j��*�B�q����V�7�\��u=��DM.��`�d�A241 ����T��#w��ʋk4;%*�����*�$��[c2�0f���+R��4�_�l?M� �Y�;��
��\׶j���2?h���h
&
��Ôv��_e�w�Z'�U��k��2���Tg/�2�'���I����Ŀ=�������j���q<_b�.�ZZL9�Γ��=�,�a��Rv!�c#��*j������C�y��@`N��hvl�]\��m�X��js��R t�1`<a��MD\.�0��]��Lnt!�#�!<�<b�Y�<F�m�I���$.�?2v9H�mQV�������x�Y���,@��¯}Z�q?�[�{�ȉFד��yiL�,�N(L�* ���0+1Jբ�97���V��<Є{�T��
�#o'ꭌ�����T�nq���Ɲ�}�q<�C`��+�a�̊ÖW#���~�K)>Z}6&"F�"�0U�	P<�m����������6��������yt�6�h�~Bcˆi�6sÔ���YN���-� ;�� �j�	�ddx>�O��E�C�F�%^�q��T��;�NUP?2�{Bmd=��E�M�3$�ޖ�TpVa����=I�y�?��ٛ��!=w��	�|����%@�Ur;��"Aw�N�+��P���u��үQ$�ӺZ��DLe��EI��N_��,&2�e"o�.OMM(��]�)4����|�E���|�74ǽ�xT�TOޝ�9�i1E|��-���.!�/[��Z�}T��	d��x*�ƤA����YMB,Keψ�����o8f,��Ř�
{��Y��ƞ�@�ۗ<��.ɂ�w��F> ����B� ���~�}ce�%��OQ'(Iڥ�,lЁ��s�
7=��������m�Vb5a2���ZY�#�{��VB�ɠ�L-"�q🆩:3�ct]BIs}�M��k��C�3v�ſ��y��E���#��{v6��L���:2ܢ����󸇨�� Fɿ-&�2�ch
&t������X�ܗ ��(h\�SЫË�B��^��]HO�m�F�/������3���Y"�<�n�ʛ R]uu.{\S�?��&g���m����b���Z}�%n�L��u�L̌�E����?f�6h��>��ܚ�!�F�@^�$z;�+:��$%�8|�=u9ÏT�����yrQu>�S2�A&�F����4|ӫHK�JL�	����V�����D�h�k��w�`2�PU[[�vuS����ЪI�?�H���졎b5��p;rm�|�yDu:)}�}i�+R9�Uc��^Ǽ����%�K�҈�@��+�
jޘ����P�ݹ�S� ���°ee�(����!G�+�q��4%��J�lYI����шz����u�!?�� �+d�$|P���総�B/����s+���m0�!#�x�2��Mq�h���Nl!/ȶ?�]\�����'��Y�XS�j�������.p��!z�L�-a2x�tkB�s�rT�Dq�O���S������K�������K�
5�<C|q9'RR�DPW����ۑH�'
���I}�+��:�"�4΁��3L6A� ���	�}��3�3�Ī�5;G�HR��',,�Z!�x=�8�>�� ������7�6}nH^<̎�c��f�5ެ���s;�#LN��H���1
����]D8�A���u)�����#�-�2�r�åס��R���`��%�&�I>u��Q�1�!Y�n�ը�j�ry�|��a��3�f+Kk�z��Ϝ���'By���P �����Ϳ9����-{N�˜�"������^��s5F2��,XD<S�n���'�C�E������������CG�jFL*�� �������3P�� z�	�0@?�W!�t˲ܾ9�X"@����o�y��䊐P��tv���(4������{��߈&�vBsE-��2� ��
���ckh±͛�X8��=8�D�L����+N�qWri�	
MP�|AS�����M�x�đ�ëi;� Q�*t�n�ȭ�u���O"�ʜo�#��Q�3W!W�dj�UGU!�W���]�$�F�l��}۶>�=�A~�v'�+-t�tG�iBj����c�W`U�	�аGś�V���5'�đ�L�j�ݣW�U]>�s��W)�N�w�k����5;>R���(�#���@�K���խ����T�_s�	n�*8��L�~�-�}��gp7���U��h�a�æ���r4�*� ZJ�0[X�_��~�++y<G;~f�py�i�_��/]͆�P�K�	"4�����߮ܜ��w��}Dll��u���jv[�>F�·T���9�[!�ՑM��OYv�Q�"W���[���c���j@o�O��n�	H�DB}в1���5��1%��^~7G/�?HD���ҽ8:-�uP��M��/�k���~.b�P�Z�^3�`�R-E�&��J^�ǎjt��5N�����أC�s|�$5B���q��_ФK̂[�x��)� ���U��5?��l�Et�X^�gᒖ�bu$��A�:�8}Tqd�@�	Cו�t��"R/6�<%�$K�ū"�~�^�>Jb�ۣ�&H!��<�Lv|�zn	T5����x���r�UC/�j�a�J�ϠFt[ó���v8a׋��vM��ʐ�Ǎ����~rГ�9J��{�i`G�m�qc��d�L�c�uI�;���i�H1 �2&RG����)��{�>tD_��Z�2]���Q6C��ig~�'P !�*��S)��cC"��4�T�����z�(�� B�g"�NtOg��2�tb;��Pf,]k�;�t��τ�4�FT�y��5C��{oʊY�J�X)Y? �X7���}���%��'��6�����yI��jș�W�Q���k����]u{�/� �.�p��`8�>t`߂B-X/�T��
��Y�AC3����u��$zuN[�w}q�j�H��ߜ=P����t\��i`���e�!�p��v"yL�������G�=˵꓎��3�����o �)8�N��86wgE<���%Xn �Z����Cb�HU��Kyn��*�7�����.�KmCj��G4�p����O����DC��MJ��h��K�֗,�k����u
����2lqJ���]ں'p'5Ro!l�\�uj��<s����>[=9T��[�x���*�k+Z0;�Ů��g�a2&�Z��j8�b���UlEI����D��V1���S��{i��d�n���BY��k����Ž081[��6ĺqi��E �mvGU����S�#^���Z���s��a[�֠6I��e1�x%��k���U�+�uB�_��Q�#��]�F�k�M@/���Nu��TR�R�<s�`��b֗���Y��(�&���楮-Y������.�zdlh�8���2�75�����r���{�!K{�Q��vL-Bh�{���.�h2��K��+�6��/j
CQ�)W}H��S��[���B%�r����5�q�:��I�*�����XLM�����щ)�}��ŝ��o����V�z&uE�o��2��=����X����^�כQ���ʉ�Z�'�c�M��;�$Ҵ�5Ǆ��^�py��)��I:Ǣ���)֠l �#�T�(^�6�K�x�뭍��	�z������r<w��gG�T�)4C��o!v:1�U�tl�\Q̰uc߱(b���u�u�2d�Y��ͭ�*a��v4Cyu��/p��ԼPE�.�p��6a�k:�&v^�5��ڍ�&�?^��nhnd�E�YH4US�,T�! R�B�<pc���
z��l��c�{(Oy��m�����d,.k�A�N���c��ʞ�#2]{��9bR�g�h �i�Ζ�����B���S��d?4*��+ �~�Ƞ�Z�4��>�o��ѥ��r��c3��m/���-�e�$S#lƽ�۸F���r� ���{��b�M0" �~`�`Ď���O�M�j0/��.舟�E \��JJ��U�H꣋��ȺRP���p���YT����|����������9�S���𦨠
�|,���I���  ؏�#�,���{���鑽4��zr/#���8�o�B����j���0���u�&9��N��A�q>(���2�dԧ�i[X^�2m2ץ�lƔA�ё�dHa�YB--��T&�F��ː��(���f�D�BiGob���X&�����رݍy�����C�k��}{�"���z��ˈ��S�i�������ך�䷬zn�!L��M�m� .�<��;�QM�
fsn$S\����O�-�5En�#�M�s�&MbT��oª�н�]�;�"����f���M�/_,�F�������F�����`����I�������=ӿ) +��n�J�������۝\�/`/���k�)��3�]T�b�:�dO�y�� ����޸�P�RPg�����盿�r��ɕ6��un��F��WaI*���u<6�1�Y8�iS/j>7��go���_�7��[1+����V�]UVn|�@!ǥ:|eNV��|�d��W�>�}�K�[�ѡ&���,`����$�Kb���!�Rl��[q�P���Y���$�'վ�@^������H.82���U�J8��l!Y[0.۳�le��+�1c<B��G%� �@���D��WsЉ�:����������P�{N�=��.���ɴ��@��Pp�W�p׀���E_��"o�m�>UC���S�l{�}�!�h�<D_�hY���G��d������~G}0�����-;v�0��ag��������=z��@�I@��I9���ULhU�*����t�/�0�=L�{8їh�n�7�I1DQJ�Inϫ���/����DH�����kl��h���F�'����N��q�e�A�,��I|E׏g=��P��(С���f�S��̕��P�*�LS'g����T��u����T�F���+��~?v�S	\qi��yx�ȴ��6�$/��"+��դ����\�H'd���oz��q�^�D�Vtf�`��B\g�gsA�V��v�J�ҟnF��Pו�X�������������x���{�ŀM�M�{��$Z����;�����X�ƀ��e�v���l&�CHŭ���>�~i��^�H)Ȩ.��4wf�������I�W����O�I���bQb��x�T�UnN�|��JD��?KTl�2�p��bF��g�E���^D���N�\O�� e6%h.���B��$i����� �Jz'Zܜ��G�؀��협��!P���YǍx�cn��?3 ��1*%S��!��I�3�@��eݫ,S��j���:��Ơ������r����W�v7�V{戈@��^�8%����q�:_ʷkp�ot�ОZ|yX�u�x����:g�[kٰ�
��/N��mk�>�~-׃r���8��TQ�RE�-�I���?�o���Lߍ�������-���Eu�(끁0s� �d&>k��������$g��T�lV�I��t{�,k_�Yj��Nk*��g�̿�¥��P�T�,uV�Ό��Y��=�ϒsU���Ā������Z\t
���A��� �q�P��H�r�!������3&��A�Cc���Y�?djg��}H�d�{"%J�L��D^�[b^�"�u�C�8��#���v �){e؄��S��R�5� ��n�n1=$*����)d2|c�/����|L퉬�f�W�q=d��ca��۔��K
lr�ݶ��l)2�l�reQ���M����Y۞<�닼w���a�o�������vqF��i�wF�y�aOs�����&��������J/�wb'm����8�`Txr�õ��^(�dfqN�Pv����^4~Y��rDx��'�����ֆ�{J�v��H !G�&KO��Rr�5����kN�+���*喓B�Q��O����e'�̵�,j���g��5�;�[�v��
-�q�4|�t�0� O��,�4��ݛ_���|ݹ��'S�U�Z�=-?b�emW��cb�@����4s���KD�Z4�l
�R9�u���k���e�ԭ��H��e�f�\1f3�3�;�@���cF�Ǌ�o8cq����Oφ�;-J4��d�I�],�1ً���*��U`28RsGj������*�;�A(�Vq��7��Q4U�op$o�� \��@�4�T��{�v#h��(��	c��i��ɤ�2�N}��Ѓ�{p#L��wy:r��Ȳ|��AG.�K��/�p��)�q�m���Oq��*�>��e��`(#�(ͳ�����ze�#����2S�J ���WfF���m��7�]tH�h�f:���&�&��VFp�4E���笍����֟���=l`k3/�x����Y5�_�JT30^�ހ.C+�YAq�|Ł(��g(� �{�5k��e->�܉�~ө�\3{\m¿HL�O��[�BkH&%Ύr�wml�?��ӎ�8[�Ȩ��?�ʔ�>���,�n�Y�����Ŗ.��Ŗ�7�5F����ۭ����R�-��˥�O5:*Б��M�C�� j֘��.T�?'*:�˙[F�6l�������dNL��'��BV���6�����y0��e`�# V_�K��������P/ �	�/a]kG�|��Z��6��+���֔�:>2Ώ�I
jC�\�x�*�cih�J���sٖ$�wh�� љ׸H��m�퀲u�P���ix���}���{��(���ׅO�s�	ƨQ���P��S������n�����1��A��r��T�ћ��U7Ӹ{s�?ZДTG1���;�aꌼZa+D�j�^7��(�$�'�����`w�.�{r����j����ӊ��z{�\U�+�|�_�2���f������H�k��n���D�^@̴��;�}B4���hΜ1�9@a��%�Ȑ��GW�s*m;Kе���q�A�n�	���*�7mW)�ێ��-�HO0�O��������}z\Dds��x�z�D�{8�s�����]�c�Jʙ5���Z���p�ϸ��ґ�da�`��,�ښ����"a[������G�Kσ���_�z���Q�^�����of(e�_�����k�W��,�.�kA �%����R׈��4h�:�]���ğ��~~���(�>���m��?[�x�+�4�+̞|6����++zz�> a��cbۼ΃$$A���d�UO�lB�����{U�a/w������ %o�NUd�1�N�4"�.�'�z�m����ΐ���s)�����!���_��d����L�@L4�u�{�V��~���L"�5��[k��P����mk�RA�LmՄ];��M���#r��:�eCX`�Fr%�Ϯ%3�^~~�8�Х��u�瀦�""��1L�o{0�A"�n��(}m�a.�����m�@�K��^�I�94u5�����,���V>�寘�L�b��u�X���\4N�3��R��>[�]��sh�1��	�x��h�sF�6F.�9ttzz�&R>7��"}���*�[;QG;4�6�G�1�:w�uƙ0�S�V�6���넚�jbe#�o�.�N��߭5V���#:ٛX?�{t�ͬ�1��o�䑕�;.�����] @�f)y��.�3Vn�H���ՓA�����c�O�jk�J_Y�Ƭ��"M�#��5�ʗυ�/� �+W�#`v���ba'����~�>#�-���(�=v9�*.8�I;{tᬈ�7Q�'t�;��#�f�"G+)�h�(1-/�&�NQ�7��~����M��<��E�i�����;	�����2�?�+^2�:P[� BH�-��?�Q��Y9��V��Y��J97N�b�v�}�'w�X!tmu��ۤՒ���¨��K)��F�B���vޟ�.���)t
=WѼ|[u!U��Ɇ�i������J{� 
��s��KR�&a�׻�z��h:�9n���gL*v�����A`XD��6�v�_c�I�rJ�#g�2�I�eƥ��'˾́Ώ*%1�҇lT�v#8���"�X�d<�g.k�ME�:��\E��.=*l��ۙrjI_��0g
(���� ��"�t�����"��Vrmlq��r��Â\��n?r"ȣ�o�g�bH���:S�k�2x����IUNxĔzqWݓ��+� �K�Y�[R��@W��W��[
����9!�?�$6�Zs)M-�t��1
hf��(�$�q]Ϣ�uD��ކٓ7J�\�"���ϒ,� ���-��;�C_���O��-q8:�j*�/l�Fw�~献�Ę��Q d���>�4e�`@�o�4��f�]�&p{ e&�]���L>4���T�3"l99���S�*��^�m�1�9>��:��B}�/"�P��?�͹9�~�T��<ƕ��&p����٭���fԐ��y栞�ҝN��u%����M�Je݅��,�>Mn#[������o�Xw^-�"�ќ����/(qQ�i]\ڡ+����L+�\3C%��^�q�>a����/�R��/�p�%`d�����j}�09&�{��CK��DG}����A޷M[�
�?��6��i�.�1oo�۞�#L���ާ'l[���8p �����;�-j� gvt�g��_�M���
*�%�"�2i�m3�j�M�v���e�wr�f�۸���=r��S3��i!���}btY�g�x+�[7�"N�w�z�+���D(�`r+����lo6�iK	��9c���Ct�w�)i�����vS<�KT�m�p-�t�*a�6���_x�����xQ����'zB�OX\&��"��*��=˒��Sk��X�,�u!�����%��W�z'�V��x�7��&b	A"@ 遽����ÒM�S��Ť)��� M��1�NM8`��;R����Ro��[���R0EX���V��}-���B�T�KlQ���1�Z-��v�zq�"��Qh��|4�4���M%�T�{� �>�@��4v&�v�����4ޖ�=��S�݄�BP��?�d������}���	x>����B��cZX���ߡG�@�7���^K;�cM�)kМį�]ox���ēi� @�|�ࡹe�F6�M���p?��	ش<#�����%����7P����1ܜܱRʿ�vG�I8��x�TM��n�|Oί\����	�����HE�w�zoD�He�]-��+��������߬z����E�ݴ������ȭ0ډ�Z�i����>� .� �8�s?s� �
� �
����<�k@��Iqd0<}(
���~v�P�p��Cri���xl��g���]�l��,�r��Iׇ���}���`�mx��:h��ǎ��)r���K�x��l�]/"}����Vt���u��^����s�
�1�[T��ES�`��LT�\%��	��~/a��q~>�x+8`��{VbQ�4���V��!��.c@�a�#��pa��ra§���+�z)u3�����I�����c>�T9{0w�\R	w�LO������Їy�vvy�,�3�������&�()���cN�!f���j�Q��(1P_t��&�D]�����0�Z�(�c���W���t�1�Kg�o��I�ߚ���;^cq��z��Ϭ����q[c��Z�-�Q�X:�#��Ad�g�>��"'
f�LLn��:�Q�d#��K@'���� ȷM9~���%�vM������>O"��S��� o�H�I��)��s�dY��+E
+P�Y��_�h��\	��%;���샼��X���""��7 ��X���ȀMp�D�$�~)���gWezU�Z�<��R�����٘u�\}�Y�קW;��Y��͘��*[��!�'��&O6|T>]���vU6�.�%g�k�\s�q<G_���ڦ���A�{��Z�A�h99�2Mv��ka\��5*��ЏvnH�u�����4��ҟ�AXo��߃�Ĥz�Ϯ�~oy{D��aχ� Ѓ��}�P	S���^� I�<���Bѐ>��r*��3�u<@l7a_
��G�|a�����J�}��'�NWY�>����|����T���i��t�s�{�?:W����p1���܎��'�F0�����Dƚ�?�[���zeN�.��Ց�p�x�)��FY�6�v=0�`����Y��B��e�Div!�V�I�`ݐ���<��oE��Oo_���E�p�L�����Rc�3���L�M5�������{���@N:o<�8k~Q��>HM'��$\��|����&����%[��L���p{��p��kG���8a)��"���u�m���Ͼ�
���^x�a���5)�^�ɣu��&�S��<R� ���y�@(���Rs�p}R�j�]��wN�S�=�i�H�H5�oDy� �3�Ӹ�Z�`z!(v�4�d�	n��%T�˼"y�d�t�{��9��H%m���w%pC����o٣4.F���r�vE�G�����b���ء?�Npq�ZE��(v��a�AjKO�����`�v	{V����A�`�w5�g�}7��~�C��ײ��va���/�8��ꉘ���}�4�H�C�g��g�,��?[�`]3��<\�,ȟ�Y�O~�@/-�֒�J��t��qf�XW᪙��0-�N�����}:���rk�_i�}K�0��i2گ�%\n�aTA�m/+��C����!Kt)���5��J�,X����tT�����)�Fƈ��`��I��߁����
%��9=F�('�u[�å8��8-L,���q�0�Ѿ{��b;�+���
��?$w.V�Mj�;�w#Q����;L�%5 �)���hI������7x+�ñI|�ۍEU��OIW����!�=Bb	����
�BH���!1��ߗG�e�Ԙy��G��9X���+��@^¡q~�
��Y��J�eV��oo�{�]�zrҴH�o���䂮)��]%�ͧ�X�o���'X�f3�/"ݘ���Rm��0��ɆC����>��x�����N2ayG(u�аOlhX��U}��w��[��`bdH��N8}ҎDqP���a��¢�t��t:���� ���]�,)���ˮQ��߀�U�1?�=cG��'�G��iY�HW�{��L�z"QL�9&9W�W2y(�k��Ƹ|87Ͱ��JǛ���J/j��{�w�ﳳД�1ښ,���^m�d��t/9!5*ߍp����n�Y�о�N�f�<|�HJ�b�~�����4�֐7�.��zZ��;<�(t���ڃ�����G¥>{�CF���rЍ~��&ť'�V9�o�{�ۉ�b�}]V�A��m�E�5Q�8�u���1���,��$����y!�Yj�K�۝Y��}�{K]b��P�_�Ez��~p8��8/�u�~�@TSK>��J}@���]Ί�����䓩�j��M��|�>|e)�C�H���������$įJ��%�����*�E� ���g��f��*҇�&�9�Û:���݄��g�Z0�� �}e1�xo�ڙ�E�S��@�\1��1m��ܚϰ�2����t�=���p0wm�t��s ����)ٴo�#lE�\5����yuN7r��r���>ώa�A�8�;_�^�= �y���q/-��$�m��ʪ����v�� �}�҂VӮ�Cv�?*zł��/L���<�E��ªN�v���o�vj)׏�m�d�e������ʀ�'�T�C�0�<#"�E3�Â�,淍<_ߎܴa��sH��-4̘��"߻g0�\��������K��b~�%�qԵ���
�I�J�WR��̈́⿁z��)ak֣��	W�2�/���Wy=�{}+qC8	6���{�%�A�<K#w>�W6�^�/$�]� ?�|^������w��髨�Fvc��m�l�0R�`��V���V��X����x�C'��r!v�C�ׇ�j��nQʮ�8��gi>���1�0�k%�
�mJ�n�t;�c�0�}K���tf2Xe��I��d4��g�(@K�n)pPe�L@�j��)�LkK/�k�P`�9|�k�`���%+?H+p�r�l�Gw�P��Bb�;��$Q>�[ ��^��|��E�5˰��,�	�aN�b)��VT���=�D2���']�����Xea��%3��㥖�P��?�i<�X^x��<U+��S�6�c���c\Ƀ�}��q��JB�19�btM�YDX�z��_ʽ�p���$�{
.Kp3JAW}}]m�ū���`��@9P-�g������_?��}����1�xN�lJ�/O�O#o�
e`�����\	/��>`=3��c{z�* ,0�2��		�B�P:�M��x/�v���>�[l�d�=d��j�/��5:g�jXZB�5����'��~�8yW�|0<Tr�I�./]B�FJ%�*�/���8<�J�\Y"�['�]�uϕ�EF� d"q�#i=��ۂ��&�N��)#2(��@ �7��9������V9�)"�`�SJv�w9v�Aa����,�Ό�䯘�@�Bpmjhry�B�8q�mӾ$�J��ī��1بY�[F���NB0Zpt$$�d,��|�R��"��U��g�c0#-����9��� �HZŏ�����M�M7ˊ9�e��=�_�Q��J	�>Iz�mIV�q<�Vb��:�俑��!�x�{�1�;6�^&~��Jl��{�g}�F��9���}���X�ݩ�R�+;2ʳ�@<N���xK:N�����P���}� �3EQ��O�*�����P3�������/��C�!�d.K��b����X�Q(q�h���pd�2�2�z�㏕�oX���)�_���Ć��Jϥ��0l�tg�Vuh�͟�ٌQ����y�I��%��
��g9����A�FrgU����ke9C`��ªyL�K�`�e�u�,��鱱k?vÚ�*9��R�_Gd5tI[�0�-��nZ��ut��@co�)x#Qk[]0�ˋ��Cdr���t��	pL5d4h��a1�͸���eշZ�G������S�VoJ�cp&T����a��22mA�Ӵ���"p���y�Z0:L{���<Z�� ���wmzx��/�|�ʳ"�|5��N������2^�b��	l���t<�(;G��q���*XL4l�^L�O����2�c\�g�}����@ ����Æ]��H���1��}ݺ,�j#RX{`�������+4e]k�@�n�V���ٮn8���ۈ�i�f���C������d��[�<+y٦Wc�BuSfC�����NC0|���JE���������m8���2��U��l���9_�N2���\�y��>n�M���5��h���ʮ�n%[��DE����f�&T���J�d,w�%L�Q�/�1�4����2|�2�TKM��&?�F�`�v�})��ZdP?dN/���ڽ�7c��n�5~l�yݐgz�?�u �Bo��D�A��c��(��P5���ג��^1������+��i$k�{��ai���f7n�^H������3J�������9!}G�i�?�RII��^c"G{�g�1�[%	��@��7�zt�`j��ۂeݓ�����dE�đN
�y�@I��x�ZN��e�=����T��?�3���{{*n���i(��w"��Q(����:����������dc�/џ��t�i	�4�t�+�&��t��h��,�3#�����coI��?絍��MQ�`'���D�۲�O�uz&{�|��=hKAmȏ��ܺoBB9۔Rz�Z�����-SҀ��5���
P!�hw�|ͷc'K��}S����U�u\�q�Q���u���hv@�qCO���i-*�h���*�o�Io,������ڌ��̒o�Y�J��u�"�7�
V�[Xbc�A��G���ʟ>^��p���H��O|�x�
����B@�@��Xf7�����Е\���[K?��?�
�sH>�?ē�]�#�`(��"	�u�w�j1E1䡼�
�x���C�7�TV���tm�#�C�
|m��~S>��Z����Q�Y[gRy��kk�i��ĺV���;�h`�¸�	S��<�.?��}��g�T=�C��-b�����fm��2B%�wm霱c��'��{|t��^��4�C��@��y��#���O�G�%�Uޣ��C�t�"��mI�<%��}3�kk�
�d���\,V9���Q��߅��ݐ|OiY��H�{�0_X�M�Z�w�w=!DDBwp�J�"�x�e^$�.�a�([$�B��W�'`0��E��?�?�\4?��E�a�P*��Q^J?�?)(��t��dr=�޻RfƸF�N: �Y��� ��-��xy�iA�f��赨u��l�OiD7{Q ��o�ss��1��+*�V�K^=X������F�5��kcm4�9�[tI�j����m��ۤ"�?���;C�A�?`�j=�mbW�@�š�z未�+J�/���1G�#���W�}{\ 0�r-�� ( "c.-]�ޫ5��`:k���BƗ���uv��Y���&9]V��өQ��rc'�+�������i-��{@O�R���B����Yf���|ƨ��?Q'��(����N� iT,V?�M��.��X���r���Yj����=��,�B�9����hM�h�ڲ�<�j�t1�V���
����t~uM� p�8�Q
��_��J3��?7o�vc�0�7B�`�}�M�we����3�c�*�&��9H��Iw?�rO��Ls��7�%}�O�>����$@ߍ�߱ɜ6XW{p� �<�s�^���|�Ew�[y;3s���r܊4u�T��<�����m��0�Eҝ�j��]h�.�S�)�#�N&a��=��bU#��p4p�\s/���|I	��ܬ���ha*�����Gφ��T'�.'D�L#�(�"N#켗-�,+l���kJ����z&#�Xv#�(s���[ 7��_�Mŭ��0rN���RD�h��A>#,��ۇR(@[b<&C�߀\���RTU��f����vB����4B�nJ��Р���90�Bug���
Ƴw�^̟�k�'����>I.S!�`7�h��vf��t+e|�3����nr����5�W�\h;��D:%�1����Eer�I�~ں��
�p�>��w����IѼ��}�\	~�2�>_� V�.�4��ejA�O@VLv�zIE���q�Wt즡�MHF>�p�8����A\s2a�7Hg,	��1�ˈ[
Ž5T�|��H�
q�(��d��$�#�ۅJ��d��xjy+o��:�s8,͝�E. ����K�g��}��A'݄퉘��oɉ2�k�l�ۅ]��%0ce_����9�@F^2���f�ٛ�U���2ݜ��Ҳ��r���#�"��l��)&x�M}Փn��ۮ"���_��<c�@o�P���"L!���i����0R{�����(MT�1+�H�$��i��^k�	��L.HF��>��v���a6e��~7Ξ=�h�a��i�Ʋ�ĜZ*\��0���%08���8hF��^�a8�q �$�L+c�7}>6w�(O�oM��朆�]���5�� ?��7/�w(e��=��%z��+f y��eyR�	���I�-��ȕT��t������7����(}P����7d��N1IN�%C�k���|�H�ޤ�N�8�Yں�?mΒ�j��E��W�%+Dqx;_���W�4j�J8�o _v��� K�k�c;�tp"Kw"�����B���	_#+
�;b򞧂[(�X���`��h<˞�A�ն֊hGRK����L[�E�p�߱��=^4z��A�e�T��Cn��x w�z�`l��{�g��+-=9����q�%�Z�;���� �V�d�@M�i�ɠ�c�G�%��
��	F�	��M(JPB#�/�q��דT擧��[˗�Z���YzvZ%�6�]5��4�CtYP8��E$,��@93{�sǒb>�o-6%���u����J�Up̒)�0s�1�\�|B����nC���Wy6�ih�	�!a�6�P��]$��y���O�R�΀��YT�Y��6��D?.K����7��K�W�]���|jP���%2h���>�&���:g��"�oM��:�7& �<�߄G��r]�_��(���*ދ��+wA.	|���X
�'G cj���	��v�|��;访�0��M�D3E���\�p��.#)�N%厫&B'$0�?f��}����&./��	��Wp'tk��'0��rzr���gc.�/V�9����螊QS&׵y�s�q��(��pP���(�ne�F.�b�0�G�#�NV�"p�5fL��o��ͦ�`n��;N+�P&f��!�2���E�"���$����%�-��u��T������x(�7���.��<�=E������f���f]\HC�0��_.��vŋE�H�ؗ�̐m�sc'Q���N�|��н2ùh�~Iw(ʫ�8�>\�S0�2�������V#xe6Aft��dp���L�[�o�<��d�u^���0�xO�6�]�+�F���^��'C�d[r���y�L���t'�K3�o�����������k����5���)�c���ޑ[���R�`�>At�؄�
�
��:f�hj�'\4�kZ�0֧p��t�w��D@7��1ÄQ��v%�h+FuPc"�|�3����s(�&;}��x9|ZgCd^�^K6�� �F�wM�4�D�������j)e�%�m��A��
5�}.�,�0�*��e�����e�j�S��|��ܬRz���� �!��L���Lq��Z����ٶ��t���葆ؙS d}d�JޚH�A�)�@�m,�t����j��8��ѭ��[{�EX��e������J�(��B�Iw>v���;M��K�:I�hݲ(L���d.�-��&��JƘ�W		��/#Э�l	�͓h���.��5#:K|�-������R G�"w�="���WG�����t�r%���i3����f�Hۤoy��%P�@3�9 4��4��_8��l^scP<��W�^�>(���B�@�j�O�>p� 	~�	"���9$��^�OX��ϝ'��*�4McG&Fɀ=��$��\�K�.�º����'Ե@�V=�m��G�:�BˡPx�?S����'�M�>-��0≯J��]�������EA���y���u�mB&���5��H_�K��͓���;��>�-�?t������|�S�W@�H4�\���#��n�G� �PR���i��T��Ez��%#3a=�@��6#E�%����x7��VnU�n�4�F���o��|����_�ᲓpH���<�5�� G���*��!p���'fSK���6�	�K�Q�����X�"��ښ���5��#��L�ڒ�k�M+�ٷ_+A� �1-"��d�[�����ߞI�� H��7����d�r��}��)%3�5���t�c89:_�p�Ec����@flL��j��n���h߆F&(��
EfS�t�}x>���P�A�&H*s�^J�/��J�z�jY3���!���٧���3z����糃d�;:����0�ŎxĤA�+�*���蛁ԦX��7��2��p�P��9J�e���!�6�v�j��=�.y��}��k�ڭ��A�P��!G���;n�7KU���s��G��w!Gj�Cb�,��@;y�<x@�{�h?�zq�y�n���c�a��Q��m��F�O_����!��S~7>mBs��a(\��o,'�ھ�����T��5��n�0a�[��z�Ȉ2�ݹ���(G'"ݻ��