��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�? ]r��j�p�V�d�����띜�7���{o|��hg�EbVS����K(�k|@g���)��i���7�b���&nDo�/7���)�&	!%�Kw���qi����N�c����S��g\<�e(͕-�T�d�G�KD��P�j;��|#r����l�|�ݾ�SQ�w�v���|d��2�ښ����g�Ti:f�G�Ǐv��3O�o�d��*J=�#��IX\�T������2)�En���3h,8�Cg�-T���9�αI�4;k���N�� T�"u���P�aT3��4���F��x��r�gav�m� �ᡟϴ�^u)].i[ݤ���*�X{���db�#h�ϟ�j���(&>����,���1=�<�-�����ơ/2A�_ o½���Egi͡8�Ss/�S���5p��A�H��)�U� �aI�Y���C��u�Z��j��-��19���r��WbJV�������1��h
W:��u�a-г���D^p�V���l�U�n~h���ĩX�ӿ�o|�� �J]�d_O��V���G�>�!v�}��b*����?P_먔o��e���a=�d�C�r��&u�'m'�Vi!21��h��|~���Gk{l�?h{ۀ���*`X��E���q\� l���)� ;��c���߷(��q
�cl2"f�t������'�ɒ���+�3��;�����-���2���a��4S^�w�)rm����>�C��(�O�nV����ww���͕��ˀ+�WqT��
P�6FT	��V�����5����	�wK�9/��'��_��?_ra\d�ll<s�5��8�ɳ�4.	�PO[u����z$���F-�����ٝ�eBc�g1�=�E/��i�Q����asO�=w�׻�.F��F�^k�pk� �ք�?'�v��K_\n'b�u 4�G�oגџ��J�����\^\����F֕��iJ��͜6�Ҭ��0��EІ%$m8��3�o�����[/O,S�D���
�z
$��#���sK%�\���7y� �
ڽ�u[�V�<0�؎�Y�W��N�����9�d�̳��t [W�����
�3�K��Ð��� �Iތ0�F�xs�γ��u�?2�{؄���Ě9(�D"��i���3^�y\�H֣˳�'�I��h]��=���S+TBM�al�m��BR��8(t�	uM�4mYڶ%����I�@��hG�ϣ˩qG��邼U3�X�lp)�E��l7}es?��U�%(!Ϋ!������{C�z^�s)9�"P ��:�"��aH�ڶ0�R�e�c�mP�P�� g�'wt�u�6]�
��ԒZNӅ$bĥbe��I�A�Sʆ0�w݅'t�C�L�ِZZ.�l5���]�ؑ;�uB�z߽"@fE�*V%��dc)T� �*��fj����)�I��o�Q�W��+�^4؋%����*��Yo`�ﱀ��t��a�nΑ`�r�@���b	w��Y��j�d��C�D,��EH�| �U�Ѩ��SI_tIe�-�K�.<^}�]�>$�W��oK��(�Ώ��:�Pi煒p4w� ��ey���^��|H�L8a�v=�Б�[�a)���*��<�:J���9_>Z,���f�D�>�]yeuf�΂k����7'���TQl�
�=^�.#�l)H�4�CK��0�� �c� @���hEG2��p{%��E�U����Qw$&Y25�~��CsU0������Ӏ�SɃ&SL��E֔��ff�R ��q��9VEzn�z���B���{i��C`�$�����t�I���`�ȝn�T���+����>K��z߻=zHzޑr�h��q��T��/�wf���Я��}`;�(��#TZT��{���������<��*��fXs�j�����V�ގ�J�"���XK0�s��zB����od�i��U��i����g�H��4П@Ll>@��$����.B�W� ��R��{�dܕ�Z"�`l:�si��j�,L��ߕ��U�"�kF��SI�x�*"}5a��YCfWl�#lc�;��7��o��Θ��|(T�Y�p|���"S�}n���U����
eD����:�N/:��Y�ז
�m+�eN����o��\=�L8�������ƥ&�`��]O�����w��`�vh@ј�4�?N�N� -q����4!ʺ_A�1�`2�
ba�Y�DN�EmxFP$�H{s����S�6���@f�@���#�k��d�~��&�&U���Iz/��hI�W
�S��ܲPv��p~�G(�[��0��xV��'&v�ѣ\1�����a�,���"eSPn���
&6R����u�C=�o�];�H��F�
NM���
��G<�A[� v��ɘ�!�y�}0I��7Ћ�����^qO��]at��.v	��G��|T�YM9��4o�?��ŶB��[u[ˢ�a8�RY��F&d^3����МΣ�qb��r���<h1)�[�Df�ΔeI���%��]V���|6
aR�N\Z�"��5�8��;�N�ߣ`�L�wJ��Jvn��	_oX���B`��au�Q��DNʓt�OO���쐱02����hf6	��]>א1�=�D���_o,���B�Em�8G�Q��KCw��P�-h���7���mDi�rF#F���E m�l��eNZt�O�A���ӭ1ݕ�Y�ژ�<�T�vtŘ00�G�
�y���g�=JDQ̵�����1�p��6������h[�M�F΂����ɴyD�o�v����	��!�jW��]���	�mKxP8�/��L,a���g*�"4�����u�h�O���~��,w�n��1��L��v&��L��������,��T���#z�c��+3S���>�ќ��'��!h"ô��3���r�����[��R��kWr2�C����;"u�op��zY�8m@F�P�QL/6|�2*��̫��+�����`�&#�!S:\FL��DZ�6�sj��Z{�^M��S�T�R���_ uu
h��_N���]���ZI3�BFDD��]HA �2��j�s��U���>ـ҉����K���6�Q�W��C�d"�8T���� �~��LIo�q&u���6D�������W��E^�����!� �`�홓�Qx�pO���qV
«�@r��l?�&�ip���k�8���o	�ܚ�Z�Z��H���Nf�4�q���mM���4��pw�������؀W�c=�ǣs캅��?�:yÒo�'�l�/�	���q��
5�!���g����ci���ȇN�Pm��X�J�G6�B�D84s�!��z��,�S��v+�jK�l@�)~{���+�`�m�S��
5�V��ٟ�gq�����<h
4�}۠W�S
+����hy0��<~��aMZ!c$N`c� ]PU�x �A��
n��-�Uy�fzX���bھfn��i��m9����H��3#M��/�����-I���|�$���!��@��S ��h�AZh'�z���!V_����}7�����xx����o��g�]���U�Ȏ)�6g����<���%�K�<���]Wwd�N}���%��u\����6x�vgz���n�DŲi�K���?W|��a����F����o�GO�w)6$��*c5���ʌ����2�/��̔�b4.,���=;f� ����|^<�o��'{�b�%W���&`���� �g�Y��8�Y���H5D��e|�
wZ�J�1sg��~f�FB�����r?S�vW$��H-�Q��Ge'� ���d�����ܟ���]�kE<ƻ�@��U8T��R��,)E.��qkJ����7p
|U��2L���e��rG��h�m�٭�	�q1wT���6��*@�hdN(Hǯ2NSΔR�n����
Y��1��!�p�Ss����(�.���m��d~[�� �D��^���v�r+Hc���1j��
+����+p��,�U��h����T�*r��槖7����H5^[q+o��st����z?��|��E6d+:�!�$�u\YQ��2�=O3���K)��]��v��S_$���S�� ;��NE�[/1�|�J�>����t3�N���r�jԠV��#�ǆ`�x�G�]����
̍��l�n��68پ_�����i*�m�Uʽ|fzbJ(�q}�Ї������k�ͣ,E�c��>�.��"��E���l�a	R���U6(Q�ņu�w��)Z�|_.���j��֜(��tX�hQr����31����)�'`�}L�1LĆ���#� �ԯ�/�W	�G�d&���s ��8dV/x~�)�#̃�Ղ}����f��CaeNC]![X��mx�:O���G�����Oc�KN2u�=�y���?\3���ԕ۵����n]��y� Q��$��wH����ք,:d�Q��"�������j.ڤK��I����J�t�ѱJv� ��}�ϙ�'����2��Nԓ�	O��?�n_���w��@T�CQ}�����3��U�	����j5f�8���w��7F����7��)�'i�*A��k���dZ5��59��-��'8f�V��u���\	8ܴƄ��ټ�	�B���s����]��r�?���e�T��ء�6ӻN
E���$����3��m�HB3^������5FJ������g��CAg�1��_�Q�ہ�{b<��,:���tQ��������n@Fa ����Q�a�ȷ���%9݌��5����P[��S��=��lr���}�_�Gm��S; Z��B��
"%!��y�~'����P;[�q���wW� 9FR��������ߵA��^X�M��g��@���N���A�~.��Ѥ��~���lm�#I;\�~��p�,K&F{�������J�L�6ٹ.��9Dmyb����a@ي����$�cy1$i>Sarb!�+D2X
�R�3zzbph;a@G~GG�@+�	����Z4Uv^N���ub�Np����)�>c= �EwFR�_�2��-\�7}Ap�y��S��n[r<�4����P�t�;�O��U�����R虄$�#�|�MS�T+�O�Z�e�A����x�`�m���1��gƺ_M��|�X��U����j���J�O���N�@v�]��9���Sm*�T�ͬIJ�3@��T�:�#g҃�@�Z�<��{ؑ���²���`�Љ:��\ �������2��eoKl��/Y1�vҩ���ke}n�8ܘ4?}*$#����Ctz���t����8U�
g��V�#Řb��K�iG�I�r,l��!-���M
��zZ|�vy�^����:S���wWڪ�T�#Ix66R�<��3��g�оHe��F[@1�� p]���t��n:�AZ��ɪ9T���0B>O��t�p�孄"����?t�Y\?�ˤX�~��/� �27-N�����4�Α��������t�Y+��<��\A�L�����"[���䫌bd) �k�3�v����nGOy; ���x	w�[�Hv���;o�mB���׌���Y��FT5<��WP@�@��-��/i���	�~)�s$�X���V�x�P���kb����)!JC��J~�P| ��q.�Q�*�:%�|zP����Uv��y�d􉫸XdP�ٺT,3�����y=H8��UF?7��!��u���ZA?�X�H5T�
'���/�K%��Q�!tJ�}K�O:�#�	b��in����7�p�3o_��#���B!T#��������Q>�̽C�)
+,C�6��Z�"���e�vT�;A�Uk�Y�����$�(8��}늷���U��/�V�T�����&[4q/���^�-�.
�@��I���e������̭���zb�Z���pl�-~5�P���&�8�'�6����A�|���eͬ�*XƦ�Gnq�������� �O�u���e���옪�>ݢ�scZK"�Hx�~K���A��Ρ�}~�x�>1�L|[!��~� wCK��Bv��A_-`�[����F����q�¹�Q�1���n�Y�>��w� �9�@ub�����7bm?G?��\����� I�6��fРг3j�[��h�`$N�Z��D���ܸ�F�*���x�h뎠�ļd��Mר�YD�������H�pm�W����Q�D��A�6�E.��mM��a:ۢ�4�I~e���Y�)����5S9�ؔG���s��kv�N<+R�p+w�iѕ��X���6���Rlx��(70�ۻ���+�V+t���G�����P��!L{w�O�z�\�&�蟖�?����5Sϯ�ucx�@�
��%�P��Ouv���'�؛mi{L͡���ZA����$��s�g�[ f;�'���.za�L7�HC������3:  @�������~����uh�)�イ�����'�gq T�8�1	��(��F�z��Q���T�`cʉ��V���T���E�N�R��r����꯭�skj�P�%U�8 �	n������!`��<N�-�$C4�
�]8�9�q��~s�z���Z����.i"s��b��#s��Z�4��Ȳ5�M.0����ОB���J{a���Y���+�c�8Ji&K1�Us˪��ra�1V�h���^�*�2trk@����Ǔ�F��JGH	=��\:���4$�q�X�U��8ԯq/�Ng���b�ªr4�]K��8/-��g^@�$qZJ�rT/��[V
�F���_D����&�N��R�~���=$�Q/�Gюj��|`4Ҳ�pIT�0�6&&X{�X����#h8�(^��T�
���!
cL�%�F�2Ɖ~LfT/YN��v�>���4��lRޙ�&����l���	R$sf��8
���dN�ǺӜ��w�X��RՄ�֗���!YeӋ?E��f�WF����>´+�3�왶���|�4�X��&���(��oRû>�b�� ?:�@p<µ!��0ik�|0<~�K�e�g��2��,��K�$z ��.�2D%�n���:��!OϘ����Ʊ9!�@1�E_�\
'���}3'����g�
5w�~RڮOm:ۄ�0�ж��,�;�X�=P~�t��N-�+ɺ�.rĮ��78�ŕ�ک����I�s�;���Ӑ=h!,���:{}��4՝�� Ԉ�C�*ir�
8���?�曶l��Ox|dm�lb�����I@X��4��n�L���af��Mk��0y��k���Z��̗�Lp&�z�ͤ0�;��;�/V��롐������z���^:�D��;%�k����4�ɭ���oS���}�?���-��5bJڸ!v��\XʄbK�#��hݜ������b�}IMT�3&'x��"켈�υ�
��dͽ$Y�����a�{�Ɖp_�;���Ń�����S�[L�"�hK�<AK�ͩ���kJ��s�a:�ϗ'Td�k�[6h��}��޵���1����a˺����D�/Q_w(T��A�� J>pO=��M����$���>���p铝�QFw�g]�q�ݸ��`-1*���R1M[�7��2�_�F�H�œ[�k��:v|�R %O��B҆�.�	�dńIX/��?�NvJ_05��<zg��vo��dk�Q$#�����N%��0�W�Ў� 2�f����n���fWү
O����Z��ȱ3�1q.�޾����o�h.��K�')↥�;d�i�g�x,�Es`�-/K�:\?�f�{��@���gs������6A�p��B��|������)�Y=��ˋ����=a�K�}\�$'&W�Ő�t1w]>a��Iy+�����e|H�o�izƍԼ��sZ���YQF\ҤG>���������M�Ypv�F�O��\n��ICF��ʤx���N���p���7�<�@M�T�u��f-Z�����Q���m��q���sI`�yp(
�;ͧ{��Q��z���T�:���IWn$WJ���T �u�$�6��4T�"p5������_�o���='�-4($�e$Ʈ ��L�3��$뚅���tuG��mG����B�y�p�G�ocz��7��ށP<x;*m�e^����8q�(�s�[�ߊi&7��=�@�ЙM2[!�OQ@���S�eJT�W��e}�up@()�`v��Ѥy%��������G/��B*�o�0�1t�X�/��WZ71�g��V�7=�X�.�E��i��63v�I@Ɍgf66���&쫙�J��m�0+h��˧�wLI�|�F|���%����՝m�C�+��H��>j�,-s�!�z��,$uF��%�с���a��`��u����n�B���i?�XqO
�;��F<d'�!fQ�;c_`��~�i@W�#�4�M���t�x�h΍��e�qZ����Yw��l�.��_e߬8t�51hn'�E.��e��fj�[�a٭k\y�<���8Er7��X�i����ճ�;OamG�;�>iL8�(\gh����;C;�N7�E۫��;����/C���iT�NqҞO�'�m��ef������֌W�La,����u�h�
.-oHލ;3aI�=��ZPE�?ἱ(�#ʦ@�fB�-a�o���m��1ky�/����.r�1���JoLVB���QH���e�N��,���wnBfX~sh�,G������;�#^��-`wd���/�B�D�8�u��or>r�G���Ɋ��bL`�h�����suˣ�D�~��WO�
���dz+�x�2{��ȏun��X�rlNO��NX��;j�W�[<�m狑h�.���}t�����I���i)z[�(~���d��F�n}�̀��������\�{�1���_�h�+�v�˭��p�� �Ġ�r�2�Dӎ�f��x�J��*�4�g��b������*�z#n�Y�@v���'��WRt�X_�q���EPC��FF�(�
��<F�Ρ�׆�7���t2GH"K��x�G�={�����_���|�����P�y|ej��{I�)z�7�Uu�N�ظ��zp��iSfR_������D?k�2Ż-xKh�X���Ii�Ǿ������A��NQw�,Eg�����_�LI�A�tI�S�����#�e5���@4�����f83����1jK# ����"�0s7u��� 2���>�BX��~h���mfm|6�Zb�#:趔����g	�w��vu�m�ǕY�T
��izGRι��t���Ru$�N�&�V���K�v����l�0p���M���;�yG�M��u��(u�����Y��N���c)BE_�ZyH$5��e0�c���,8���g�/�S������ ��\�"����q�#޹%Ɗ`�Td�(\�2�b��$-0ʅp	��#�_��r�5�ܚ��U/:�Ce���L��{�;=��v��'���K�(�>����6L�U��aF�-I/�u�_��!��m�,_��(�*ŭ�`E6�TB�Vi��v�z<[2w��=��$;I��.�;�YC�i~q�����a���f G��5�/��l�9��.�3#��B0��������h&+�[0^k�;�ِ_$D��]*�ܸ�l���q�{41�4�f9"f��b��b"�����s��H�J'oK�d�$�)��L����d�����C����fd��&�`��L�q�9Y}c���x�Ȼ��`]Hk�,؋!2�D��JB8K0|�j~/���9io|QlBGݎ���}?� &s�RW���1ތ������ ��*Vx	؉i ���E�,���[I`����f���gHS��.x�s�l}�[���ҏ��E0���Y��(Z��kw'�$�c�p��fB�E�T���u�_������m��V.�ں�]�����7+Ͳ)�J'@�����m6r�!fn�����m����$�˒��>:�U�ۭL�w:j�.��o�f�7���s��Q��seڵ�y�K�b�,� I-���ؑ�������a��[D"}��v���?N��m�3����{f�Z��d�}~T�Ǒ�I�?ZIJK�C۵�R�� �t�{���?��Rv:��$1�T9�$�"yB�W���i�E/�}�^șE���L��b� �T^��0ܧ��}D� c^h1��@{7o���7-�(�yel6��dǤ����0��6��:����(Q��0��8;|Q�h���^��W�	���毦��޼�=G����M��>Q�g�o��]&�����x2h˻��Br;����1�{����_b�Hb�����-���懟0J�g�]�kbp��V��p�KL��lwp��Q#�0��ۅ ���D���z�B��XST+\!{� ��b�}	��H�ph�cنGá�� %)�
ݙJIG`�oc�䰻��I��!�G�d�PB�Fyk���;?X,��MI�PuY�"n��FB�M�))[�Bo����|!�Bj�;�L���'\1)Q����!��-+Q����Ҷ�B	�m>�V�#wY���E��#D��ZB�x��'
L˜��i'"�����""@�D�:_ͥ�wq�&(�������.������ܪo��+��ϣ�p�s���<��m&�`��L�M|��qik#���]��eD�Yyҫ�l�}�2A��h����:�U�W�et�}y�����a���J��X�I◀o�9�U�}0I� jb�^�PQLQIW��[%dS��s�&xd��M��H�>a�����]FЮ������X���h��Z�M<s���r����8ϣ=�Ȝ�]g�جi�~��eه&`���Jh�&k��c��i�8�|���hQ���t�.J<�.%���JK�ע�<����Wh�T�H��=��d�஑���dI���� tm��axJ{J��:5'��~\�Lt>.0G�@	�5��1���c��i.���"�V^˧�H*���Eb�qʔ
;(�ɠM�Ol�m?���O:A'�N�S������j�5��w\��hʽd%��hI>B��u�̀�B�H��;F�'S�j�|���nף5�,�� X��XZ���b�����8cG��N>�8�&\�q}P,�4�R���T������Aˠ7-K>%Օg�y�2
b�U�<o_��yzYx��Z2�wf	AY�@�M/�f�:0+��n�����m`Q��W;k@�]DՀ0=�v���\���@}����o"�.������_3��p2�v��j�خ�?s���h1��������Ƙ�K�
h[8��l�Ü;U��?B��mwH�D���©�7���zD�||�K䆎<��@���w�S�s��&��h�}��&Yu��'�9T7����#�B�O�XcZkd��e?�is���LPH1/���P��P���n�E�6ׯ�pUu��xb�[����V�X����q��K;r����]��by`�f2Ct��W�+ q��,���P��a��h�&s��r�/:(�O�8��A4�M����(P���3~�Frq�V���#�����}��Q�E��B{�g��ƣ�3�wP[!%T��.ޜzWi=4���j^���h\#Z(�j"�3!牄-y�{��|X�6I�n;[R2�!#���Bf��P�=ҩ��K��C����9Rk�W�(��a�b�I��g������Õ�>^/l���y�O�N�^@/g��W�-)1�����X1��,��o��FΪ& �	���Eo�����xL����n]�L�o�nT?1�z�c��Mٟ�ov�Z�˰��,>�Ə��i��l�|�t��)�*�fp}�Y����	oA�x�A(+���X�K��"�!G���y6�ξ��d�xػ-�o�7F���ͷu�w�7��·xH[FLNJW��}������m���|u��3�$u�aa@�B}���9U\����ϩqM�Dy���)q��D"����ݡ!�}�3������
��lf�pM���C�*�P���x(�Q�Sn���]�k�ĕO^#�A��&)��@����˃|���
7g�b\J&nB�.Ԣ�ǖ���������s���r�?/(��%�(B�Mk���lCh��x�J�ͪw��T��UH;8�j�Z�(��[�\z�I�>F�+�!z�n�?�/R�h ��kY�}]]���t!�~ED�g!�*���디)�G�S��4��-��_��'__�� \;�L/�#�2��~|��l�\�S#������Gog�����G��`قB�m��!Â��W�9-j�jɟ J��E��x�`2�,�_�*�`���f]thQh`$��[�����&�[��!f��C��	�6�aQQ�����f����s�W�p�x�"��DO�.�x7"�$�ցƩ�$��NT!1��}��ck��xk�4��=���5ԍ���l�8
�'ns�_-{��c�'i�I6ӎ�λ��#*�`l7��һ-DuMѦ��kfr;L؄�'�j��k^�w�{g*�i]�m��f�R���'��[�c4~|X�A�}&K���/�󒞅���<4�I��Ks�%�1�~a��{�y�a}Y�̃X�-��2| ~;�t��?�g�C�%-h[�t����K9�i�Bfr��L�%� ��P^nkz
��횳����z7�����(\���x �`T[��bׇ-I���%(^3�u��x�����	XBe�I�a~���s�$��sN�H�.��?h[מ��gV��A���E7r��4[��"x�Jd"�)O�Y#N��L��y�L��[�R�����=1�O�	j$$
�Z���-�.3n��c��ֳ��͜�&�)����G��� R.kt����q��ud�2�К��F6���J���}q���i���l2s�*���&S>Ss����*��x��F��_3��B��{ K[�k)�v��*7�*���I�<k!v�)ݽ¥���.���F�Uu��"���h;k��D0Cj!;w����`/y$YP2����Y6=��)-2yR�d�S�-?�MѲ_���u�P�����ZW�T�0�՛Cq�1��C�b��4�����-ٓ_����;������y��4��=Z4mc<�kVXy�?I�P^T�4r�jU�]!O�~-��h�?�9C@�fP�Ht�O1��8!R���p��g�]���=�DU?��^��Z2��&�іG|GX�{"��e���U��L**�^T�%|v��5�J֩�6�G.��x�7l��Z��y�$��sTYb;��+�3�hw�B�<��4��碉��#��.VPs��S	�R� �l��D->5��:���
f8"�Xi~-D:���F���\@s{Yr�ڐ㇌�����F3{�P�^�@e)ĹqI�'�Ϣ�kX���@wx��j��2�}�Y�A�T"��
��	q�,��T����2z�(��A!�=�i%��&���t>Oj��O�(խ�/��R'�X���K�K�,�bSl�f�;�������I<�Hw(��~�G�Ĝ���Z�e�Wt�(�&bbi�"���Ga��(_�@T;E9�D3�XĔok���m�ąMku:\���(�L,�(b��k���c��n���x��t�bA�wN~�!/�H��-)!*�#+8gi��C�c�H[����E�{�$�h���q5��=:�:N��!���N�w�ߥG�m/�v�� 9����af1ն��hV�S4�V �fƋ�piQ�<Q¥��T
J�e�%����g�G���*�c ���/�
IǑ�����K��lV�+�ZLHP�  �
7��q������
�>>�(����)%�S������x��������9�ޞ���s��9�cX�e�<��Tɢ��u�ѪI���,�c���D�.�7���gf��M�*���;��h��ļ9� ��0H��D����Oz�=VSv3#���'��B6g�9��L56S�Y�N���U�-�\+�dvmrϞ<��l�k�ِ�}����󢟶j�ya^B���:K��X�v��
�2h" 
�ovN��y�NY�%�*�I:��E�?�.Jh��6��zm�`�)�_��Y�g/7O��C������+�_}�W��^)��V6������E!Ԋ�飑������(�������b�}�3Z:�_�hP��4U�,EC���&]�l���'��[sL'�]D��N���[~o]3�e/� tJ]�':��T���ٹ`��s?����JԦ/��[<��zJN�gC�L|�y����f��K��i�9�CB��2ia�5�$?�ۀ�FkO�ud��@�n�K��뛒*�nNb�˩)�����%hxO>잀����vN;�
;�Nͺ�?� �Z)�� /�E�3���ٝ��+�ͧ��v��r�ű�;��F7x�j��ÁU7Ԏ��7�I�F��Y		9�v�Qo��4�_A"�7������}�hZ�Y�a�: K�Ũ�M����ɇ�;N�Xmܱ��*J�κ^�e��EhR@�p'�S� n��������Dn{�|���,��Ʉ���"�f;̳{����5�F��B5�	���9dk38��Q� ����77���b�������VQp�ik,-�L�ZU�}�(21m���o��|U�0g�/��+P��cR)�,�ኀ����(4��75vk/���L!�ʶ������3��1~�`�py;b$�n�tBy��&����ź5	�0�Sco�8���L�"^���O,� �S���Z���AjP�Z8h���G+�������g ��~��Oc�"P����� ����֗L����#�����o_^�֒1�V���_Rll�Sl�%N���n�`݃���j`k�1�������۵��e�I�C����b��j��e{e����	�����ɊT-Z���Az����w��xJ��u�نAp��t1c�q�$yM��ߘ�H��&/Hi������Vfz�{�u�+�T�]mL��u�\�u6aU�Z�[]G�F!!���V1�Pݨ����h�X��4�0��F쯋y���@>��wL�'�C� ��ݴ>꓊�w@�:�A#-�����o%V��/��&%�5�a��,D��hF�|5,	)�����-�թb�Ϋf%kN�3�/�z�?#�� �ѧ�<:�M�,;*��c�X8e�����6K�I��,�V���������/3�(��x�D�m͔y��蛽l|"�iA2��O��<N^�WJh�O_h�N�M)�_�X�1���!���\�eQ
M�d���^��uC
Y܊E����0���zq��(�f�o,"O�@|�@�$�I�(+� �}<)D�#+���иG��=���.b�ٴ?KŕJv��X5p/̉č�����u�m.|*�0h��ĩrH�6K� �~v�+��-����f��!�y����u3x�0�	`z5�ommOU'd!�@�k绸;�AQ+����W�-L�ԯԴ��{�3��V$	�(�q���+���嬰�@����a��OÆ"B�2�Ṕ�S�6iL�vP��y�	|�_���H�sR��CK_߸3
� ��{��v�>f�vV���_��'G4̃ͯ�Q�J<Nj�6`���{�Lю���d5����v��^�:W��@�jZ�O; c�2�;Ō~�v�	�1==�Kup���t��l쒧ٟ�uқ�Ȯi�TP��us DV	u�-f��9|�\		U� )�	�+ '��k�T�V�(M��;�ռ�B�� ��uq��/��(v�]��K�2+�'ri�=|��a][��c�W��fӲI�9���b�qT�r�9�!�X�"L���}���,/����pS���Y�b$А!�
��
�q��JV`�9�phS����9�eW������*�P3����Z^J�G�F?�Jxd|�r/b�;uMW��wd����nQL?5V~�ʼhSU�}�I�*���J��K���U�I��t����&�������k�#�G{ƭ� ,+�:����;��ɯ�5"��F)g��p\fICX��y�^��.���G���i�aLsIIe=dk>A�,R��NR��j@怍+_T����z�K��TG����*�� ݝ$D�4�y;Qр�y�R�	��	���z.d�C���,�3��=^��;s-;;�#���	Щ��xJ��!$zN�F���T��t&��f#!{y��j��Gĝh+��컪f�HîR�����=���'��1��p����cV�+�	��n[�&�fA:�	��q���1np~��{0=��h�t�����=��݄�5#��!��W�<T�C�If�b�ӘI����7 ��2��b�J<� }p
g�Jj)u6B�B�G��GM�A�m�:$�<v�i����e|�}�
l��	�%��x<�&�Ѣ�,h<�T����ũ��]��`�U�L���n��=�f6�([���T�s��w��
����=���s&���^��z3���i���/,Ug��蘋���\���!�{l���`�e�H}h"��Y1��]S�2�|JNG��H��^ԥ�ǳ/�����i�zV�YlKx+��#zњ�����bfD�ikn���*>���N�9�ʀٕZ3��C��'�����<�T���5���"�	���V>S6qx̇Y!=���R��s���kr �!>�������>��(K������邟"ZD�<ٛM���8kd��6L~�s��Dn��$u��T+C�휢��<�����A�:�s�f,'rw�@Tdx���a?[�-���)'�x��Y+Q�#��dі��"�w�Α)���$�õ��<�4ۺ�$W'NW����xN֒�Z�v\�F�euy��5���?&��