��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S������0u�ҽ�s�!���ةt�)�o�Tk�i��m\���W��
Z��>�� 8���9�|
Ce>�22衣��\���"w�Q��=>jUj���-���]N�\��ԏ[��8Ap-�x|�0�5sH�ƾe��3��Y���;���������E�Ȇ�+ʮ˜�!��-A��>�8��X�Z.�c
�|��G�ػ��1����$	�-C}��Y�1��X�hX���E���6�R)_!��)/����Ġ�O���z�¿
<����Z5�^9&�s��|WQ�������N���M��4M�sиl�8��k�k�j�:��-태r�/OR�^��[�ا�o_ �@��µ
լ�>��/��R��u��p%'n�q^���㚄 �Í�*: ���~�w�?A���II���7�q �ϯ1�"i/����"f�r�nY�S�b���P�	��a(�L���V7��^p6W1��y�#�b�!��[�� P�ӂ����Oky�_��`۳�c������L`?���nzJz�9/����195U�GIC�=QHDo����u�ʪԦ��О�&j�	�&u!�t�3�Hvlȭ�Ւ�%�xGpoIB$텝J��[���D��(�>'JQӂj�����]���&F��*D����"Yw^���c�{�r��"�>�A��6w�^��vf(1b��)	��.�҂ds�0�t��V$`�����(l�SǄ�'�!%���w��������8ތN�����,(:p�����^�J��l{��D�� �D�L��������|��i�-j�Г�r�W�R11��Vlbq�B�0<�Z���e���<�\�ڜ)��Ŗ\� "�{�h@Ǜ�R%�_����)K(��:M�Dގh����76��=��І�i��I��~׊��7�n:�R�n��%^2��HV"����U�%�ݒ=x����$��C�B�焩���b�sWӰs3�q5la�,�@�h<0;\�[��r)Y�BgB��S� @��@�V��jE�D���tu9�Pm,-g�s��G+�����u1wlq��I��u���ą����jvOU�9���kʟEߡ�W���2z����;�c�)��u Tl1֜9A�h���yA-̱��Cyu{?
D��rC@�{�#���	�YY�P�_��,�-'�}�a�A`m9=�%A�BCF���t�P`qPq�70�EY���`po��A%����~�um��b���o���K4��܄��%��pw����yMX���)/^9�UI�!�#�9A�	,¿���͹����W��+!j6)ki��si��UՓ���4g���Ll��U*-Jx2 �f�<�����(hk�F� f����oY橆���ԘcBm]���~FbB�X
����
=1�8�vݮM��{!��/f��m��PV6�a�b<E�*X�B�0"����V�E�B��C�3��p����4t6L�H�B`��?x3J 7f��T=���Q������pZ�6of'��j�US!n**����~Yr�P�hb��f�m�3`X
�ۆ����h"#�V�YwKbه�ư��%N<o�Ւ�+�W�WxN�{�4�.2�X��5Ʌ�R�3��G�#^+g���װ�{7Ou?�:�{w��%@��=���J>�E0"�6?�K�� ��X0�̨���և�:�cޡ������(�?N�=�T��0�@��QE��X�X������(�ap��e[-mb�Z�չ��>Z�A�dB����Ƨ��_���|�4��B����׾�߉��@Tdo޴����4|��h���Q�SO�� ����E����v�v�H�l�*�*)�ɱP���پn�����uowƉs~�iKh��J7��5_=�<C����[�>t>ycNh�w��JMZ�g�c+�],ۗ9Wp*Y<���� ��%��."oD�^�q	%B{@�s�tr|��nF�����׺��iD-̦nf�e@N�	����c�������M�WVA�؜���Ɂ6�ѱsI�境���'~�8�d�����*̀������A[	�7�"%Ԩh̾3l��Q�}'N����y'u�4&G.�s�\�9`��7s�&�D�<6N�U�,��{�w������߬��e�U;J,2%�V'�=�ò�{���A-/����ą��P�|}�Z`�Ь�On��]�69�h�p} ;N@�m�Z����
���a��=h7��
}m��[��)�
g*Y�Q��(��z�	uW����&A<�:B��RCo�؍�PUa���kq	�;��8#�]�Rc�F�����۬,1��,t��$�{�g��}��,�v�sU`��<2C�Iʖ��}�kU��0�3�
R4Um���\��{��u�(����E?���UJ߳w+y��^"�Y6�&�j{Ĥ�'g��'ˁϥy�o�-����ԐDW~����*���D�J!9a?�8���Mֺ�<ɀ�w����\D����o�q��#O�0f��sw�����B��6~�a��տ��P��^^_���������8�Uk���l������.��i?�����!q���a"̀�xM2���>`k���D�����n�0�K[Um��+ș_����)���Zw��a�Xj��[7��Q�3���b�u03�RB��Wؓ9p��r�xf�����	e�_�-��#/����6#d�o��C`	]L����s�W�(�;��Xt���t�_9��+��;�Lb�h��QJ�Xh���H'���!��\S��B؛#4*#�Ͼm^����a�Z��H��=�8�wt1�
8����Oˤ�Ʃ�^��a�fO��Ӯ\?�PW���w�̔xm���@ݛ����C,�Ζǫ���K@���[3D�Z��"��P���*e]��_��N�U�`��r�9�L�^������!���X,�bX������{7͚��tw�uCR��*��.*�ZS>>k;Odp�k;�a��L�c��� �Kpic��	��<�����F@|jVLO�������l�
� ��k��Y���\֛�?i��l +�	^O=�	n9b��Sū�?\�d��qmZn�J���Uc�%ՠ�D��<�B����^��%�)t�7VuՂ��W�ϛ��
C���8��±w�.dCFЦPʱ�d7������@/@���W�������6�"�,0�����M��~�
۬9W��L�A)����ur�Lxg��t�J���b��߀�����ш'��{�8�H�vO�Q�"����	߰e�E����q�[4n�p7X��Y��>26Z.��N�#y�~�9NM�s֘4��2�#NT�����֎C�����ъ2ufb�N>қ��P]�f@9�8�9��ԒKV�/�_M��l�6i'B�A�i��D^?��>-�&�c�6���t���Id�]2Y���,��]M�3y�N�h}�@{,�91��Z���Z�r^���ky0�'&W�o��|J�X(��_�Yo�u^hB�
�rû��ㄖ�7�R_��&��R�蔩�wm$>����zkf&0�6闩@D�v�C�P���w�o1}���K"o�@�v�ن\��%3��a-���t8dЗ4�~ﮫHJf�Ѩ@CH��QP$Q�]8R]f:�'\E?��<��Yi�zPH�_����=���Z ����w8��=�3z��w���Q���O��
gKdw/H?�_�2��ёD�#�JE���5$�'���@�{4(�|��Yq�{v�#����Y�kF�f���*}EHim���D6c�zP{	 �&G=txWZ�߄�g]�,��}]���~�.�l�9��x�2�P�oz*�����y�v�}_6��"H�of 0�或-*WEQA�ad�i�H)[v�����r�8�s�%���p�������Ԣ7�u�q�g��s`H*(f�OZ��GM��p�Q+�Ċ��3�^ؐ�i�v�5�)-)ה׳W���[����gB��|h8�\<(����?Z��Ǔ?Q3��\U�i.���b����CڒMՎu�ؘ��5�������G�a���>�~L�4r��m�!���{�b_ �fk+J> ��L4	Ӄ�,1z{Ľ��˙!a��N�J���)��dG]n�@we�6�/�&]8�r��N/>��t#��jMY?-��DZ�Rǝ���O��yi�	ٹ{�H�Ħ�ȹ���~�$��A�$R��Ф�(ٙ����'c@H���'л�殍m�Kx\�#�b�C�C�Ґ�мZ�;�ˆ���]+�IA13�%�,X�$3��I���,̢������!W�^z>��Am��@���u1��!��UѲK�q�	�+� r�䇈�o��ˍ����q�P��Z��/��4�>�%\A��3��x3*��qؽ�V�P9^~>��on��o�8�=,��2l)�.���E]�+'�e�����sqb�D�2���V|��Ɵ� [��Y�̶qA9� h��!�gs��
`e�qj���C}�����' K��B��ēh1���>��(m��]�l�m�O'{�J$��3v�'�}�#w�����������sohlLm�+O�A�n���/��b��ϵӂ��ƒ�[��O�璑L��v����05�ٯZ/��Z�B<�k���cy3�E=s1P����(�Zu1���%�W�\Ys�1<[�!)[�~�/v�{4/��/���������3����|�����S�=��ˑYu �UGr�.C�p�F8�cR���̂�]��;�,������:}��xu��^5��G?�c0�g��MV?�"�HOK�*��4V�j8px�]���?���NV�i���v�`�N�F\�_�{��'���������0��/0��n�V
��|��S�(�G"��KcS~J� jSy;2��_'��\�e�n�1KAVz؋7�����}O����gϰ�J�ʷ�Nx��6\� ��O����P���_>M� �{4�f��]%O����������j�ۢXz�V|���սt�[��u�P��lm�|_��dp�Bl���<"�R�= gf���j
�ߛy���P���ɖ��8ׅq��������o���s�s2�����:Ո������4���Id��Ԏ�İ'�<�q!E���[4��&_޲�|���'z��X��c�bP~�����@��>;���e�[�N��S��ԝ����\]O���رt�;��W���,#��U6�˒�a��:�{�1ڪ�f�ڧ�T�P�H���>��h�H�T�ހz�-$��U7�tNy;ϥ��E�"�tw��9��û��-KCt���6����Z��0=Z��B�:�6���q��L�E��Ym�G�E4yIpHG��/��h�1NQbCv�I�|hKϒ�,�*�{�:���֖1�/�
t��'���hZGp4��c�W���-�m?��ԙC�PŲa��w�M�٩Q��gU8��V#�̞����]+�D��Vk &y�*t�L<V�rσ�v�H�?\�W�F�ch�Wc�Q���|C�G�D�1��~D7/ɀX���G�~�����������7�y-X�����y9�m���{�1Z��!�	�[��U����;�hi�l.za.����g��+R8�	\�C�l�1��88Y�c2L�8ڞɿ0�A��1���"&�w��&(�I�G��E��|c'��0���A��A!�|-�z�jp�]ہ(XzE�e�:򹟽�ɮ��jh��]���ˀN4��Amu[[\1O��g
�kof��CS���~WY ��uy�wgZ6���vg�!ŀn���=�G���[��TW7UT�#���yY�k�@Ka�`AgY-/�IM���B�-��q��� 
\�����j�=��W�����/�9��'�T��q���t�M)��Z$��]t���)ݺ��Qby�p��05x�[,�D�j2�n�El�{L-7���5��C=T-g��R����7�W�2B��˼���ɣX�C<J�d��l�!��ۂ��s�e��X�t:�ш�J,�dX���ζʑQ����#9�+>!^ܜ�:� ͱ�T�MH���h�
x'�byĺdc5��Ux�����+��J�B潃���7�\-�/��r?��7@;;%�x���'���ju|���
���!ǌ�9R��6�aL���9s�h@ݛc,�2� �y'�y]��C����(|ڠd�q��f�_ּ�)�ʗ����}r���Ei�V1
���Ay:�И_�u]�P&e9��W�ģׂuB��{9����cu�p��_�ѥfIGn�n��-9T��̸�d =_���W�wjF�HS��ޟ�XC�ÄWl/��I�ǙQ9���ܳ�S�%_T�䍀&0��i��Mm�8qk��.$�9�?��R�l��j��ݯ���xC@}[�RA�d$��՝�DfE	o��HL]�p�m+�Ɔ�/\��Tny�!Gf�`k�Ʋ6Jy�xI�B�Ug7v|Q�0汸�:t�҆E��:o�uA�� ��j}s�֤�Z>eY�T�F�+)��#��My #bg�5m$v��_y���.o��6�b�[��5{N��Gh�x7tc`�ڝQ�`t�b�sY�j��o:�A��co���bG���E�dC����$��ՠ̷Ja��ӊ�ڥ	�g5B
��:�@�O3����HA�)M�|��I�z�EdP6}%����\ϸ��d�d�N��M�u���;~Bl6p샾�O�[�"�xi�N���$s�|�M@BF��s(���]��?��I�<�g�u�͏�~.� PG�5A;c�6f��u�e<4���{��4����s�bf�Ef��T%8��;�fX��6���`[A��5���4b �u�I�^��rAu�F�s_�J��\�X_@;�5+F�z���`��JSd�T	djOC��X�џ��( �dSU\�L��k���n�;v������Iݪ�M�&r��V���UzU����p�Mp�������g��^�9�}�H�9��F��^��ˇ�·R���l*���O����͘���>��޼�C2p|�������F`3/iO2��ڿ�o͙��������o�ܻ�W<BIuԸ�UZaᆞJKĎ�RaĢγ4�>�L$s�α�C�����Wȇ?�H�!�Qs�ĉ�{�H�D�߲��]�����V@,[�\Go$�h�,�˨��h�:���*�?����ٔ��O��_\��&=����ܕ�ԋ��Lb� �[6�����l��p��r�z�Z{�5�>5�3P1�띗���h��\;>��٩옻����W?0�Q)��P���W�9�!AtA��Ud�0k>0	��^Ōo����[e�ґ���1_B*��L���)��������c`�
m�v��s���ҡ;2�v��5�pQЎ�dlm����9:�A��9�[o��`v�p9ZO��:~í[���p�^'����\S�6�ھ��!v�0[����M���I%�S�#�別���`\���]F�M������gwTYF��ͤB�G-I�_���#9���+I#ft��x,�Z��`��F�P'e�P� $n�a�EH��ɞG>h��کkZ���g�3d���>�e��\|-6���r�j�,�[��B��� 6]�ȅ���[�D(t���+T	#�s��J(.�!)`��^����#c��4:qtM�̑P2�!�-��(ܬ\��,�!du��]^�݇cU�8��)a��94��)�L�S�SM`f�f�ۆO�SB�]������9��݊�S"���������-I]�7�H���6��\�3�� f�8�ˉ��eh���s�?g�ل��v2���OW�}�x�Jݵ9���\��k�:�Ow_�#����_���qb�sf5v8������	�����,�Q��m�������;�p��|�h�d	:G4���?�ꇚb=�ӽ<���=N"��:��ѣ���$�����ZM�K<ǏkPZԪ��F���lx��n�pe�H�s�'k��XE�=H��H�(��j�Ilƈ���lzR5�X�q���(�zt]�b�6ٶ�%�\�I]xʤFj�U-)��
�����xǠ���E.�mĻ1gy�,*W��8dd�j{u��s��Ȇ���&�-���%x`kZȎ������8AC.��
��0=�:��铭2 � ����z��)�u����"�(�$eb9T�$�~�E��2��%z��C�z��4����%lJ:w��a�mb=�z����E��y\?��_8���*��9�6�,6��3��0@��b�g�2l?���i�u��8��S�s\��R7��ؑ��'m��K{�?ia�|ǹQ��O���D�w�,�ӻ�	h$zf���	_��[�9��R�B˯��Uma
�뛂޲��۠�S>��<���f��2hrcxD�����NZ��ty8�LU�5��SX�Q}*�t�!�~��'f+��Q=O�g��|	Ӏ+�٭-X����%�k+D��b�3Z���>�)K�pIܘ�ʨ�+ILM�k�RF(=����oHd"���n����v7(4\�}��B����mcJ���ͥ$�o��1.��+*g�.p��f��"�J,��W��*+���y����i�[LA�H���n��JvihA
{�2�Ɖ�L��y�G�4�q�N�����87��H�E��߬�G�#Bg>=�c�n9K�s�1��+ub��r�X �G�	�/�� 0��1�C�;�S J[�������0���Z����2ܣZUY�XEj��r��g6�+�䞄��0�>�S�:R�/2��xɯ�C� I��D0Ԝ`=�/ߝ����`.׉'k^�"]�TI���t#%WT�gˇPU�
�e��6�2P�ŵ�7O	������*���'���C}�N�\�ǩ@�	�[�7E�>�Ŏ9h�C`Z�ɡ kEE60���=�/�a�Sg~��վ����(eX�Gk���I��KAv@Z�=KI	ڻ�Rk���}�f�e/&d>�nx��p��}qv$'�A�(
3֐�Sw����ȧ7`���b�#��ðW.7ʎP{�,�#�Ҡ�c��l�Wő�ŀK?>�R�����}a�_�c�:&�0�b#�ֿ�����~���5Y]�)��0FC����j��pn0����x]�l�%W��_둆@p;�J�~`�k�]â�		hc@����u�9���}�v���t�0Ǻ�1J�1��eqH�&}��ZѦY�)�z��&��p�$��BYS<�86�Q�e��NvР�z�"0l���7<ק���ܚqt?�/EMY�Z^�^)Gv}i��a�Ņ���XFo;�o�T�h��&�/��Zg�����!f/�j���E�B�
��V��v{��B�<��/��O݆�@����mo��+��X��í�1Ev��P��ȴ�������RMbo���>����%�ͪ���]�e����!�cYq-�y810=P�Dm�!O1�fy�c�,o�!�8���g-C>c\s��ˑ��O�ZXL��H#P}�]Է�H���p�.fX7\��8}�� �&8P.����T�<�:S��fǚƋ٤�jS+�[� ���3��B�u18�^�Y\����I�D�/��!��za����� ��'��V^Mb�Lu�?j|�:c�o�x�^���}E�R�hj����Ovq�9*ʔYŘ���P�d�>N����U���Y(w��

���Q���#��C��U�!��-[8ի~Q
͸��uZ$�,+ҟG�yL�'9�?��&� B��ӄ�t�e{2�@S�a�g�����j|_��/;f�����Q���2���c��?�Z���1�~���K���[�>R�kJp)�#d`���B;���A����Aޖ	���#М�4�(T�S���D�sz�N0DZ�t�G�����8�N<�ɐv/��]�(�U����)�W�H�sK4/�'s�-$R��lS�Ԁ��6+����I!O!=��Qܲ�l�1�Ep-���#��RT�!7����W/�9fo�3�dY�8g�t�ji�
�P����R�	��]>�X����e�p�]�X��]�+��e�}(��ӱs�%]Ue�D�3hYT����X����/x��:f�qB "1f��|M��T*�$q�]��ˇ�Y����	��hu-���|+��P`�x�4��zh��S�EZM*��C1y�C�!�C�+����]'@��'I�_z��`�2��/X� n�1�Ф��s��h����(_�c�����t�n�P��h��j�}T��%|Bv���j�K�Fnr�>�Y�br���q��0p��!A�Cص�ۢ��"NLR.v�;2�֌jN��K�R�X�ᐝY0��ѳ���?�;�g�ѳ��{��
���W�#�������T����.������"�~V�ŋκF�x�(l�k�'��Yv�e=?���pg ���ڪ�Δ��&B|�;�袲}2���>�v��U�xk�0�VT�)�� ���R����r��� ��\&�.��h񬭢{Ġ֌](z�*�<:E����5�(��G�]�.A�d��6�;�(tJ���P�C?]�툍%�!^ʵb��@�=�c���ǹ_����I��ߐ̂p�&es���������nI�;�Y���<)$��,�Ejk@��s��w��851� e?HaKܻ2�/����U#Qo�,SO%�*�
L`����׷ǈƷ�1X��l���A�Gv�B�u޼��؍��P�"���L&(��r{+��`1caY(^7K@/3҇!H��W ��Ҁh�A�)��r�=��m��;�%���U�+:���[Wb��@�&y4�h;)���@C�[3�(�a�3�ϯ����s��<��Gj��C'Q���V�ն�>�l
bb�0'eY�Y�D~]:k�ޥ��)����i�\Ѽ��ڽ��t��
�a$R����<�'(�I���^��l_ԞS�1`�؊X\BK'�6����Y�r:�79�gɏe}��_��v���-푭��z�w�i�s��d�8�Ns%=f�I�Qa�/|q����]*�"W_GMN��T��)i����=`O8���Ϝ�Wc�U_:����b2J�11��PLM�����d�B��ٻG,����Fm�t����z����]Jj�?��ڹM(ȧH�k?��-��I奣�w���5/0H�[R{��M���PEP�9�p*f2�6~+�t�>���Z��J��W�X�Y�'��XRl�>#�qVg5|H&�	��N�����?�@��竩�>
�u_��ͯ:��/���?��Λ�>�>�-4*1�T��~��D�/U@�aXM#�x�9�z�Z�f�;����(@2�-�SƐ�5��b�Z�A��v�d��;$�F�ZL������@ev�����t��B |3��>���z��~1���U�r��wC��a&{����@��Xg�2����&h~F#L�K�
����;�<���V
C3K_$<��y��&��N�͙[����y62>��+�a7��~S�����S�T@�9��������~�?�����7roéu�ё��E-F֙X�A��%�?y@n���D���[D�M�-ǮD�b2�Jo�is����2y��H�áN8ڋ��LJ7�ѣ��Jv����`���,�1����s��/8�Z=j��
�y[�N�+H�g���. ђ�ȕ�bR�	z4����f�IF�����a�_���}�P�%���_*��*�*Il;�L��*��B�ϠP���s�"�>��z��k-^}���!uG}�,>��q��$q��X2��DY_�a�a���n���ƭ���kS�}����!瘊�	�F��Wf�Hǩ�QxT�@�{<G�G'���!Z�X���NeUdi��+X�$�K��3D�@���oوYa��4Ɠ�(�/*~���/(�ۍ8I���ESIG׍�� ��0h�i�~:'f��
���Ľ6��AF��9f6��˦�^sڹ-Ӫǲ(�<�/
W����,Zs�βrܚz1�p���.��*s7��nk
"/C����b����4M�_t� ��	r���A�|q'Z�?����w�� j��,�ϷG��E��R]�l
:�� �~&�܁gT_X	q��V�Σ%��p�QNg���~ο�bJt� ]�v�;�E"��]
5D݆��*tG%N�;Tj(�=��r�f#�̿�.��e6�p�U�X:M��윉�,�\�6�@�	j�� �O�ɖ�P/wA�&k��m�r-�o�i�@	,��V���W�	�ᡛ�ӣ�G��A�e��W�S��ΉIV�%��~��0��M��b���u�u� �Kx�V)��ݻ~�G��oC��ae�.a�U�.8�����X�Vp���N��]	6��-�V$��Kͻ� B���=�6}���.V揝ȟͬp�kVn���2��h��x�:KԢ��DO�ƘTM�wP��Bv������Z
�4��ISyC�l�@��x���M�$��_Ic��ማ��!Y��E���6Fq�/�&VV3`�;_�J�þƈ�>G�xX�D��wn�	���M��@�G���m��f��u�z���k캄N�fw���>���s����� ;`�/l��55
I/�i��?���W�?V���[���Pa+��&V�<9JpJ�Oב�i�������!N�ta�&�@���bF׾J�����|�!jV�����D��7lUqc�o��×� xZn�,<��#�ڮP��z�1�����p�
Cº�ZDȶ���Y��v�7���_�N��@���.�,]~5r�2)5�1V���-J�a�r��~c��0\z��o��2�s�ϨUsa��j�_��;���7�]�+���q����j���`DF��P��O�>�%G�&�f�L����,���Sq�6�L�sw��f�z6	_��c���'L^M����ف�@��鱌P�v��������#"�-���f9�����e����;�ua-#�><���ARG
�mz�E����� WDl��f�V/ d��(��;M��޺�p�����*^,�J�	#�F8q�| G���4�/�r	.Rers���SN�9�NK��o�T�3��@��Y�Q����~�ґ	X���(�ae�0�?�5R�N����-�iv�� J*?���K2A��1qw�_h�$b���#����-OG�"�G�;�ϩ���<`�X�^z~��4�y��􇌅2�.@zX����W�Jg�1!��j��u�[�ftύH�����}{�l}/���s�><���qg��b�24μy����˰�u����+sq����Ʃ��l����TLF}`K��~�xHtbӐW	��_���?�ؽ�Te�X���@m[U��T&6�� �;o'���3�/t��H��퉞}m5Qx�%9MMZ?\�2��.3�l�z9�+���Av�u����J��,�M4��5��X��gc�d$�(��}8}�����`�|�����Ψw�R`MT���8��dܘުɮ{�B���X��f9��QP��"�a���5?B%��	�vQ�%)�%�@+��������JN��J��1P;�;Ү��t�����ёS�+^�B�����$���nL
>�qh�m�b��Q��)K|�S���ٯK�i`�Z��T�s9/cX4͵�	���Oī�>��:x$�k�z�p�V�F����ç� w'���0�+ж^�b��+�K��7'������arؠ�`B����⛊]7��k f��&��r�>�2��ʕY]Q_Sf��N��ƒ�cAՈ縠J[ޖa��t����+�גJR�?�$+ÖY*ߐf���v�c�K2NɊ*\��~�ؕD~{4�����'&��q�T�)�b�C���h_PR{���ɴ�u����E"4������z�_�/�ҰWo�S��*��Ғ䎶�E�0�~�q8V��2.�k`"���5�)K�ȼ��\c��Z�uB�.l=X�P�ʤ���Q��ۯq�I�r<{��o-�w߂b���K��D�}y�'�;,�Hy����SA8��&t�f��!D{���J3r4�%�#�	?m���5���A�aˮS�`ƹ��*E䝦~��d�����c��.����P@����t���3�qh.��(d5�m4s�F�LwI�jp�
��=�G٫��p=n�u�(O�w���A3�I��<k���$,�R��(�����j �ҁ�%�&��&���뽒X�:ό� ��7;�H���wJ�TIy2�9ߐ�5�UT-˝��;�U���
�q�߯�7X A�P �++�[A��I�b��쬜�8̨փ[}�J�b��`���h ��x�t������5ox�4����ƒ�bSY��R"")���%?M:'�x�9P~�n�ߊ�b9rNG-���;�� �e"%S2q&v�T*���|䓑Za���_�K<��)VF�6�H�-��D�˭{m,Uv��Z5���e#���mxy��3<,fP!���l�|�=e*^�����	�C�,������8��������c��H;U^O��MK�y�N��\ѧ���Q������y2)��W�������`��,���%c��zC]$̳��4�r1b����ՒcR\���3�5�e9������ �M�ڔ�a�����������#�P|*�RQ�݃��-�gm�Q��[G�T�"$?$Og�L���5#��%��"�{1\M�^�(��0N��2�:Y�Q2�W��k�51��Hf
DP٬�h��+��iKE7�~)w�u�e��8�x�EȜ F���z��G��g�����+U~�ra,�B��0ᓦz�TQ� ��a��k��<W�+���$���ڸ�X0�	����I`y>b���f>�!���p#א�*ZvC)�<fFp�k�[C.��>g3�ڲ/�v���AY��x���r�����\XSw����j���1�\�<���k*�+��5n��c3���艹��Q&�C��\����ɗ���&��J�U���<�����j������M�&?/M�4�0n�4i��M��N:�F���
�Pxq��ց3�(�q�{S��R�"���ٜ����x���P�,�dsIt#§%�`� �}-�g��|v���m��ڱ��9�Q>0���n:���I�_�7�/�$q�3G�	��E���g��گ�kR��%���`$!��9]�\����E��2!��<����Rb;��9��N�jp�ؐ0�<���)5�UM.9ORw����q�Y��>3[p�_��s��\�H��1�2�䎇�F+��e*����)��R�p�i�PB�LuH뇓"�Q�4���׿���/�ع� �{�P6��nA��Ą{�i	�lz�nϼ�j	W�
!���7��%�-�@󺫙�\Xɮ�$x�1[��U��s�5ӱ���]~�f�6:e�a�t������dL���G��Piۣ�1�{����!�I9ٮ_�p(P�Yu�x��?w�ʏ.fv�䘣�~y�����5���~���(Fh�A�2�~�Pi���y���^��z�Fu�x�?v�e�霱��:�ԅ	('�̬����(��N�@)vZW"Y�@�(�>�ԝu�q<�u���&��x� sq�|�9=���i��E=��O��4?�%��L�ɿ�l�� ���L9�����{���T>�$EqK`��zǊ�k�2��y��������c�Sl��.Km�
�R�y������؏�I��|�/<9(�&w�6�'���Jp�?��x����e�Z�'<"�Ap��^P��@��[0�`%���b���up.o���R��J~e�|�I��Ǟ)gD�(M����d.Dj=��c-�R�Nx�;��i/IрVAt�JRV�y�Ϸ��B��5���a���V����]O����˖F��Js��Fg �n�8����������s��ͤ�-k�«C���k��H1�\ܛP+�����G7��Y����͕�l-°�m � kڀȜK�_r�ǰ=�˹�$AB��2��}�jn�71\��Wd>��B��ܿtR	dq	�����q���V���>��-^G�r)��1��!�ќق7�=P]�W��$/����	A)V���"dT��+��NJW����I`���,	��csR�+*0`�(��~�=����=�O*V:j�2�.�p��N]�+��/@a<S�<��ڪ��!I��W��3�w��*}B�H ��P���t�h�0���{�Ү�PJ�	�.��o�`�ud'`viɇ_��/�N�w�ip�;�K�
��Ki�h�<��6�gi�:����ţ�_�b���B~��v���4�<�O�ΐ��b/i+Aޚ��0'D(v����7��
$F���3)��f��	Pkz&���w�xOR�j�-��o���@}U ��BT �u�K��ꝭ��rڮ����jy��Bo�U��s������� )ⳅ2����1���a���mpLr�H:eq�
��ParVm�s��d�6��W@@{�J�YE�;qy=������ð^�P�C;�.Ĩd~����Ug�4D�d�Pʟ1m�x[�;P��%�V�r3n������������S(�c&o�~�tl4 ��4�8c��d��Ծ��ϋ�DQ���G#ZQzW��~�$�=���5W��@�A`�K艧̼2[�Xu�8#b��	��D�N�vPc�N:MR�m9i�^|�C�<$�7ɔ�.[����ঌ�%�0\����;;S�����k�?D����u-n�^q�5�̋ͦ�pLw4�7d�~���S�C�!�_����t�M�]��dh	�M��WQ�4�[d�?��<�	(O�}�/;��'ᬌz�	/�E�hU��!����y�W|c�^������D2#���׌��&�@O�i2�M�B81�����[!,�����[ADW�r�RZ�#EvA��_�eL��A9����%��.i�ax;�	��w��Q�:�Њa~a��yC����kqvbʚ��3�Q�t�]'r���,I藑n�"�Q�óv��Z�e�%讎=�S\�=�_����ڻ1��HWa��!��e�&�֣���L6
?��#�J��_׾.�rY�u fm�9%5�)�,�oou%Re�:2f���Zy�} �h��C�O�Ov��i���Y4D��ۋ#맀"�l8��f����@�s)���Lf9,.U/~S�Li� �4a]��������^|��`KO##���N?p��p-��&�k+�|i�xv�(�8�L h�;,����}u��""�sP�P��jf �C���g�q� ]���3�VV2"{~�cnUo�b��x+c���wIe���i������{oF,�=�!@v��"�K�?�ؙ
���nT7�"k����t�ge4'C��]c�#�N��p�F֒E>T�=����-�?���h1��?x������<ˋ�7�8�?���e�e,�����{|��<�ޟ����3��J)����[iC7�� �|�OFt@�J�1���WdUm�� M}Rގ �W3��h�9�G�U�8�A�])�
�})�E�1�jh�lƷ��ٚe.����R��[��d��l<�T�uz�{����߫�V5\�iMy���� �::|��j���$�-j9B����L&"���$Q6GO�|(퉰%sk9k�!�諳R5ϴ��m�&9� �d���V��X�bfuG�Y�d;��E��Uz?���w���M�g�8�b��su3&�F�l*F��ȓ���>3f��ơ�+B��Dd��S��T���U���Ʋ����j��Ĝ�e�����k~��.��:p� �t���������+Ld]����,���Ꭺ��;0�m��w���*�_���#z��>_7,��L�HM��`?0��gԑ�u�	^�}�˰�6a�k�o�\��^1Ǩ��+I���?���>������7�B���J� ��9Ց����_+(�"�n�����o�4�:c���屆�l";5�� sś���R�8)-75P*z��[e/ ���A�Ց4��:I��%�)q<��+��ZR�����'&fAP�x��s����V�u�`���J�VXS����DX����B�jߙ�A��;�(<�v �®�2�����(������i�d3�ZO��0S*o�wE�l��oR]�%Ӎ�Fǹ�m9�����9�>>-?�+��8Cq4]E)n�s�)��"ʦq���L��������I{�4�V!��QL :FS����K�	��\�$�[	].�1���<����'��}�1��_^i&d$D��0�����⩖:<(���X��ӱ�y��v��g��Xb�1f�Z+3���	W��t�+�x�w<h��.��xo �-.�u�fl%�e<���H����L��Y��;+=�e�����&C� ��\�����JdP�JDY�]U��Ҩ $P��a^��m�vn$�Q�So���$߬:����<�_FP@�O}��Ra��,�&�lռ`�M)���*oJ��i�mqã0�5j�3T7.a�ENXؾXj�S�bΥ>�����9���|tc�-�:��=�!$�gxe΃���k�se N"�Ea���|����˴G��Eܿ2R��r=Ȭ� 1��3Jj8*���q�ph�onqw�o��v���lC�eb���Q�xk��!�/̕�Jsf�W�KR�H�/�]��?�P�)i�ս߹��/a�YQ��ZJ�:�Ch#%hAj��_��g&�����Aߕ3A6�b�z��D�+`|0r���M�+�0������rn �u�a�H �����wqO�`��*�Zwkɜ��g�3��91/�-N�-�_�G���qq�}��ŕ�zZ�+zޮ|�_;t(�0�+���\!l�o;�e������Z���O�6O�uK|�8`�5U�J�څϥ�(�С,Ptw����.��=��i�&�=�3R�������x0�o�M��_:�qh�� ��Q0`�?�Ux}��5f ��@���*:�+�`��95~��9~�BR_)gT�N!Fe@u���(���7�m�.�R7����ۥ����	Hh_N2�R�����`,<����4�����z�������&�	ƺ�AK&�U��� ���>U6�hS�"RtK��,+���ɷ�uX!�X����O� ��0K�J���9)��B�G~Ƿ��V�F�9U#f�w�Q���(�V(��%A�&��U��.�:�5�5J��lZ����Q�hr^F�f۞*��(-��wG{�6�J�t�v�g�]ZG�����x��= ��b��ɩ����oJ7�<M#ϟ\gh�l��~���pR�_G�f��� ��D&�=1����䪧^Z9���r@���#SEܩN��X(��Ci��Y�r�9�YǑf1�n�y��?�-�}<���;��F�r@` &gd�=: �W�n'*Nu�4���#�z4O.��/[�2y��^�}_ ���f�ʺ<��l�Ji�%�h����hUjv4Em�"
_�փ���� d�^���
��)t��M�>�Re�M�܋[�k�{���x�+q3���~z�s1�*�Eā�(�&i!�Ei�8�\v�؀�wU�4i��A�j5��)�-�R��9`b�0O獈���1� ��M���+��E��]z:tk.��i�|(3���Â/3=���8v0M����
=�7�U��hFf�T��E���Ќ�G�a�za���i�EBS��
Ӱh��3��Ug�YP��KN5��|(N��j/(Z����D:��o�-��=�]*�zǌƷ*Lh\�
���?�~;l�5�O�]��9P�>�unۘ�۰�6�54�c��7��˄�ߥ6B��D�R]���y���~& Z�3�.w'�Q&�w�V�Wl�х ��֬�N�7���	��K]����S��|�K&X���κ���gpΝmq�ob���k���9���vE�������G� ��k�ꇛ �돶����l�ވ���Z.�(��ñݑ��v�3����Rk+�y.�ǘ���P��H�����1��[�@�u��Ͷ�n���w˓R���K2�_c�N*W|�胟pww�f�
��pt���u
2?����:د��_,�P��yN�����c�4�%�s�}~,.���OK�"�)4T��K�9�e�������U@6��_A�
#Xr�S(��mԫ�w���Se�&���e��#a�2�acP)Ӷ#Uo�{KzɆ��:�4�R���$�N޹��:�Lq�vql�̷	7@�� S}	�n�����RfD��Hp�1J�g6��a�e��I`��=��}��գn���R�&s��!�a��~���z��M�r����yӾW�u�O|��t�����/w`��䥩�*J.o�hw����i�lY2��Q? �����+Ԫ���oX�Eg����f u��.h�qN'~[���=21��@{%�D��|e�d�󐚷l򭣂z���m�j5+A�F�����-����-ʑϖ�l�F�SW�><�����#)(H� �3$�|C��y.k��@�a����5V�W6�$}�/\O��3���?$���$��d��*��'O<���\±V�5?15�@}?�������3I��=/� �S
������G�"�ź0��F7췉����K�xD����B����<��zI���a���SV�w�2L���KW{a⍥�{��7(�f+�y���(��~�1��9MEy�__��'a�_���x�n�0���7~@S��$�q�{���~���������W��[*):~�y�N6���_�;H� c��o��R�$ �[�q�B�Q0r�@��7v�e���[u-�U��~X ���hH��A"�@��"��Ix�}��Qݺ̹l����v�x�D�_����Zy*8S���+�Q����	sa��Ac�`�4?O�4�K�b�5��(�':���`|�$��Ee���d.7:�+YH�T�䲻|K6�e���?!0�FT�U1c�8�Ą͎ה`�#�"Uۢ�,_]�-zIb�5�n������4V����E�2r�(2�(���'�
<g�f�^�����i��!퐕��K�3ŷ�� ,�w�_4%��c�5~�'9H'�ɇ}^�Ca���3NOIY�y����W�"0���_�a�[��-�O�1S`�ai�jw����l��f����-d���Mt�;H��^����D��N�^ms��b��V��TI~���s�{�k.Ec�*��Ǘ�To�pX�|�Ł�t���	ͱ�>�!����\����J�P$2��fGMZ�	CFQT��t���\6Ɗ��Hs#�U~=�F�PF��>�)0�p���25�
(ϱ�5��K��%�S��J�����м�ii����XC��� %&��A\T�*��0�[t�B�s��\��a���t*t��M�?0��;H�������¿j�X�Ç5Z���SL	��ͽD*�g�B���3����g��ڍ���I�fW�H�b��JK2�v���-�0���x��겴餏��"��b�!�I�pݐ
���.y��?�:��kk�� M��+z̩�t+7$a��/�2���d�E��Z�oO|��j�]�I����)��>��A-�E��E�J�,�w����f�o����H������RFS�0��Ev�0`y���2\��?�G��Ke3�Ӝ@����6� ���ZRd/�:z��р��vk� a����h�s�Aܧ#�J��"Ey�&%�4���W�J���d{
;�Cdg�r�M���ɟZu��}蓋z	��8�2������_eL�����qΣ�����l���@��y�������2����/C՞��J�^�5�,��#��c,P�Hznl�5���	jȰ�p&�/��Y��r,��Mwa1v���ǎ��F&��:0b ��d82�3��-�� �ث��`?�0X�<������Z�>1��G�^��jfv�LY3��K�)y�n�J2�ֹ�c��(�`$UF�e*���-*~cRp~�5!XѴ�BdZQ�����e�&�7!
�^˘�$�wW�$��$�1-�ǛX9�Lg���{�������!���"K��}���!Yg����w���H�_l�5�����5��P��H�Xl=���<�4�ʏU\�8Q�b>P�K���hk�9B�(=�O �fōQh�|���y����`-���T)����s�_3̓�[�/����6�0e�Pͩ,Đ�{�b_`t���Y�7���*�tt�ᕈ�F/1�]�z7a��a�	��J�z�1g���N��(����-�+M�]��.L��\�����>��63N+��g�GG����ke�p�ܧT�Z?V�BQ}V4���x	���(�h{����nэx�aL7i-ty�by�45���9B$7�T�/hұ�oL{c�7��7V��b�l����Q\�	�F���]F;�S�
)�8�F�Q�@F@^��g��(��8�2�@�P��)ۗO��m@|X�5b���"><Ҟo{ݠ���JB[Z�.J�-�&,hL�uRbfMa�6�x�v�9;��|d�v�_�]�r�\�Xq�V+�KT��<Uu����礓���M �~,�o�f7�a�6�u��y`�3p�����[�w31\*�{3_��LlH�cg�e�gw~�2�xn����������Rc;���!��I ��,�-6N SJXᷮ�`�@v��	�1�"GdtpIm-E�P��{8<֩�Ql}�ۭ�G2r8I-���Y��8TH�F�?��E���5��N�	�x[B�3��������U&1l��U(�p��3�������k �Rˠd�£O��ٕ�����U�s�w���~�SH��~���]��O��U�u�\*����F��:)ϤX�7jgXՇrX��nx41q@T����ebU �/�\�ס�fvR#k�B�?��#�t�L�ծ�}���xm��7�c}`��s��<h�n�Kt�c�}Ҫ	�F$R|!Q�^���||7�Iŵp2KL�7�Ŵ����F:����]<W%a�(^��p�{�����4���p�D�<�J^�'$�TN&i��Ě������}1 �
�?������g������E�m��N�!S��Έ��!P�z {�O���7�Z�&I�4�r�@
S�?P,��4�pP����Ax1�ğ&Nߍ�L�%G@C���*����vxU8��I�Ф�sM0sܯ#�P�%�a2:|�tv���g���1�����^�^���E�Xld~0����&j��
���s�K�������F��ݚ�ߚ#��~��?�R�܋/���"����dE䘦���[����.�b�����l{b]RD���v�+ O׹8N	n_�]U�*v�d)=,F`ߚ�{Z��.�ؿ��O�e+"dn*Ȍ��r��0��dI��0{�	�0�y���Z�?������Ӆ6�k���l��rBM���(c�n�QӅ���{���y�s�Y�z�t�,��|�.qY?�RxDf���tԷ��_��c����uɤ�;Sr���+^�\O������	H�1-n��^�U��J���� i�ae[.A^]�i���[� I�Xϋ�N��l��<
(�{�ʁ��]f�A�#�t��B��qp8����o�Zy$>�B���J���r`�@V$I,Fo?�l���u�����;-_	�����|7��O^k��߫{�`��6DA�k��
Z�XTH�������u�X�=�4+�	j'UrcP��nϤ���\�ڝ��0�Z�AC�׬�5��K�2�/��H~�` ߬(��z������:Bϒ!6�V|Y �,?�5H��n��ni�� $�f��L,�x�u��9(�\��od�qBA���=^�[_��zgv�c|�L:�L�]�Hq`����!q���5���~:�^e�[�7��$Gu��-a�A�<���t�H�Lu	n�q_�*m�"�.�r���M������N�s@Ms�ó����o��$�d}D�S���A~Eiً��)���Ay��w�>KW�j��8�l/�E��#��U��������vv����z����s�
	MY/���-%���ɾ���P=:>��GS'�46��x�zP�n)ϸ,"�Uـ�����>��Q5`�����m�\��`��P�R�x5J$<[t}�a��7�I͵����D���Ӕ�1N���u�)>(���0�+��٬/�� �,B@|nOV�W�̬ЗMn�~T�*���ٖ��j�_�N�=_1���Ccn�9��9����T5���y*�T4=��ϫz��yQjyc��][�"򭁇�Lp$��-+Wl�P�Q>�FB��
���sA�d��xa*�P���Ǻ����#|��́���K��D4���\�X����%����E��0.�3���'��#D�d�Q�;ԥ����O�3���̺��X�uWM�� �n(�U4�qAo�p.��r�������_���fu��,2���c����5i "��ߑ,Sd�}���$P���er�v���b���"�N_vd�+�@�}���L+#1��a|���a
zp��?)�q��M�H�� ����.S������W����6C�F��'�5ROE��E���vA�WYO���?�n�1���G�c��_ͥ����Qn��u�	B�6�Ч��8�$t�Z�n5muz3�����^x]�y��D�גB�r�Qn}S�e��Pʍȥ!9hw%��d-�OPJ1��g��0������|R���0@J�u���t����!	�I�$;Q�y��8�A�g� ���w�+����k�K��gݥ�N�xC��Y(�z
f��l�>J�p���q�-F#��g���?������� C�z�;���3< ��=���?��{�%5�	m�����s�M�lކ��v.�h���S<&���"�ND��Iڶ��w��Ks�P�j� ���{��R�F�p�3[NBC�Q����7��UѼ2�٪'Sy�՟\���哛��1HHZ�z���u��SL�WE(	��xT9=&�f8΢�D���)��j �眷�4ڗ�x�u(�{���(P�A��m����V��٘����T버
[�CeV�6Ϋ�eY�guߖ͖�����>���<QZ"����3t`z�2/�8���2nx[��=A���Û�p>���f��IEyBl��.�t�u�)rd%DL Ye��V�S�E!n)2�|���Jd������Q\�KW�I�k�����d6�╮=mᕍ���߷:b���K�2b��k̮k�,s ǈ\�^-�`������3H
����ۜ6�"B�2VO�PRq�<�(=d^HfM��	eoqN�XU�Ya��h`bL[oY*�����Ì����#�ә�jǨʋ��9���S��,��\P1�H��b�R������+���4�(��0�ϋC�+6O��l��/�>��Mw
oC�����7u��k�z�~�f ���
�d?����*�(a���
�^��XJ��w��fY7GwK��6t�yL7b1c4�ŝ�K�d��$�E�D����Ti�!��&�*��XbYP8� �!׃���w �8��h�{��(��(Y3w��G��8�<F�غ���^��Κ�n&������KeI����N��\#m�Y�@�T��;0�<
#�+�d�*<Z�Ob�34�~���ٷcD!�$VE".�z�2N4�qZ���x����/ڮ�kq�D����<�~4��iɄQ���x�<�~��mNq��~�@-|
vo�{E)�Y�Z�B�UB�Nu�p A�;t�R����̢N#Q%��N�/���Q�O��6k#Xߘ��d�T	߲�Z�k3��t
�W;t��y�7��U;���A�[�_]����f��Rqf־�%d��_\�q �Nx�:E$�q����[����70n����ю���%��(ݫ��'�TEZR���Y<��>N���{+��b��le�)(��:a�ݨF��A��q�f��(r�zP��f�5�K�p��iۼ����Z����^��fH�9
%����^���U��S ��y�`g&6!���O��R���O���As��(l�;	���W�V��oS���2�������e$�+2�J���U�ܚ���(��k���T�		u�r%Ⱥ����K��.�g��e��F���R�RiB���3r"U�%xL1<�#�i�����	���iT8����F�n�sM^��d�z���������*ׄ%��>$��z��⦔P�k'SԯP�{R�7�x����$�^o����˂�;�� �m�"�̒X��Px,,���G��i_�^�Vp��lUO�1�m�����<�j�dAG�DEù��|)ϑ�[+>Wؓӏ}���x��� Q5���ǏڌP�X	j�$K#|��3͸�*���9����认�)�[�ˡ"s�)cx��<lw
sY�&�L����p���A�
�ͧk����ƇmFVd�B�9�zͥVu��X���T�#��4�L>ͯPڤ�/J#XV�BFuZ�#�f��s�>�W���I/�$�!9/L�"����R݌�����f[r�c�ȍ.�wL-t@��]���It��x�%�o. K,�K����8Ɛ3�Tu�3��}�%M43Oݝ��m�}��SS��+��-�ا�Eٸm�7�wqy��o��-����S�����몴��V��ƞ�a<�_��
���O܀y�\e/��u�΀bmҜ����F���L|����4��&ec%���+A�ԚK5<[���ks.��@�oSEo�i�/��Ci?�\=z�THOc�	N�zW_[]jRA;L���s+%#����+�,g��9�Nw����gD�
�W������}#�8gsn�ųv̍��������@.�����L���'��|�Y_�oJ�L�im��2ѧ;Uk�F�����EXy�Y:c	R�;����%��C-qe
/\�pS��68�e4�~�!�>+숛��r�xgh[�߁"D�+��C���&w�k��	�U��0B�n��`a6�����y��l%����R?��jH���C���"�[��3���j{�/���0IT
����-�F�`���K�)�2b?(t���g*����~s�#2ò����b{	*����̷E9éO��1��D�(�-��S��gza
	PN��m?�	 ��*�@|@jx��x>6Qˊk�m�%i2o�w��P��-e��9���RG\V$f9]}<���v���s�>�����eʹ���6I�\@��ޘ'�#Nq��n�1Bh�y����	!�8w�+?��u8/�ص�>	��q ������~y�&t�Ox��Z?%�7�^�V��J9ܺP$_vKe��c�窏���� �B5�ݏAQ���	9�,��V=k8�`~�;�F}�Cnf�8�5ɀ�Lry+x�qD쥔�JN��_Qh�Eܬu$�n׹����1?C͡}��3��c����.�o{�r$K��y���r��3.`T��k$�fd_��_Ml´�9�_ңY�.&�J_����.�zM2/70j�C�^��	@4��>`K�xny�G��~��1�pPS�.W��Z�;'�<���g�c�u5��Mr����C��8�����y���JPa�����c%"'����%߅r^�c�[D!��Wf��"�6&��AD맿l�}��	z�L�;�a��:]��vn	�T}\�c�8!+?�d��ѫ2uB�Ԕ:^i��IXN������,B=� �>[2��TR�eˏ��Mϳ��W<Y;)�3�?!攛��� J��|^w��L�f���`}�Q-w��R�RR�Q�h�k���e</e�F7���jZb��!��B���,$��C��eBNҲ;�NE`s�ڽ�<���,s,jcI2��e�r8��&����g�@�a�AA���5��5t���1�t:&���iT���i�F����(���ϕ�Id�$��08E�x�TI�1�׷�bj9n�8ޅ�|�Ǽ��;��"|6e�h͌8X�0!�J�=y�6L
�E�58�K�L�C|բ���L��L��0�<�$&��L�*'
��C*��o!�!Aÿ]�Ѱ�Vq��>�����H�e�3��p����BVKC��̳{i 3`}�R��;+�-����A�R��i���{4E�\(E�*nM���2��x���F��W�j�HA��&'qg;!tde���*f��Y���?�+G��l���,?q �30�e�s(qDkpO�iZ��O��d����VAV�0�T��� \&(o����6�:����$��Yݚ��qNh����@AP_�FPmK��|F���R�Б�<T�5;�Q���+�YL1�Ȍ�7+}m���[��H�&����^����!vf^���ȍ�C�P��S��XS�!������0�?x��(�M��a�KH�ت"p�Wߣ ��`.bT����Ŋx��x��ݜ�*5�R3A����ސ�-X��U��SC�'�˪�F �,{��0�:�}�0�:��vމ��Sb�� ��&��} |�ہ�p��Ql�R\I�GC���8��i%u'I��,�2S�����cx;~�����F�����V��L*��6����0Z#��,Ga�<��n��W\$T��W�b-�z��3�m����PRt2�`/�����7��86 �ޑ�v����t���j��n��Y,6��>�'�2v�5H�k�7�z��3r��]��M$�{X�d�m�~g�M��"���o.��*։e�㩳�S.-��4��i�Y~};�����j����؟a�g
h�}�U(�.ra,:oҩL�D�MXzm�J>6T�ʽr���,N�3�ε��{</]�����ȯ�"����5��o�	�
���Z������ɭ��Ψ�a�zi��j�A�]B��2����&�� wN�"�]3�d�L�Z�PP��.pno��`(����
�� �fʕ�uwE4�Eh�ܸH�7�daGIʾ����P �����\���ۄ'��ǻ��q>�xg�}O�3��^~����9k~��U�u]ި B.cϚ"¤5�b�� ���}�&�_�/Y1�.��L�#vo@��p��F��o��],s����?���*8PŇ��s�^plT씍C���� Q���.���_ұ=DO���!D=�V�C2t7���U�0�v�)psSsÖX�Ec&�0��������5&������@��84�w�|���O�pF6U����L��z	�%�bAR�3h�Ҹ����&v�~XI�o������8�^��*��;n%�=v��� ����s}�����?͑]��U��-�No@��G��@�|�����(�Uk���d4c�>��6L�������u�U� �o> ����s6=L�U���m�6N�/�{i;кAQ_��c\�R��UK8{�$y�G�<�Z��+�u@Z^���e>��&� ��ASjC���C*�X����\���M*�v=1���*{ۗ�����Y�2=���77P�1����u�Ux�>�*�i���g=[b���+�{�'��0F���}l
�v`OKɮksn��J{5�T�)�_�0E���?�/J|*���oo�r�'�M�{Rmz,0�^���8�����%�/7ߖC[���*����&��'�&�3^���_�G2�9�j������
�
[h�4h�k_U§���Q�aC�I�5u��AF��zn�AO޾ʜt�d�����k��p? *���/'Õ�'�X��nY琓���y-&�$:��/����XM����t�z`CR�S�w�����m�K�� O��SE���=� _�F�t��\����|b�xM�a�)1���vf߂��.�B�xz+�Eh��e,N$op\'t�b&����*uQȺ�\�e�OU�^4,������S
<]g�;�E�.��M�tP��\��h2�$�4�٭��`g7F3Ȋ);���y��M��0��q�=�H����m�՞�Oo�I��Y]��f�����7�i�6ڿYM� � ������J5D��;�+̭�E����}
_B��W�c�|M�� �RU'��~f�$��i~�P�mor�K�G߬J�>���]s�x,@k�)E#��AH�6����S�T�o��qTr�+_�>6��P�t�m�(P:8�_�{��3�OU���!�yrx�Ǐ��_AE�]���^##ׅ�bk��%45�;���c=N������=c����N����4��9�� _���K�N���+��ͱ=�R%&�SJ	�5��@9��F���q32K飪�o|� ���4�"��B$�-��Q�;S�CuT}�ܦ�]��4��_hf���l���)N���x�b�* h*
Ọͼ�-]�"��8�)*�j�ӝس�]�^} �a��uU�E��Y���qRV�x��TXN��8� ��f�����a�e�3C��*xr`�&X -��J�~b���v����X�J�B�$�Y� �s�t4��^+fvA�#uj剮lL��HJ�>�ݨǘ�,�9�;fRtD	���[����pA�n���6��\j��k�,�}+�ӛ[�"�m�b��wF[U,@���\ʘ�����
��Ly�����Fh����\q�gx]Va�Y��x%���Vv�[hǇ . ��w�S��wf;��r��g�L���a��ҏ������X*>����l�W�0ߟ�ꈑ�)D�1��$_��g�i�#�f�[8@-�`�|��CAֳ��4��$��0�k���=���<I	�OY.e2]�J�D��;��C�N���7�~��Q�����t�Wg�8��P�������]\3(�@�fUmQ@�Q�@h#B��[�(EP�L<��Kn?�n�Mq�Z�]�P�h��$[$�[y-H�k��(�#��]�6<@I�����L��զ4��.�����ˍ^l���,g�X�,�^��c��d���ª`o%)��`>;���s�"c��T�o�6$��[z6c�<�l'��������l�Q���A���ު'�-�����?���Y>n���{^H�5�W
U!%���s�����EW�[����!���9X#�d�����<h7�,n�k�3V���Q��ۇx�Ǌ(��=�-��1�z�؆���FY�߽d��eDy����g�	�8��D��f�ʚ�i�_Qs
]�����IɲR��ӾΕ���3?f���aʩ�tS��fo��S{̧�����������K!�w�w9(���T')*��.p���h]�/�9����mii����BʱR�U^�����*o����L~:��b�w+s�Y��;r�"�#��\Á�S}�
�P�`]2jh\����`���0�\����,os�^���O�e��)"ICI�uD�e�D[���$P�qT�ۊ��!�{%��yʱ�����c��I��o^��Da��Y����ˎ]'�RO9_B�{����<��(ue�~�H��9(�M}��l�����_Em�ֳ�����V�-��b�u!u������ǔ�o��e�n��q�ȯ\H���)���֫^k?;+�2?���OX�D�]���@�;+YM���L���Y�+=2s^��)����9�������hH��:�sN�Q���z�t��
#�����E5�,��	*0`e;O� ��7��^�0yA�q�+������Nj���i�J	wd�/@��IR��+ֺ��V���Գ�<V�D�0��&0�=�G�=�����,���3:B�L��]5  TY���(�Su�,b`���]P��?@�iS��,�#�	[ǭ�H�k����~��X��#'���ęW�K�O��e:W�^��FIH���ɑ�v�VE���\����A����TJ!-��d�F�;g�\�hb`���Fi��(LB�d�	˴y0�yw#�X=}ؓ�r�e[��<��YB"Ȁ�d~ʍ�0R�d�s��3���>�Vg0�f�������!l�,���R���!6(s
�WvX��/�<#~��_�2o�F.�C����$eM�4u-@��c�dp�(Lari\� �&H݇�\�ܸfw(��*p�rh�,�voC�O�}<}E�[t�˃��5k�]T�ET����L��f��!o����ޫ�ޏ94=1���^Ώ��a���3�AZ&!��c*P1�O�S=Л�a�@������l�/��Z,��u.1��ZŴ�,d�N�r��w�g1�^|��ʎ
ab��/�нԌ<�[�N��ɋ~��0Ev�BJk���wq`����S$V�#H�hjXNeҖ�&��0�����2��(ݏV�`�+$�O�Y!�+=s�˓E���n���(@2>A��p�H��nOz�U�߷r�s���i���P�|7�y�	~�F��G7�4�P�����0T7���Y9����[��1�ʝ����%Y�#�֥��Ԛ3��i�*p�g���9���,�%T�{h_��q�Vv��A��xv�QZޭ�0Ph�����޽w界�Y�&4`�&���h��bOw��8n�	q�Qq:r���q�M�x�ҴY�{W�(s�)�VaeOd	T,g�$ir�myꄫ���F�K��Mee�S/	���;+K��Nݰh-�k���!M�X�ץ>�D9N�{ߠ%���^?�DZ�_��բM�ܮ�������A_	0�X��T��i�*�L����G��7�Ֆ�ˈ��yDl9 ��y�@}�m�mo\IJT�q��X�־�r�+�2k�]X��
�T.�ܱ(�kگ��v����%�	������}�����N:�T�CXS2�@�eI)3�����������)�W��ˬ�'au�U�5,EJ��{ݱ�=4���
RP
�I�k���QE�I��vI&s��?&1ɺ��Ν�_�)K�i���^�C��8�m���׹(E�=Wj�-�ڱ�	�iJ�"|I��dW̌�<���P/MϬ�O���œ�NC��f�=�iȁLnw9�홹���TvC7R�G��6 }��=wl��h�����G���f��h�r��@����t��T-��n��:�3*�i6�CV�V��34S��)S���ӛ[���oD�'Ӎ嚨�[c�1�9G�S�U�L�DԑV�?q����g(?�p~b2E�q�f,�w5�:�VӘ�D��B7��ݰ ^�$%��un{�y@�m����Ќ�?��[.60��X�5h���,���Y*U����i��k1��u��o	iX����V�L*�}���J��艁7.d˸₁oh*�?�-��S�;�������o%�j���f�s�9m���G��ڲF�U�L+����6�8z�����n����l4]=렖p��31�.���@dY���#�%��[md���9T/�ri�d���xwI
\f|���&~�Xb�S��T��k6]U�s��Y�=�@���y��E�'��[+�i�ID�[�Bp��UQZ.מ�Ad筞��5.�����il�،7}1��#�3��RfZ��C�&���c:�`;��%V�⾎��=�t�]OuNS_�Xx��54MJ���D^k��UY�ލ�qH��f8 ����� �Ҧ+Li����(�U�a�"^�>^|:�W�D2�
z̠P�0lV�Q����6<�f�6��C�Җ��!%F�;3?ϡ���̗�����-]-���7d���H)�j�"�c'�XSg�_E��)��L�7�H,�N�:��X���W�"��ۣ�?��@1[������'o�_\�CSKA���6�����L�!1�Ё���2�4]{���问�MI� 5ȥD8��h�_�Ha��ĕ�?Sڒ�p�����{I�Fl�ʴ�o1�tK�k�%�}K��	=H}k=�E�Tʈ"-WĈ��� �¯R����0��\r 9$��@����}\�T$>K�?��ޖ?�C�Y�$�]2�b�5�!��"�L[D~*,U�9�Q��,u�H{�N�����({��0X����E���l��H�U����:�� �512�!�z9�td��Tag?p`����qO��?����Y��R��H�~�x"� X����,��=���VF�i{XX)�pY >f_4�S�Z��7K���u�υ��M���}k����4����H��Bz8�J��v�����.)Okf�����W�4V�u�k&]�xb��ۊ�� ���P_���T3V�;���0}���0��p�W�b��z�dM�I�m{`=.���X�p�v�Ç�u��%ʦ`�w���	Yp�a�aI�����}�-�W�!�D���yM`Ɣ��-��[��P:�xI_V[��C��.��H�j��;Y׃�j�%ӽ\�F���R��7u_�_R7±�cbӞR��T^�P�a1�iXb����__�M���3����$jހп��BE�;����>3$���[NcY-�;��H0�����`��(p����@�x}�]ɳ���=���Њ�QPXք����sVf=qGo��)��#w~�y����yol�t,�G���N��+|jğP,� �	�Hj�Ro�n�xH�;���&gI�0��e�q| D-�J�]� ����ƍJ��F��A���\���_�[��펃&f�R,O/T���;�9��v�=�Y�Q��h��J���"��C{���.�Ƽ�(g2�R&A\S�RiN4F.���~&�,P�cUk����t	l��~_L`xC�2����A[0%5&��>ޞ�*`F7�N�7],��5��º�-��c��!'�b��Ȇb%����F�o�=:4@�)����x�$;w�k3��fs�Zc��8J�򹻮#]����߄�\�<K
���A,�OMٵ�P��I�{�:��y&e6ņ����b[�m����W�j�l���KڢA���'HSB��t	�L�dv���Fb�8�Sr]����`�̗iE\w�P�F��I|��^�,�Lt0���١i�_�-��<Z���v�N�E/�_���J���/Cq�m�xy�����-F<�2�T�Zv{��cͩ	��C���Z��W$��^K�~p.S@�5q��x&N�C]c5@��B����&�����T&�
�ܤ�G*8q�ߋ��@$ O���&EJp�{@u?��9ۈ���ȟ����b1�d�2��i wKi(oCZ���'�,Խ��'1�V��M�@3�@g�ҋ�� ,'=��X��>S4ga^�Lſ���8<]{�Λ��o�xXcK�����#�r����V$RK}^��x�|���R�����?��3CVq��6�l�{�/(\�����d�������H/�\M�u�f�ݳr
�'�|�ɷ�n*��MV�\�l/��������#x6>s�߁���Ke��f�D!��cU}�EOB�}���Y(t����]��25Z�-��(~O��������0���?H�:\�m�lS!����{O�S��E�{>1ysĶ/������,ʻzM�����n�2���wf|����1 ����h�E�gqk��:��Z��
Y>z�A�.�a����^�w� }�ٷ�i�;H�Z�]�6�@q��g�Z�~�ݶu�X:���=�ca��L��¨�3׾2<�|�9��5�Z#%\��pԯmU a����T1�G����8Ṍ��^�*�n���!���4N6��@|��b��n���=r�"̣����yĕ�m��F~D��k���<�)!�bO�P�B�)eW�W�0v���w�mh犣H-;�6��/�\L*8��"=8:.V�Y|�T>���\n|����F-����A�,+H�z��R�@����T��٦��x/��)8~�;���+�:8������f�`�/m����2�{���ߧU��v�(83_���z���3���x��涒�n�	����JV���B���vPk8��q�8�x���rY��:Hl7�&�i��L����v��h�T�� l����׺Sj	_
h�I���u���k�7X3v\��v�׸������d�D���HM\I�g@/�P�roP�y�j:�>�z�����Oh�Jq���uT�=	(����jO���@6��6u)몆N0.<>��r/t�����߼��;Y�c�(���:��ຖƼ�ե v;���S��95�W&��ߍd���$}� )��Y�P�cH�Ӷ
$䓴�b���Srq�nA�#�������\������~f�E��m ��i��a�w�c]9��[��Y+�?t��{�Yo�X�%�Û2�Y��i�W9�4�m��H�[՝uR��tKJs���$�5H��A96	AcC`�����jan�7���P�/aH����FIG9���ű��J�A#�� �+���
ߦ�XZi��m�iM}��`b�::{��}T-�N�z>��eK�[#*����уS�"m�$��@��N0���ghQ-İ�JI��YX�!�_}h��^�#��覩����e!	v�� 	H��I/`��Y9W�����aY��;@&@���b5�Oq���¯�S�%�m�Vc�x_a����I���Ǥs�2y�zdu/��/%��®@pL�mR��Zz��8$ȁ��Ya��I���|�p6ʨ�v'�kʡ%���we�|U�s�~�p���[�G7x�,;� �rDv�2cA�:sz^��$���̗:�5<w��S�����̫{nwH:̋�L�g<�>�]����LO;�+� �KH�R��B�jU:�u� �A0�y����k�9C/E��*�l�(g�BK���/ܱ ���)����.nw������*L�.e����J����6�ұ��~���K�����(��*4ph[�ۯf�8�EHg?��ذ^)���]P.��c�캏�7b�i��Q��i�m|Pb�f��/��� mЛ������QY<6��+  �/��G`�D���_g�3m�S-�q�Y%��g��$2[��B���z�q���gr�_���K�j�6
{�±g�^.��-|)`݉K���(S����YRČ#�o���T��)<�R� 6I8�	�Xa��h�O�A����I�<|�Z��'lJ��d{� ��2?~ϩ��ϲA���?Mδ��m1Rq��H�G�'f���4�/-� �w���=��j�5q`���Gmx��[�;��]�AH�v0�ɫ�`��cm��O釋��z����:���G�?��a��0uӯ}��#DC7��}�Mj��	Av���lhA"j*��& .e�Ɯ��B��j�4��Mrq٘�%ԢA�8�]*�I��؈Q�c��ЦX�*Kҿ%%5��c�KN��Y�p�q�W��ԫ��ր�;�e拺6	ݍE��|�剋��-�CT_�_qj�vL��#��ߞ9�0!DgG����q�y�C4, H��U)]KP��?���y ��O��Ҕ<>�?�06��4	�s�!#�}��M�ݍOɔ�Mg���������Q��Hپ��6��0��&�>i��6�����*����N����q�g�eXǠ	z��Cz�B k�-���]n�[����j��O�N9AA����iEҪ�y��ˀ�T��Q��z)���V������0�k�������P�X?�|����,��t�jD�4�@.WҬ��[̀����|K6ҭnV,jK��;Vizl
mo�s�SK߸*`U��z�s��*2�u��I�Q|�T+�e�P��rEx�H�Ŧx
���n�����]'w�x����.���\K!�Ɔ3�  β_@�A��\+�;gP)|��tk߱�1�E*�\�F0x77ψ�2N��eE�pz|�֤:�L���_��ӞlO��W1�
���_kS��c��]c�H�<���K���� m�a��:x������{j�}F�e����lv1}4n.�l�˴Y��� sX+_��}B�u�R��1V�J�����F�ī�!C��H�rs����h���>0���Q��%`�V��흰�s�=ò7��	b�z"*~���6q ����/ɓ�X�
��ʽ+�����׮�`Tܘ�͕I�
d�`0p _`40K�zH��wI����5J&=���L�d���.i?n�����N���,�b��Fo(n�����R�<S4IL+�����8���F�խ*:�:B$}��S�
�B���a7����q��s��(2,  ����>���� ��2I1��K�1��8��aL:3����Z's��	�+��=A��9��ؠv��:���	�@�y�*� �@	`M���+�z�VK�
j�\XK��i�;��I^���N�e�|�˅��O��qᶷ�$���(��lg��D���7��a�Ƭ�:�vZ���V�q�����3Q�Ḣ�8y�A����P�	<6 *[��͚�u�O�������@�V���K�񊡦������]ς�.oQ�/,�z
$
ӻ�[B9r;�*hų@} 3ȭp..bq�,��9��� ����Z����>����fX1䣊�'��v��i��U� ֽ����+{�"���v��k�G[���hڧ��cV�bW���r��[�	�҄3ؕ	�^(*��~���<�xEa$�&�yr
O5za75�SQ��N�ԭϫ9�n;�͏��(V+C[�A_�j7�����@V�;
�|��Ǜ�mG�*�x�;���W�T��051T�2L�Sx�!���Ts�[�y��XXˇf��;M�3W޿`8��d]{w�mc(x�ϲZ������{G�BR�0��4a�|3ÿat���4����������1���1�_�,�[f��OX5%����J׷ȧn��]�f��s8.��ZHG	N��zĶ�[]��IBgLM�8�xV3\B�z�+u5��(�H�r�	�����(�j��b[��~�ޑ"k�q���2�@�ɦ��m)�f�S�~j�,o�%�z��Z$2�
���+R�R�jh#v/	�e�5<�^f�����y��W�_��w%0"���pۍI,���y����A�f��	x����`QͶ��4基m|���T�@T�y�E*�R�����G,�o�q�e�{��@�L� �=���]�hu�L�A��V����h�}5zUʐ��l4�F��J�;�(�F�+��Ps61�Dk�R�Ô��z�'I0�T�9W̖��������j0��S�d8u4��#����1b��5� ��"@�����+K��Q�ȏ=*ӿ�t-��}���^b�bIk�o%F��ֲw��OQjh���
��O�<�y%m�]�j��y�~�����6�_���~F0���n��($FT�R?ʧ���vm'��ڷƛ��{0V��ߎ<��������X�J���5��3yE6����2%���Ґ�'�dYj��9o�g�E�I�B�tŷSzҝ�z4!{5��#XXՂܔJ���$�����+���Q��mYϔp��kꪗ+o��G?���`U�yQ@��
�v�TuF,�i���$�Z��<�e���A��	��n�w���S߈d�qe:8��%� L�&]��K�������h�G��~_�'���t�nt6'v��x��!�Qr.���6��;M��d�Hf���P��D�1��L'bZ��F���Ņ{ʱ��N����{���y[E�=rT��V3��=���.��>sE<K��Y�3Dyʈ;���'�++[�m�&�B?���0G��Uio��	�J�Q�pk���[˶ 2]��'��$pR&
=k�g$2$�Lޞ��� �ǥ��z�Ғ�kg��~�m�R�ؽbMQ)u�Z�l�c&�%۰�U���'Dm���t�>�@Ǚc����-��Q7�ҝq%Ը 	��H-�J��\@��o��ZJ� É�7q�"��+���OlFT���"^�0����POP)�!��L&W���&]�+���5t<�`�S�y�{�R�W��I�5��V=����y���������Kj�HA�^���ԍѨ����NkPI(b)�s��ߙj��J=v��X
������=��D_.GIf� 1u�N�_K׉��'�'�=��I���/M~6^�� Ӑk�v��(���[8j�h�1�	آ�& l��{��P_�ķ#�c���/�q���,��or�(Yc���m&�|�ıEHJO����Zi�<Yd���C3N O'���N��\���M��� ���7��0G&���6H
���*m!�/��{=$��
�hI�Qb�UT:���0�
��Mt|�h��b(�%�jP�zG�t�ΐ=n��H�� � F� 6y`����Z3���P�͓��Y�J�o�Ֆ"�_V�E�����x�jÉl�2���<VC��¯������9�	�Jk^�EC�{E��s�~߹�t�O*���M�eԠ:�o=C����<�u!�G��6yw)�W-F��ꁢԡѿ�O�w�r!ak�!��s��1U�@�`�xZ�dl�J��x,rLW뉨Ċ�����w���5�[�a�j�^��0X�9m"��D�	�F�0�i`�:h)|n,*�3�r&�P��A������Ģ9�0�E9�`_��2M�|�W�����B�`~#�p:��* �	���t��)�j���apz�@�?Q�-����a��J�V;��B$�V���/6P6?&��J�A����|ag+�3�gq��.��Hn�hV�#%�b���w��;^�$Fyh<H�yMs�?;�2Ѻ����Ǻ��Al���hcFT�!Gb9*�V�֪s�
���%����/و��hF��"���L��{�P<�Zw�%3��N'�1�L9��]��S�r�ߴ�!�ST"��ڀo���>��|ß���|T)^�a�E��q���C�Td��Ţ:j���G�-\��zʸtq,a��N!��O�~���q��a�$��*�۶���wP"�x�y:F�]�#8�x��݂Ȑ��s���A��ӕ�Z=����-I)��}�o��P�����y�Y{!��iV!q8_��*���-��p���S<�~��-y$~�b?��DdkZ(퍨)��k�~$F�*҄�%j3��P[&�h��h*�I���S���(�c�u�|������(�����$��C.��L�=�����/�����.(ߡb0Ҥs�";�("�Q����m���c�{��\����o-�!���r�����v0���q��8�z�;�n�m=�d/�sFf�J�'��~�?b�(U�b3w�PbS��W��v5���:�A�Iu{�#v��p�i�_�7�F�m�N�ս���jn>"��<��/�=���g���7�%������}h_�dS�W9�3o�%�gy������\~������\�u"O����V�`G/�R�d/]z�D�����+���]�y�"9�?S���H7�(Ro`���s���?Ж�F����҂s�/�$X�y�k>}�CיRfc���>Ni��j�|���Ɉ�������{�f��./��?s�@ "]t�*Q�����n/�)&<��ܹ�`B�3�L���>dy ���:��3T�ذ�?��-m�H���D^���d��m��2�i/B3�kBB��{�d�.��3:9yF���!��;h2��S(N��2'�UVL �^<���sU�'��6��G=T�9�:�G����6��ǀ��]��!��J9髈�TYR%�l�����fKh��w(聓���7[��*�G�����H)Xa�m6�a�w	:-���q^ɗ�o�o�	4�`9��q3��z2�L$�'v"v�A����B��Y5�Ѳ�?:�n�"�l+A��z+��l\ͪ྽/;�����\v�G� ��OL�@�!�1�p#�P&%`�J�J����J�%�%~Ð!�D=��1-���퀠LDA���/z?{y)I��)���J���V�As��N'U�e�[38la�ɋ�n��YѪ��m���P�ެ�"%G`6�����ev�[��),kфS�{� �h�Q>��E�Du���U�{Dc��/�B$�d�+B|ltC���wG�p'P<~���]��2��������߈c�0��k�B]+��	���K�u�p�gw��K��C���({SE����陛��D�a�.UҋN/`�8��t`@�FҶ��;m@�����3`�]>�RV�����hL7�~ֱ�t��:�\fߴ���� S�XU�Й?>ډe�	��S21	ZS-�b�R��V�g�S�m$'�h�ۍl�CUV�J�X-��&a3|��t���c��w�(��efIt��\����N��g��u����������tꘇ���.=����X&(�-��C(F�7cI�n{���a���g����� 5��~1+��o01��ҷ�,ˣ|-
����S.S~�&̒�V3�D-%�G��W�f«w'/G����9�Ҹ�d6zĆ����W䋄"���&	�<Kg���`�Nv�7��
��̫��R���	�uk#0N|�X�؂�&k��r�u�?�4�TP����DU����bI2���ȷ�4��S���G��s|�<z�(^iY6Q䆸�3�z��N��c�_�@��iS_��
n,���r�R�lX�J��\÷2�)�6}PVb��c[�b\.U&�
�InCK�������5n#1FAJ��r�{*�Kv��S��@H�ԧ�eWx3���9]h"�iZJ*ݳ����?e2L�mDUhU���^i7�Lg����''xw�)��c�1Vl�w*�CqtN.�O��RT���F�-�:��ϐj%��S+���N�1eM��U@��1䄣��Z�{g�ݥ�����(�gR��uF�1X�xհ�k��R�5#�����@��&"�:?m��EPL��n(�q��]�)�-��3�t�uZֆz��j��x��,�"J{��hc��8��s,�/���8/�V��*����h|충!��h�P��f��?_ϧ�n���|��`<����ؓ���e��}|z��y!r���߅�[�\#�-�j�*��ř|��D�F�o�ȱ�]�E�~��7��_��0�%���j��T̰JH�{?$i�`V,aG�5#�S�Pg��#?�I�����zS~���*iR�6ڽ3����l9ƥ�B�u/{O��c{�B�F}�$�'#Kz�ԝ
m��A���[�Ʊ嶜B,+U�g��.뱠qL�[�[ ��{�JQ��R�WES�ׅ)E��{G�=o���盐% �Cԩ���r���r������ư'�T�ږ��I�`��rS�߱~�I�$�	���8(T�]���%%U�D�\����ī&GP�j./%o��J�}���%v��p7�1w7tF[:�!��Y?=�Y���ٗ`B���}P1�Z_ ��!-D<�{*������5��H��:c[I�y}d(�-�!
���w�^Ѓ�_������G�v�+��
��� @y�K�4�Wd��<_�r� ��Q�-�b�H)���JtG�P/�~�>t.y>�o6�Ұ�6��� �]���Qf�=�c�*�PO��^ 5�j���vܐ�@�W�Za�3.���Q��*�8���+�9(,D��d�n\S�J�!�.� ��x����HY��������OZ�d��x�OS�g�L7P�ɳ����#��e��а �Q� ��_�Ps�ۺ��Y~�iX����+�x���^3J
�u�����/�ݓN1��a{7Zk:9g�`P�#D��mN[��J�կ��fQ���$��.��	�������j���{fg�a������m��;O�s��F��j�k�ț�@�*�DSڽ�D�ȹR�b�{�C���6����!����P;z�q�A9g¬���ڣ�V|�]�b�Wڱ��u��b$�p��L�F�E]��U�O�u��QM_Qq����H���PWl9��3�N���M(4�����B����K�����B~K��(����=G^UC&�����_G�5H�e_��"�f椇u�n5�7�p�X�����?�6���l�1�;���Ǐ��m��~�t���0��;]}o�P����u��92�@v�A3���O?Pl O�P�픺�Ȼ�Q�f�L�|�}�$M�
�	�.怛*����!������<���)�lFK��B�:T3�c��oY9;�r�%�W����y������K���W02�n����+I^4���L��5��.+y���fO���_
8�6@/e�VP�_�iP�� �5�,����0<������m��"I� p�m�"�bٮ���dd:)^��G�q�[b�oHh��CB%�P���U+��{O��I̪l���>|��:	'P��B%�J�p�E���7=�6�~k�*�c�^;�U~ M�*�^�d#��~���kC��x?v��p?�[lTn[F3�`��J�ڇ�KVΩ)=C-�x"�Uw^�3�I�(I�N5g��zٮT�H��A�'��.�������BB�Ӂ���\����ٙ��#�-_���;d�}��2AӬaW*~�Ei�2f�,���;&��6�^聅BM!����j	{� 8Ѩ,m�ğZ�9��RS�2	/�R#�2����:���܃���4}��������^]���s��M�(b#h� O�4��D�oE-���,���W#�-,tQ���F��X����Y����Oy���yZ�6ˮ&خ	�Q�*Xa !�$���;��F�_���n�(!����9�`�ɈL�W�Iխ3�o[�PO��qS�ڭw~��Bem���L��\c�6ne
�uމ�5g�ߴr�[b���3�'`8a)��8-����b��O��5q�:?s��k�%��*��H���-�|�H�-�N��v�v��i�ᧂ<b�5菦<T�]�9�҆��<�`��{�i/��%Z�榷ÝJ��@�ީ�nޜ6�V�k��'�^�fܨC�	��ǉ�0L�a�BI7:WM��Q�/�f�d'tJ�Z&-���!���UTa�ܑnlߋ�w��7j��؃�tiR���� n}�-��n�$�a��v��RG��K�ݕU������W>���8tȽM8 ��8�?f�a��f�k���tz���:�*�O����h��������A;͇�\N�S���]y�ߦ���GI�yڪ��Ԁ���n��kh7W�#�@���,���wٌHEO�D�����/f�����,�3A����Ҥ��t�'�|����*o�����EY���)���|o�'���d)F�h� YV|�ȡG!G��H��Y��2���d,��e�R�w��퍘N
OVA7��1��351���X��S�ҳ�"�Ǩ��Ǟ ���+�`-lCݨ#�Ǫ�mYUa'�GA���TĨ���_�Fv} 쿱Fx���>�9o��dC�y�H�N���ԧ� �4ݣ��s�0�p�����ξ��HK)�h�~�ʜ���jb��?b���ztT�Ʀ��y8��B�cb��v;&3˩��u�!mD�9*�>���!C��84�A��h�|�p���k���W���\��l�n�W���m�Ɣ�^BX K�1eS��L����(\x�����?KK�G�!!�Wj"w�q�b�`ݴ��@i�a����, ��P���D�dj	u�q�f[H��q�8(!�D+�ݡr��|���s�Ą����}:�O��g��p޽�;&
�z�*�`�u�v�~������x�'�(*y���y���ew�DV��!�S/�����[�ֿ:E�}�9�r��o�c+�Ib����jЖ�,�|��:�����2Wz��g����P`��θwӁ̎�/>��V�H?�9��(�)��fS���Q<3|�E�u%^����$��u@�86���^-���{DӦ0
�z��vQ�!�'���yαz	'Ꝯ����'���V��Xc�*��0��G_EN≑�=�Ƣ���7��A�֫�BP�R��\Ɠ�"�~H���q[����"�0�"
����6�1�����:6�UA&�.�37���q5�J���&f�GGB�?r��S�vm|Ս�m� �N ���|�\?�mbc�.��������5R>';Z���<]<I�mB���WQ�9׮ᒧg��~�yɝ�=�W��ǟ4���jL�	�Xi��gyz.:�//d޿� �+���*�G�#���z���̏�}��mw��+�`��E��σǳ�&����L�(2��X"�"�d�KA�(���%7��"�����#����;��y�`�{����Ƽ_�QT篥�%�'�q�
 ��>N,Έ�&Z[S,Gۨ���ERL�u}�؊�JzS�:i������#@���]�;���R�ʘƜ�o���9�y���~��
M��ځL�Dyc-�v�S��$&Fa~�;\��[�wR���&�'�pX�}_Z��Т�?� ��z��K#��Rd�Ï!��ߌ���) ��B�7�##���;�֬�=��$��:J��/������k�������M�7�G�l�
Z�����x&��K�H"]#�O�?6U��#4/��A%/��N^Y���U^���L���ў[{i_��/�`�t !�"x����Aeܴc�T�r�2:
��:�v�\����]J'g���dun��H��@�#���$�)=�����eI�p�8�y�?�q��9n�@��ۈ�AU)��� �&@l�*-(����eIk|�M�m�Y5�5�r�w��{�&��� 0V�3d�'�_~d�P$��er���3!��z)R�D�.��k���Z�y8��g��OAL���d�T��k��q�����D�9�-����ԍ��f|���`
.]��'=d~��D;`��a������L�sB�6 �6���VM�<j9�Ŵ'�jX�����,:��=���߿]��Wu&4���+H�M�39���"��-=�v�o.�~�����ddI�
�R4��|JO����i���^G�LC �OY�@���UrP7A)@,^~}�R��)BAC�8d�-�$!���n5:H�(�|&����3V�G*��q6�!��a}�:jq�q[\�r��0hQ2{���خ��-�#���u��V.�{c��(�e���fXT�C>�U�<�ө���c']r�@� cފ,�����ʄ9����}}�8@nd͒����f�ƅ�@�S.w���36�_L�/�qu�N�Y���D+z(
q2*���C����{c_�m�F���?�I��v4����*�t�yW�;Bͦ^������1\���ȭ���)@%X�R�,Dt.0J�=s���L�Z��X6���5ʮH���E��<t]��N���9�u�Y�R^M�@4ѼD%p��miv�$�O�7Q�Gs�s{PAC_;at6l�%2�����~y�R�Aw��>��84x�6�
("�T��J�q�F�� ]�̈́PT]B���\̭�C� ��E'��(T�Y�����v�_��>��9��ϡ���k�hz��:���ce-S��fp���	�F�F�]�i��L�*��7tĴ.�Ex��ߢ��X��m1^4gF[KUQ�蠬!n�����?/s�,���ύ�֭迗4hl���Ө�\qQ��<�����~�ܽ ����˸���Цn�Ȝc�$܄7O~ �6�&	��O����<�*I^$����#��1lkA+���!Y��
�9�<�q�{50N���fy�ߜ�DL	��KK\"Uyk�YQʿ���j��d��a1�։d��F��̪
){F����'6u�Z��)��jՏ�a���ʢ/�u���
@�ŭ���{h}(�z��*�[�g�B���hS|�BD�(1�k�L)u,�����W�ƶm;�c<��>���������P�|��M���mh����=p��T�t|�8������	|�H�N8V_��U�lu��S)�Z�����`dU���-��4�qSu���Y���F04���Y)Jr�,���wl��ނ17J�R�V��ȅ�E�B�"cn���|y��L�pl6��ܜ�����->�*�sC>��|c���\t؞�z�wK�U ��J3�J`d��ԊM$�^����7T'�j ;��X5{�����'��A8l�z�Y��n�[��p{�{�C�AU(���¸������Mw�Wڪ�2E-:�/���ui�\���Ρ��E�k�ߒ�3g�5z��)��Ǐ{_3��㝭�7x��d�4I�+ �4�{%�|J΀�>��k��g_�ۚh7�K�I�lh⑵��ϒ0r���<Aq���3��Z�����1&;ƫ$���:�D�	�&�~�6�����q/1~1H-�|8��<���]>��YC4�|I��կv]Fc����W,�����KRT�[���g^�g-	"^^�͆��.����$i��ԟ�ւ��Ii�wUy3��gd��a�������֕��8�7\�GȮ��/��d�/��u�B��v��|��ƣ�W�%?�	1X��P�$�|�X���goނeA���$�T�b��o�~u���3���i^eT��nq|[ӽMV�mj�X"K 
_�^�ݐoqF;����/��U�WB��@_��ZO�Ϲ򵰑�P{J��,֜ ���F���·�.bj����u:�x�4�����M2Az��r�r��f�}3���\/۹�����~��-��@����M�+I��0$4J����\�$��|����U@i�lъ���A�[�<��*F�O�`@�=	� ��'����^p��#4q��d��Η���Rs#2I��dv�40"7ϡ}`��ѣ�=;�Jg��|�E�.1��Vq�GP�>jC�z8*����[q�?S�<��|ѩn��Y�y���DD]�6��=��g�o�\~u>X��vތ�"�Zp+�A�çs����A�k��(J�0��Rt�L����X��ޢH�%g�t���?�~�3�����bm�?R4�	� ���K[��y�}A�$2�XL�h\$v�~���jW��\`�m�Y"~�܀�6�|x˙����b�EF���H�5D<HX\F:���;gI�+Jp� �1��[�uKUYY"�s/!�� �Les���8wI�~����n2�߻�6��q0�k�e�"\���\4
r����l)�u��L����g>����u�)�D�6���0��{�$ے~���5����;�$Jq��OA6���u3��zcj���������D�x$�`ʭ�b���p�A��1��rNy.L����<`J��ܯ7F�}3��3��!�ƞ�s�+�����^D�f��^�4a�/��ꂒ����S��K���lG<sUM����j�q0�0��Jy��z``�J,b+���!���ԇ�-|�#���i\Ե�է�9�(W���S0�1W��Q�R�d��I{s�YB�ܗ�2����}s�À�^E]D��8oS;��?�6�}X2\�k��^܊�[�%8�B݃;!����{]�C��R@�a2�Z�d9J+: Qߧ�C�=u_R�:ur/�����z�\k��l��l�5�̃]v�T�C�$����:�W��i)�� @�Qk��+�FN��<�g뉻�-j��N���V$~��`뤻AW��-榔�'O�(��'�MƠ�yA��+���8��o�5Ew*�� ���A����	�"�r�:~�"�����¤�u2�s��2P�Q��5;̿��Dp�q��k���nl�(NK�X��]�;z�f�Va���e���/�!pF$k�8�_5h����s8������S�bhE�m�x�Xƹ�5��Ϝ�#þ	�b��"��@,0�A���{��+J�@��lV:���[G�!�`�ݜ%8c�N��N1>!|&5��� �i��!����A�3�wa���8eUX���lo@j��͖��,�"#i��e�r]d�S�J��=���f��L"<rx Æ X4��r\����cwB�4�����;0�4T!���t�8�3=!�'���d7<���YRY{^��-E�{d�|Ω"�5�ћ;��p�o[��]A[��8Np�9L��`lv��g�����=![('��4C$Cp�,Q<��-��|��-h��
.$�����|�}DQwn�R�w��e��Nr��T;�5c����(�\�}�7��=�D:�`X��O��R楗�n]�U��� ��^>BNV6�gʌ�m� �s�M��;Cju.�/wp���eQ��;h��0��e��c�6�5��W�ZG񨮌�u4�9�Lj>]��<� �ش�$����W�_��mX���&%g?��+bK��Y�H���K5: �<�{[�A�6�p � �����������)����� W����s��mބ�KFu~� S���Y�*�n3K��랑x><�+yN]�&=�+u�<vk螚( �v�-��-H��[_�J�/��h�Ė��r��Ϩ���Qg��V��!�WW��C	i����Y$�6�3]�*���S��JB{��ϭX(R�گ�QU������,��V�\�}U�T�<G�k%�t�C�+~7�H�����"�}�j}���tt<`o�$�Z�GZ��=������X�A��cr�K���&Zi�Ƀ��<.�(	�8wӨ:���L\5��)��;V��޷���10���@>��@g�<�X����GZ�3{W��>��UE�Z�e��Lqs����?k��=����֙:X�)��*p5׭��������:�_;���q,�=	���C휄X�ЇP�sit��Q_H��8�ݧ�թ�iI��p��M0o����
��ShB2A�^��k/�ԥ�����  �D���!ŝ�PZ9�X��m'B�9�_^35`��;�xqc!��r�c���H4���brZ<�b�5ɴ�SLGvI��m,.U�+���O2�������n6 �J�v�dsg�y��H̭j�a=�m5<¸�������c�H�~�L3B�>�	�7JMp�t8��b�3�+�R���� k���v�P��W��љ���ނ,����Ły����mr��ه��v9��
�~0�L�߇Mފk��¶�mM�x���T8j}�x��N��.�ţۤڠ����sI����3� �$|��>W�h�f����;r�(Ӹ��Ǫ�>��I�ؗ��}"f>W�LZ�k������O_ԟ�	B�Ȓ�/��L�R������өf��]�� ܸ�y,⢄�5�wG�٠��F␧�;�@��+~�	)S����v�6��WD+�<µ�w���z�6�سN]���\|v�z��Ҵ\KBG���'rKl��,��wڌ�(u��dM����#�ۺ�o�|%6�1����vRm�۩�l#�9©�}�_�-��߽��Q]lfT�W�E���T�W����M"��r�]�f�N(ǒ�UK�tP��;�KE���ԓ���]5vk�\`�i�[f�ۉ~��^)2p	�� ����1�H��<rn���"���G��˟:�oƛoK�)����.RTep>z�ܧax�27�O*��5����f	�-��m�ǒ���xI�TUV���T�P\��3Yq�Ee�3;J���	w�65���zhNP�b)�HMʑ�7���:�+�.�ά��:�	���eU��~���o�W����D5a�������e틿K#:�VF���LZX��q_ji�j�۴�9/"�O�cLZ<�=�pid�_�#f"f�)�JC��v��h��4���ڑ���J�<��U���b~o��gݣ�ś1v�B��\��W4�kr���\��X�wF7�m��vc锔3C���sĠ�(�/-�ۉ�+�A�:S�vr�X�R�!���!��W����wX�G$�bVP��������q��N�cC=�A���= D���%!i%�������t��A�^^�7����8:�~�f�3�~�#͙��<�Ƈ[��Y�7��m]��g��.����wi�>�U��T|�3Ui�'�ӵۀ�@�樞gy�%²�J��fa;T���o���N���V&��VT��ya���qSem�*���}"���~J@%��F�;	�9�b��b�r�~Ң��W*~j�iuRw�8fD��P@J���*�hJD3>Z�?Ȯ�cG������D�=CA��x�B[X(~-ʖҽ}p)�5��z���֊��FP^\PQ��/K��d��W�����B3]�	6$��>S��M
<����>g�������-?		>�hR�xh�	�o�]�p �6њ=rDk٢V˜]*;2
3p��KXO��v��D� ks���n*��X��ylW��T[�q�W���๚\Y�/jI�B���l �����FDX1M||�5��ǹ>��s&\IP��g�|��
�h8X�t`tY� ��<~��!�u�h���,Y���=ٵ6C!�;k̟c?.����3���ab���op�YML0.8��1�Q�ԟ�hZ`=�9~++�����ps)���� ٝq[����B\�8X�`c�������\����ѳV��݉�~M�p�� �
+<6?�KQBY����!��V"��7�P��f$8 �٦�,�')�dR�M�nt��� ;=�]_�P4ߎ�42���P��/��uG>����-���1H1��%ۅ?�'� }0�n�~�5c�DR�'�3N�7.��E'��M�<q�H�s�r��Tf3!�����_�N�,��  '�d���a$^A{�djGe�39K�'X��3��7T
��Ҳ�n:{�ɟ��1�(
,d����a <ȏFd@+Ͻ7CN