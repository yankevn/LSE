��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v������� ���6�\?���������b��q]�rf��<Q fUk�â����2Z��)����UU�1��� :�^8�U�	�|�E�$��s�&5�?��w�2r��K��\�m:7��6b�r2��y�g�T��C�(����g\�"��z �����'o�/���F2�����|U8A����,����u??}x�|p\
���Q�A��Jp4��D8IWȝ����pD�S�GbP[���ݸ��3XN$Py��>����\|��R��W�����;$Vh�"�F��Yq�π�M����h�_�{U2UM.�r>�Í���`�圬�m�Hb6�%�`!��c8 ����vޤfJ��r�(���/!*�m���ER[X�+1Hm�9r�/����⍩c��[���w�<��I[�CrPID�~�]���-��{<���ĂhY�I��ٶڿ��^P_�p�<O!��&��nqE�	����]&vP]|P9� ��/��S���䪯�@Ktf״ϥy�Q��S���K�\f��!�4�l[r���*����g8��#ǒ�\�_I` ���n�������ꡣ�T���g��%Y��Օ4#b��Dc}s���!�F��/މ�T�p������	,�)@��*p,i�oK�HD7�ea�k�a:���pD�t������[s$�A*�!;�f�Oɾ{�����~�Y���z�k�d�w���i�l]�O����(A*ř����Mn~��N~3mX�^���T�/��z�Ꭿ�����6��nɴ�1G����n��b��|Eq0�?㨸�W�Lh��A�����Ee_�钀O�}Ō �S�Aa_ ����_Сo�Z&��/��!4��9��\���'U�1��m3���!���1j������T웿㶊d�ٌ��W�s-2�G((z���.����S&Nq���Ö_銰L)��C:u��{v�o�=�@�WD�UIW��_�#NЖ���I.��4��!��F=��7N��1���C�znm>�4��3+n�-)^_��#R�܁�HbG�n��'"R���Yb}��*��'=
�+d�����J��,Xc��ýD[�� ��(����O7�air��kdH酸A>1 `d��;�QG�c��J#|�����Mr�7�z\�ق�,6D�T���
N�����'�`0�_T��'���*���f�i�Iiˍ8�h1�a�qIr��L������պ���ÁT ?���%6�&q�����D�qFw^��i�d�
[��tAͅ�
?���,%s� ١�O,/���J��&�S����&�,I��S�L.J���=�X?���^�����*����k|����4]V9>����i�=*������J@��`B)��F�5��x�?-�3Vc͖�Û�K-�����\�ő�^^��;��i*�У�kT2��P��#e�%���aÀ:�l������h�膂#���񸫹Ǿʺ]���~Gkx |LB�&�
_җ�!k�1�Z��F��yZƌ�܎��i�V�kN"F�� �o��+��w]1�Aԏ���=��9E�D����!v>�CᯱOH���]�u��am��Rs�V���͋�%؝�]�Q�0�.+©%ɴ�Y#�������jr���8�3�$&Z�o��kL��:�;�D*�m���JA��� ��H�I�`�������3�󇜁S��Œ���tk�4==�+�Ԑ�k�$��#���?�e�|��&�.5
���X����s��q�ä�	�z,�!�:�Գ<�`�}�߲�MS����t�aoư�l7���=����������2����q8ۜ���������u�:Q���?3񢕂z�=7�b)2c"J�Yv�T�"���$r)r���ю�Z��	C"1��ޏ����e�8����Ys�x0�`���G�Q/��icb�x��,<��U�S'�\�T�a���.�� 0������Rwh�T�J%�Xꗤ)�z�B�{�ZD��R�/m���7�|H~����I�Yf�,2���s�-���l���gT샯;w��/��D`(���t͂���~7(p��#��5s�H�Hff	�b`�?F���'��'*��]�'l�9^��H����(�����[���0����ԫ�-��������k�ͯ�����&��*��(" ��?A�c�V�-,ԃt�ъ��R��+v��B����L�"CM`Q�Q��,��1�����T']�/�� ��Lcg�[j�]D���-{�+^nȥ� 	�8�G����%��6�������w���t�\	�zC�:>N�o3q>�[�\l�:��o9���  |}��1B;õFyU���vz����\I,����j�����V�lۂ4F	)V�����&J �{'��b�3�ɦ��.��|��$�-mZ@0������W{�vl��DcL������T�x&��62v}#�Y�����2�URm
�ؔԣ�2^ݙ_pj����ͯp%!VQ���8rbs��1�{Lڂ�Lm�+<0*��䉟V�Y=��#��$S��'�؄�����Kr��=	?��F����(l��]���ζ��2��FӾ�G�G��^�Ûج������r��=(|���=��Z�u�ä'^�{i�]�������7��Do�r�����üs ��6l#�@�\V�X�ݱV{�Ó���L޽��Y�G��k(F]�"~'*[�'	��1yQ�9t��1�М�a����ˈ&婗NeD`�wD�f� ��fB����7�W��I{�t��w��݋z�Z���5w@�}�#?S&F�k�:�&>�)"�펝��冗:�=���r�L)��h]��'�+��&"I�8�t���A��?���HqШ��C�M���󵠓�>H�.:�#n D�;�	񙠹��+�{�i��#�M�ۋ��M�˨a�s�%n���>`���*0�XͺqjYН���!S.J/3Y�)jQYv���)Q�t��˒��l�����=�O.[�R5�&nIl*��څ���fDq�5tנ��;uk8�k\2��4�!{4 �4�0!*;G���l+z�F���?i�Z���<��Gb-�]ō����[��B�$�3}ɰ����˛>�Ү�Mq�����l��n���ř�z�C�ߜ���� T���q�]��y�.
�/�Ra���RYj݊$\'A�y�)#W+{v��u��f���Rj[g�5�=���,�s�e��B����|2V~ w��0N�w�;�A��'�D�Ƥi,���ڳ�0n�E�f���c���
ՄA�p\&��j�/��Gzɂ��s�de�,<���h[�I�������:�c�$��� �Y���*���\�{�`x�o/�׏?T��
0�1p\��ؒ���i�����L�x��9DG����
)z�qB^��{��a��)~�ZS#�"�&���qG�ʞ���hv�Q4�5������g
�d7�S�o����#3�l��gF{��hw �O��~o�ל���������I�ZFFl��V��51ϩl�k�����̊�,ɭz�HP{�����xM�Mǉo����o>�&f