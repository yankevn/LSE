��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߎ[�zZ$D�H�=���3�r�-�7�Y��B
6����I?�����k�'aQ=$ X[Mo�o�����o~��P>��]p�]�9��D���M�y�~I�ʘA��l%�T=���溟q|��iN�NL��zH\M�I���u��L
�{��D 0�w��h�g�>%����2��*u��ПmX��)����/�̑蟕�H�����6[_ �oY&�,P~�
�c��~#�	�5���6VCA�F�_/�c�o�9JW�c#�Et&�.�Zv+^l��!����NB��>��92�L�'�/i��׿�ؼ`�n��H�L4K�oz�H��~�W�Hu�KN��;��E�	S/<}��x�
��^px]oaD�:.~��:��hQ�S�χ���Y�,���/�x��qy�yjZ�ڄ��<���'��X��
'������D	��d�b�l����K��!�uĽ�L$�e}O�z�!L�r�䌁�NB�7i$|5��b������*�]��@2��MPG"FA��Z��ƖJ��zoPw�*0.U3�k��^�4����T��%I]3�l��z9	%tm�����<S�$���从�<�}�9Ң�r�'����Jk���MN��}	B[:�b��d%!Q����3p��xD�!���zV�F�{p��s�niuψ��f��"��a��e|I����G�[}Aw���{y�H<��ͬ/�dg��y�����2ʠ�ޣ�?�]
e���̀ȴ�}���������kR�/Eb����ڂߟ�wm����ϱtx�)B#��Uş��ÌD�޿�<�$���
S~<�n�ZVؾ�F����Z�����m5�K.���w��.���9�ބl�8��+F��f��F���z�vW��T~����F��8�����.ˣ�4�0�Y���G���,^`?#�F.�2'��]vl�P���tn��3�#����i_����(�3bͳ��\�+K/��5�L�}����Gv/|h$�1�� �^�k�nq���h�-7TA����[����<k�ib8�KЬ�3�r��\5��.b�֯D7���͋3�n�/;�|:0�=�2![g;��tpOZK��=�vE������ъu�?ĤEhsC�p�z�܎�WS�n��̰߶����\8�CNg$޳�B��P�-�MT�V'�7�ےb�D������mU��0E��O� ��G��K�xe_
�u�BV�s�b5�+]̚C���-#��
a ��_$%H�
�{���V=Ƨ�=�M䙣���䆌D9�ʩՆ
�.)�w1"��zT �Ì����z"K.��
Tֵ��^IJ�\b9Y�n ;2�(\k6�I���~�H��Z5l���%)B������
cOo����hc�5��J�҈����X{��5;&�&݈i��S�K��p�>ސ�S�æ�ϵvzۗ��9Id���h�w�_�U$�W�y�Fg�ƺ��)�d�.@�P�r�W�у�KB]�/���x�����=k�ۛ�Lf�SY�XS�]���w���@d���>MBt����eM�s	ə ���y� #�l��1#�}z�'���G�_y�/XW���|�KQ���}�(��/]Cs�C<&6�g�@������cŖHbO���`M�u�L[�Yr�.�,J[1r;=r�^i\"+������%=3��ޱ�!�>J�ƻ;�x��𭘍6g���D�GQI�yI�Xjn����t��ߎ�Rwt�T�u.к���g���%�7(5�%�@�B�x�ߟ���X*No�3m譮so��N��	cF�\]5�� j��ǖ�F�Gm}|!���s��]e��ח;s�ӟ-�����0�L0N�n�a�g���j$(�1���`�c 2��� �B8��A{4��_�J�һpDӐ�=� ������I���]����SУ��IMzI�S8��'k��I7�<Dw#�v�|!�jy��j����asS4i�G���w�<P`Ȯg�|�<��(ӳ������I�R ~#�ZkH���Pr}�8�5И��d]�fP���ZG��~c�tQ�1����I���������j�J���$06��tH	zC�9[���]��+}Yr�~%��7�S�!�����M�1$x'�,Ym�\H�4ߗ��sz��Y�{�]
���5Z_�e��E<�=����z�gz��g������%��؟C��'Jf��ͻ�I�S:*����DK�����p8�p,�<�d5s���'Gˌ3����7^��DBыZ�6s_{F�&dvP;+	c�φ���`�k�Nt�H᳦
b���E��F�+����#�N����sx���6ם�	0!��uσ%o��R�b����C~ʐbS�~��\�R��$�+k8y�mw�8�|��.�ծq΁�W�z���8Q��?p�l.ì�a����ߺ�x���?ܔZ u}�����S��%Bp�Rt�aar#p�.��G�<a���Ay&.b�s"r��)��m-K��ܛۗ��4~�Z�#^�S�eM�ś����˪#���IYoB��1jF�O2D��i��6��$�i�FЂ���.�l؍���ϭK�ۋsGe���|Z�Ⱥ���?�:,�
��������������Or질���)��߼�j�x��ս�33@O�z�j��4)��:�ȓ�t߿����~�/��J׃[�S�i�0��IU������}/��{��D��%&��C`�*�c��.@��cUnK�j��:1�k�a>���~;� �l�"j�	��!W]%���WsQ�?
W;��Z �CgC�n��c��;#�r��4r���!� �	�C�qߨ*��V��W�[��O���W�sa,`��C��X������?�h1VB� ��T�ٛXU�;����SO�L[OX��x)y�г{�UO�*��:$
��ռ��*�ֽiXK ]��&8u����$� q��+�RLN���/`pa��np��Ȉ��?r�Y2�Yq��ՊaY�{�JY��!����i��/�?|��[p5+�M`�P��-�(� !��%�0@���u�.�m�0>M���:��|�j���_M{���e~����vIj���uGq��9|�A5�m7��6y����3��t��i��0;A^ޥy<�B)
�c�B|�Щ��-�i1�>�߭�j��"��}מ��R��u����d���pza�F,��a�͠(�F[�6,��5�h�$lvT��щ�]ө��WR/���'��F���V'�.��z��1,�-�䱜jf�����X����c���4J���@���ϻ��$��dd�ʂ�D����%���ȓW�W��ݷ��O��|Kc���u�-���r�[�d ��� Y[�ҝ	f ���p�"��ux�%�{I�;H,v�S�?t��8w�\�����f�޺������f� ��o����ؓ��.5���Nz�9�E�oh��W5s�"k��j��W�?�^��}84ź���n4�<��7�^v�C<�GV��?��<SL��#Ջ��#$���1Q̔���n]uy-#&@Z��P
Ң��䆬��ɬ��O~p�.���7ńF~I]��Y]?����)vW�΃G�v����Hł��[��w�̋k�1�7ɟqʴ�$i�!Z1��ќ	�c���f�X��X��2���"�~W9X�62%c� ��r}��ѱ!�ִ�a=���sK`5)��=��6�oB��k����Z��2�L�Xȡ���}��U_�nj�0�Ɇ�/�d���}�#�u�l���J"�kM1���x��M<�hh��:�$��S :���6���m�$O�ލ�6DT��TqW3���uA)y���"�Y&���;��_1,>q�l]\|��R�y.���`-r5d�m_��?���%�:�ʄ���Jx0��h��^|#�����6$��
�w�N�+c��ٔ�$���iG�^��q;��#_C�"/��;�c�<f��l���ҏ�u0�	��-���f2����u�o�F ?�9~��Xf�a�bU�'��E�%^i�$�K�؁�����u�bx���~a"����28d ��K]z�栭C9=�ߙ	��(�����f����b{G��x��#�����W� -n��	��-]�C�i�67E��/�J=1X�o�%�X %_��M{3ս5X��R��Y�z<����,�3P6[/)*l4��j;�t�\24��{_4��� Q}���>�����X-��ـ�4e�9b��[jg3\��{�
j��>4##]X�`��p��'�W8OV_��b8Z������e���Nae��Ju�)������b�F̊ ������c�*��5��%K�q����Y\'W	N�sL3>�ĝ�{(9k�ؿ厇������/M��΁ ���(��������j��%~ϸs;a���Zd���Ϸ�sX>.��6l�u5���i��0����7��� Ν5���g`@y��rZT������k��J����v��W)�˄��ܽ�G�&S���B�A� �;����/U������ ��P�y����B����Y�rL�{E�����u�p\R�V��T�a�@xnS*�{L�2ߒ��"G���(����v���'���${�����H}|ZC�XK��F�Cp.v���e�.w,��F����|5��N�Y3�&���gB�=B��C��ǂ���d�}?���A&G�\4)݄�(�uF��
a��p%��jl ��$:�����~�>��V�0�z��2k���? ��+�Ӓg��q�ɾz�(�ApCF���al�3��纈=�/U�0ҕ�ֈ�a���ٿ>V  OU��� �b�c%|�������G���y�1�n�D�I�� b����	�)c	B��,��eV�:���x�$5i/���?��+6/�ɇ̸-�#�x+蘩��,���0��Ҹ�`�m�4���T�@BC߻�F�uLP�	x���j����_��&�1И��<�VԈ���p�D�@���u3����`��@
m?�4�:�����G	ق[<n��Co��~�9HX��/�;���"��QRŢ �jP�:y� �X�ŕ2	e�_���0�x�4S!�C��Qz��pLa�����ۗt�s�������[�G�s3��@kJTE�v����&cjLQo�u�6/��w�G��y1:�WM��G�p<�׍�.���D��D�1׌<�(�|��T0�Z�&e�`pH���0Tz ɹF�s)�2ȅ���_�%����fm���8Bf� ����vE���*���J.�+$Y8	L�ukəPF�Q'���87�=�9��wPZ��C,K�2��b�Ƣ����n��뎅[�x������Jk�����"���9����tZ'F�ՊO�1F�G̓)>���A��Ґn�T��8��3�6ѫab}l�Lh0mW2"�
�sLC����ky�(<��2l$2���;��?��'��+}�K.1E&i�b��ĸ���Z��цâs������F�/�z&Վ���̡�U�f`K���Å�'��n-����X�I�ȇo�;w ��G~9���2�\q⒜�Ck=��(�j�����Kp_�х#ɕr�$�d�n����a�̥2��C&�b�VjaJ���\�?�&���F��9��Ck��?�xP�k��s�^�o����-���Dfճ�[�����e7�M'R�����m�Ȱھ/5-�,U`R�b{��-h��rþ�B�A?.i�[�����%ZM,%_*H��=nRZ�/P� >�~�0oh/����p:��.� ��-uplD�w�'h�	�3�	(F}�a��/�װ��{�x������7�6�[r�Q_2={v��$��>������2�zM���jj�=̓5��挦�<���������R�5I�+�|���t!�DfY:ّo��O)�d��ȳ$g��k��%�eu�m�4��8d��{w�X��E$�`yz�?s�����ė3 � �Dj�G������|�����/����k��0�,�͈�p�M��֔�xO+�Kv9#~l#A)�٘�@ٝtR]D���`
�E��J��0$��o��)��a]�c�tFF&�ް`�ڞI�ƅ/��R��r�N�l�v����ӱ�zw�j��Pr��� �D��7W�� n��rS[���4��:g玗����J���t��I�8yU��E����ܰ9�ZKk�6��'4�T��$���&���ح��Pr��{1��N�j�81'����q��(o�76<^G;4B���l���Ȃ*M�؎(;5më�T�\�_eړ�9̃�A�U
�V�� O;í����Cy� s�7�!�Si)r��?��� �OCmrLG���Y9�3li�g<2��[��1;j��ꁖ}J|p��*)Xh��P�؋�RcwM��3tA�����f�LlN��|W0,���ɡ(j{>�4��z�
�E����{0����/,� n��m�������/L�`/I?, �Ǌt��#��f+����c(�yf�;�߹6]�d�[LN����'m.�nK�qW�A�?|<Ƅů�u^��,��zUD�_��,���7ڷ�)a%n1�'���W�=T�RXP3f���w�U���Ztکȕ��z[H+� 7�E2Һ��*�����i��úi�8�ホ�)[�ET)����N�}�q�Q"�e��L�@	��*�i|�&m&[�b)���˫vL����
��pz����Q_�����<�{o/xg`Җs.�Y���s#_��餥k�y;!L8d��&?�=��V�.�ͱ�ֻ�>�4i!(�h�@��"�vv�<r=��6����}����X�!ǈ]��~�}���7\���cu�����tp�+�)���"����܏M��:��M}9�<��zE$n���T�^�r�+���>u�6��dل[C�6�#���H*�D�AE�R�n犑 �w��'}��:
ƭ�TW:HZ����j�h�Ќ�G�lugQh�!I P/��.z	�t�m� �@ǖ� � ����Oʒ������Q�'��V��Ѿe82/jx�����+>^`����M/T������1nlUTZC:Z%(:)g[̏p=N�2$uR�� �%rY%4xA3�:�9Wh6H2������+;_�
��1�_TՆ%�x62JN�EPB�%��TX�@�I\��F��Ȭ@���Ĩ�>
*:5mU �t� ��qVF �B�Ba�%#hU��p��Vޒ@��N�'l���K����K��P���l����G��G���MNn����$#N�G3H�ω�b�v@i��#Va�-����漤��ܫ�"ٖ�4j>z�l{���8��qn�x�.�B0�80F���g�!�U��z8��k��,IZ���/����z���}[n��S���;�"Y�T��8�%o��Ew̜x���Zy�jt�Y�z�@�\�7�]��ʕ�n���7�謁܁E�����b�6w�6�D���a�_�e��9���?1����%�;y&#�r$�lC*���j[�٭��t�a�-�,������y��A���QT��r���Yҕ�CUEV��`��s����a� ���f*=���K��ݚ!@�Fwz(�j��y�J�!� �wVwe�Rb ;>d��0V�r���?*x���.�E�B_L���l�*b�O�:���\��M��#v�U��V��|����_9��q�$K:���r��?���b���RZ�Z�S�wb����U}\����*��4d���xL[2�E'Og�!4$�@���i���{N&��5ȟ;��]=�?��%��j@�Poa^�lud�_Q E?��3��mf�v�o3���v~�Q�����%C��->���Z�M�`�����IZ�;G4�����awE�Fк4�s��M0%w�;�O^qe=��Ó69��w�x���&O��6Z�Q��6��Sɰ��+�Ԉ{������i,�S�ϯ��
tV7*�p4j�(���$ڵ	7�K�$��Q�}O��Y�Zr!y��UGaR�I����P�����W��;�ڦ�6��
�`�ji��Z`�_�'w|�����L�h4ډ��nj�YJ��̧�F'<D��>��%����t$i�w�B,)�"���7�Λ8����*�}_{D���<���{d�����)���7],6�u\ꢲ�����]l&��{LU��3���r�����B}���S���� Ti�O���U�CЄg]Ԏ8�Y%�����t ,���s '!v���/d�4O�O�N�=
��Bɥpͽ�!�^I�=������W-`�������R�M��E���-��oX�z	��eT��f�i{�	 w�:�A|�~[�%-�k�m�4��iX�W�����ڕ.7��թ���g�?6��4Wߩ K�B̰�����OC6��ϻ�.:kF��+�u1��iR���V���+�p�$+��ݤ�Nj1��Dw��RJx\�gaZ���5����O�]i=��� W�I� ��l�Zu5T��:lI �=�����6���E����搓�+�����#vVnv޼��ki���z�G`"���/?e˟��DM��v]�v( ������EEh��pN����j�Ъ`�x>a�V��m{�],���O��F{yA,���=�J4Nuh���Zd�N���Y?4=�+�)�����[7=��	IO;U��9���&v]��wZoO0-:j҆D��ϣ��L���߭,z-3�p���F�m3�]�Y�;%944ፏn�$�v0$~�v�A��9
�$,���.+��+�b{8zp�G�s'���V-�=m,]Jx�=0���	~f�O����q��	1��/��s,P�a=�E�z5�ɫ�'�4�AUyDU����1M��`9�H��J��&2&����L��o���bf���҈h<��T��2̰�S~��E�"�8���!�FK��=΀J��t�0݂�ff���`UW����_�Vu㱬��X��=��\�m��^�������&��5U �?}z��r�����v��ͫ�o�Ȕb�TQ��Y|i�{8L��-�K3�n�xL�q"�������-z�-|�)��`��w���<-҂��q~u^W��P���T����Q����W�,�+�sE��Oeat�N��+�;��۷�@� qeb3s\��E�����ZJ���]��E��TY�|�)v��a+=�7G�z�q�
f�6�q����ߙ���|;�ڥ��2pl���E�6�l��Ѽ{8�5�A5�/;y��u�f�.W���u����� ^ަ���$��0s��	���ˈ�Y�����PDo&�I-p��>���b�${\?�|�(`�K���>60�P��k�5�Ǧff���6��7�ǥ9��Vu~�_�/Du����KG���lb�B��ru�Д���:%��M��|$��*x����%B�}�P�缬#��$2]��e�S���LE��p$G$���]��<������ߘ��(��b8�lA�>���l�ۚ��2z�a4ŀ��(��;���t��
�,��uo/�n���B��k�ŘX-�[�h.�P^��q�H<k��5��_���h����q�+z|E��\X�Ø�[��ƕG�|���tqGs1jd�f��(�or�\�������op۱u�G%����8�Fwi�]�k�0v��r��A��_�wL9>�*{����`7�=`��b-h��L�a(��_p0�%��5�n�&j�J����?Z���R����Ջؽ�� ���F�{��wo�l�5�Nz�(�$�j�!�I1����E�5���S�H!մ����o��pGh�$&��B<�>�w�^����J��?���Dv��Zo8�.Y�������� ���}�pj��
���
���g�#�i�s���n]dm��y���Yj�ԉH+!�����XC��K_A��:6��ϛ"���0��.�U��0W�5�ޘ԰ڒ�4�V�Y��wB��^��gƏWp�wf`��9�vD�����8M���Z͈���������g3�\��w����ԧz5��$pl���ĉ���'�Ϩ�����P�l!g�zjCI�a���\O"u&o�ٮ�J��������V��[J���'������r6c�������aW��Y��L�c��h�"^x�Gj*l��^�P.������ڈ�c�?��x{x��u���OAs���<(��̨�(�x��ۀ�@��m�d��#{�R�̳���(�%M�
\���������}a&M�����d��Sy�F�D�z��.��Zd�"�(�+�F���$��$�!s�.k���'Ο�"�2`��k?�Q�2��9���=h�=��MC�
!����	2�y}Q}�Գ��c�
�֢��T��.���8R�R�kn�_C�>��$�2�،!م����F��'���_C��1�O��"�$;�����q��$4Ğ�/�7���s7�"4�^-�u� 	G��?y�]dfy���)b�K�,ePodOe�-���f�am�5�"�{��@u\��#��r~������.��M�Y�������=/p�i�>�����Q��kLRV��O\r��Am�ײ��s�s��n�@`&#'R�nϒ"9��K��d�r��ن��FV?(�M9G=�:�Y�05�#2������e@���5r�c�R�(i[�`}���/��D4����bl�GH�b��m�h��L]G���7$=�:1:Sr� z�nʽbswúm5mS�.٩wY����-��퍮������)�A�u4W�Z	>"����3���@�KBFD�*@�?n����3�t�;13�bH�{x[���4���������S�ä�.b��"~	�-U���{Y���`I0�*����������m7��J����"���@�)�I?>�9O@фdQ��Oy-�G��)�62Q~T 4
%�^��GM\i��s 2�<��u>0N��AjJ��B�@\�u5��򣸼�O�\v͖o��2�$x�(��_�%�xWBT�&�����'g�b�M�YA��vE��dj�
�_t}�@��U`j��\٦�s7�[pn�I��o��K�(L��͡*��Y��h�=�58³䕴�h	�i�S�H'���B��7 ��{����7�p�VU��KX�',�5e@K:iuF%� kU�,ً&�(�����m��P�K��C�a�$3���Ĩt�7~��%����F3,o�� ��+v����<�M�G�H{�{�ky:�OT  P��۲Fsۺ#�M��؊$���3�^s\��Eu'���b�TR�+����Gm�׫R�9ty� T�o�H��@	�Lǎ�?�MI1O|#V����9�4g%�� g�n�!4���N�N� %?4� T3�=�������