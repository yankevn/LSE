��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+��M�_<��g68�P����S��{?��
���T�B&���@{�=9�"�!��MK��f�7~���Gi�]ۡF�MJŋ�) ��"�W ��ys��=�1٢o��E.7���u2��+��J�Ҝ��%����mk��$���P�	3�#����y��c3��
�u|�M�����|�?
��-�=���7�Ȕ�ͧa���R�*�E<����Y^�&��`�ܐ*o+�k�2�b��t8�g�Hz���&lʙ��(�&˔#�i��͎I��'�P�ь�p8�PU.���+6�u"�c�OP_W8�Ʈ͂?����[d"�0_p�2s��
Ȱv-�Mk�q�y-�<Dm��_�[Փ���R�������_ǟ�U�ǘO��o��8��ؿԏ�+__���nOФ�����8p�S0�yJC�jq������I���r �47��]#�AQ=�M��E�q��l��`��C:�)��
W��!jrp)K6+5���B�7�I@� �K���v���I6�>�?wm^�H5a��Т��O]���Fm�s�Ҫ:�a�-�sd�a�o<��t�|{�8̣VlEn�	|i��-��9�*�	lg��(`�m��Ɛ�8��-j݁�ŪyK(��vQ*�
fI���5r!�V4�t�d�,VOXmFf���pm�~	�]#�x�V<��S�emj�������p��ݬ�Sz\�a,� �%��Ԍ!1X5���%幕�P�e6���AKy)p=
�u6�J ��,6��ۭ�*\�7�\��a�~�`��*���f�cN��4Q=���Ai�F��tct�b�wE�~ x�3�����^�#<�Hbk9Xj�:
P�UԂ�A��"w��,jXA�BІ6vPe~R�t�[\���pzo�Z3��5>	�Ӌ_��$�	6���|\@���C�fCˤ[6И���Ρ��E-v��^i?-����W�x5��Eꋁ���燷��Sc3ev����O3�1�M��u��2��{{��6�[S�j�GsXJ1��Ý���.J!hDJ�R����uH-�%���r_�0�ݷ/�6p3�kR)g�c����[:�:1?�{��*�i���D��,�Z����A,]Я-=�h΢a����W<?h�4#jT�nIs��,���ryl!���L�c\���������^r�'4��W�̧EC��}t�a�
�Y����\��x!6��uuַ2�t���"#�x7�@��ĺ��CBQ
���.�L�?g#[�D(9�`����%������,F���b�ݖR�y@������.�@«��xg�
�.>�ٽ�@z�xN��9����54�>����	ۼ��'յH���N:�����t�M��"-�� ��	�l���2�YM�N���(p��3�k����^0��31�@3~�Y��G!v\����e�FWV�_���c��ȏ��pŧд˔���/���^���Cq�K�y�U�v�fe�W�Yje�V�2-;B�h���ݛ���F�����"c��C�K�B�_��&���/�𿐀�l��w9%�I��{��H}�$ܹ���V���Kk�9���,�e��}؂�`+W(�*���+���P�I<���G���D��*��X)��8�?�6D��G$n1n	��J[(�e�G\Ɖ���Kd�
B���h�1�h�2�h�}V l��d���{^x�c̚�s�^㎼g�]��~�&"�dc��=S�҄=�v~8�ڴ-IF�L�M=~��v���B�D4<�|�mFF8r�r�P'�������)jp]��SR6��F�a����7�ه��N)0�3���I�<u�'<����E}��$���nMȕsj`����P�������!����
glG���l�X�q���S���)��Ӏ0/�
Ѷ�:��[���P=O���'L�;z�w�Iryk���f�9>�������9<���o��;\9���#�s��~�{q��"j@�r$�����F��`8�G2�OIbt���q�"$r��`U�7z']LI1;��Ax�"DW��E��~��{8y�UU7�Ã�"����*�/��씩[��/h��`<�U5�+��L}=[a�Ia��I��jy"'Jtaz|m�t�\��ӈ�{�R��~�"y����&�;���Eޗ�Hh�
-dhg��T8�L��wл8���`)C2�Xct�i.n�!�@5�p���P5@&?����Ds�������%���+�tگ���-+7��ȎV	�P�����K�!z�mevia��-/r�6=V�x���8\3�4���N)}M����ro�	�j�qs���B�v[Uaor��!r)���q����y�E ��g�z���4��[N���2{Go@=L������?������'��N����X��F����k0��Na^p|�Bѹ��o\
gX���u��?��;mجoZ@������H�����J�4G���}�8����Rм�Y1	�&�Z��&YWx�$�s���̏*��d�X�m	�4��R�F):��8��ÖyPZ�p�D���^�Arzi�Oe�q�4+r���@o� ]��e�K;]K���/��J_BTRN���x5����I�e�M�l��a�Ӧl����IM!�w���,F����2<����Op�q�`4��^�in�ک�����P�d�ٹ#��L>h�
Ս��"C�*�������x���p���2�=Z�m�'�]A����������H�q����Q<��W�j/��<��/��>���X��cLT�����Ր��"�*Z�~M�Q#�`��N�6�{��$�mf]�Lb��|Yi5�}��e`m�~�&�ϰ��k�O��������\)ʼ뷔�L2+�i�5�,Up��,W��-ţ4�tϹ�|1�hs����kϣ9��6u��ů�U��A߸�!����9_���f�#��ұ �����Q+#�R;�JZP�w	̈́�6�b@+��+�E`pq|�Z1���\l�������i�|Z�t�6&?
&@�����=�!b��t�iM2Ė����s���k
H�9@�����E�T3~����@%ŷ〜ޚ���*���iS
A_�ס�z�i�)ȡ?C��p@�^^gӝ�mXPPb1���-}�*n�12_>�h@���jaMU�J3; N6��w���MN�?�>>�����ЃW#��a��7k�J�4��:��Ɗ�$�M0�J�Ś��ɥ���@�~�gT|*n)T��3e�8f���\�WdvʤV�z��B Ť0�c�D����
鿥ft�GDT :���3��uu�cc�q��L\.\�x�VoՊT#$I�W/6��H�X�;�Ծ��ÕYI���9<D�h���.�A��2��@8a���	L�F3ʨ�Q06�	��ٿ�$Q��̨C�����ШB����^Iu��$�edI>�L=E8��z��G���}��Y��3Z�=�}R�	l��-��-��@��`�x���c�-n�G�E�*3��
|�K��� (*�z�VC�����pQ�Θ��M�Y��Ai��Q|�P�/mɟFBkF
�!B+�|�o#҈|���T��.��P�Y��tè�O/N�![@������Q�AC�#��c����+���2M�S�$*�C㴘�,�y9���PӪ���A�]4Z���&L8u�����k>{tw��+4����z� y����ͺ�l�n��أ��H��ԤW"9lh�O��2�\��L�啍�WVŒn�
oX���5��f��+�w�r��SLX��b�ьU��jE�ؙ��6qۖ`#!'/è0n��^1��J���P��Q@��9s�ٚv�In>$�痄+��	T���*Q�����u&xo�hI��-/����l�����n��k��W}lf�X������H$npC���