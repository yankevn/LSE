��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���{_H|7�chb��kS����L��ݲ���N�ƬK}�ڷ�!�rT��Y�������{L=���j��=��!���j���8L�h5+�}�=���jE����җ�&	c�ƴIlנ���Xh�b�bh0��w�.Ǆ��OG����1魙��
D�HA�SA[)v�����)�?�(BP桞�eI*g[Z��������7A��W*3�F�1ȧ��k��}��\��`�1{ ��@�W�9��/*7�s�[�BhՈ>�5�%�tx^� U�$zi�E0/:���#w�2��0V��^��"D#XN�U*L���t`W8R��y���qYE�6DB�A�8�=/�qw���A�Y���g�<2��x3hy�7_�?q��ĥ��2��6���R:s����U�wC}�!�%ϰ�3�������?�?UQ{ �i�n�x5'�>g��W��)ņ;3!j&�5֯.Z����w��wEŉjX^�υUSTB���n��H3�U��[gU���y4C�����꼸L�T��>踒] �ﶒ⩾S�`���0i�#�9�%�o���'J�B)z���|���=��y�+�ۍڌڰCx�@ ���!�OF`��|�1-����6�y2(�4p�դɾ�ʍ��������~�ڻml�6���#8	Ҿaʇ�_d��N�Ϡ�/�Ŵ�,�\y��$�"����R۶Gj�\}�gB���d��k�:#O��˨����=��D�ݺ]u�Z�r��j��xj6 �0��[���xDjd,ҷ�^�Q��0�jwX��] P^#;c��L�fk>�"�@�[�P�ӿ�d��K��޳J2,.�4`: )m����9%�f�d�2$*��N+zϹi1)���2	�K�c��d(�ɭu�������'���"�v�����Og�K��	����,t��c{B�)�%�Y�N&�*�W�e��0��#��O�6|�f4�xQւA ��=һ��H�v&���)����3����.�10:���+�pł��)���fb���ZPW|�`�z�J���yx�Nj�	5/n��v�^w�m��A������dH��g���=���o��Y�{2�,;��B���4�g,�'�g"ҘJ��晞҇&��z_�T��̈�h� M������B�h�ʖ��g!� �w��49�;�Qm%�)�=CXoG�Vq�jҜm���s'�-�O;@��}-�k�K^��M5��E��K���>bqJn�q����I�َ��<�A���$]<iib_9`.�s���X��ŭ�*P1���ݪ웍]�Ɋu�{�H/F��X�@������/�bfbX��`\i��5
�˨~H�s����Ϩ(5�H�g$�9\?��P���01�;�XBVy|p�&��w�hZ�h��*\�6>k-Tq����OD��V?C��	����~����[�GI0���F"X���]�\�g/���;s��EBϓl��w-��	?�ֽZqIo~
FΎ�I@4l�]DF{��#JR�)N��r�< ��aw�g��4�t�C�ޗrۍ[�$�����!G&'ضdXH��u��38�Y���Z���ӑ���5���sd�7�qdncD��Q�}�F��9�3����j"�VmJ�B�cQ�-G�ӏU��dP�V=�|�[��x���6�u�<����U�44:�3��sʝB���� �=R�R؜�3N)�^$�;���v.�[FQ!W�W��+�!E�_�H[��5��%�8��tH����Oέގ�@=`�*F�p��aA���'���ј������ϖ��	#��h���ʧ���_��R�ڬ
.�l�%`@�^����e�'p-�D2D���Tq�d� �?kM7���a/��fX]�]�*"��Yg�>��<�Y�-/w
P�4�8�?���nip��<����s�X$Y�h�""O�6��I��Mɜ��ݧ&R ��9��r*H��i$���2��9�4�i�s��t3*_}�;a���up��!c�-m:ȆN`kAqѨg6��W����� V;��6EU��w��ɱ��W�����k���}^�'��p��e�Z����M�?��舥Wk)cz�_9�dBgW��}~�`�ț������@�����Ry�йE�M�q[�;�=�ވC��YЊRv*�	�!�93���A��$��8��
����F>�S]��5���q2������[P��L��M�1�Q��)`��� �ٍ:Q~^Q��\�@��e�<m�c�#�]�l�����~I���H��Q:�ξ�CR�����k���H�u��e]U�/�jf�����N{�X��K�FfIR(I�_�~�����pC�1����K�$p��3�ݳa�α��;]ё6Kى�I��$˔r$��H�	��Eb+3���j�nO����K���m��D~�vR�^uX	�ͺJ�Y�f����$<%.D��q�8DE��miZȰ,R���v'.���-�͹<hDzV�S�-�/9 ��?�xh,���|s�p�b?ja7w&J� T"��m���ؖ.��~�tN2k���������c�X�B�y�{��q�@�;Q��P�@�����\[m'�|���������R�vko�A$O��/��|Y�7'M7&�q�#�*��q�;H/�}�Fhw@�,�).:޳*rq㗉X��ɣ�C���+�"6lR�h�}.� ��%�)7�$��y���0�VRIJ��������6���ج)���ڨ��cǠq"1~wT"6;�E=�U,
G�x!,4b�%rq�KY\��]�{|�t��P�		��̡���Q~co	}��G/���ո�n$�硒�F4��^������+C�}�%>$n�֍�$�:�8��VӋQa*���n<	7� `u[U��� 9�R��C/ah��f���Oɐɫ��%y�R�͖���*�z쁓�Sx�`ȎJ�h��q㋶u#�P��:�b�߲�K/畦J�\]`�N�4�I5�W7;�����w��H�۰p�g�"��	�O43�xI���82�3�̪w��v��r:�%�+Q�������<�{*Znc�t|<7�̿��.��	�1����ݶ����GO&����;��i�t�'��(+Eb��cK_���q��A$�Ŏv���i곹���PEb�B񊀀6B9c�vP�
� �����fo�%�5Nm� ��q����!�=�$'r���Z\h��]!w(!�J������';�h�-�p$��L�:�� ��%�����1Tn<~KM��!\�D��(?�:��g�8�@@XD��{;��o�m;$�=R�U���=����������o&�վHUd~t��m�]4=�CLd���7-�Z��"�Rʂ>��O�r+�Mu_������]Z���"�!�"e1;��9������t�p��dE��C�0�Tz���H���^��ˇE�
�$��p�:2���#���x�2��<e�j��R�zm��~g�)��������[Z��5��HCV��D7?KcUxm�N�gJ���{?#_��Cc��TUD����w������o��
�ym���vg�:
Ǐ�j$����S��pg1)�5B����?�3�|��iSc��UA��8���@���'#��ȳWx�e�Jv�s	�ٌ�����s]X�;�TH��[c>E5��j�����Q�a��w�evې�#A8���w9g�p�5�t/�����q�v��u����SI���W^a�
D˾��w�3�Zg'�S5)Z�o�u����δ��"�0�Y����x�^�������4�+�w����E����*In|��J���|�iH�����px`,Q���:��b�Р�>N%��(-ciާ7�������`&��[��\�~]ty����T��I��0�ĵ��"�
�.\���,9D7.���i]����`�Cz<��.X�x2
��,�:f�$�(�ɋ�?���B؞I�gå1�l�=PG�{� �h���q����<�߁�8�(&����U�/P"Ok���I�d�A?x9sO\��E�^������BJ�i�t��ź--X6�>n�ލ�p�`\����B9���h|M��]�Gj ՚�W���U����=��9x���!�ܡ�
�*J-�ᾭ/�c�we'�v�3Q��n��`�q�����Z�B�ΤQ�r��/e��g��Ej�[\��^�S�;3H�;�K�:lת�Q0|)Ij5C����}�Qh^ֶ[y-l��Z�D����BJ�e	��Z(��V�����lY�𾨲�vKU��l�oU�$�E'�=�-V��+e��ʛ� %/yn�9&�'��sY��؇��*�z�v�XaH��s��<-�X�"�	������Q��g!Q�JBb4�B�gX_߸"e��?27�������r"uY����Y��=��t�f,�D]�C�-��I�.'~��Ȃ�^���!��ʋɡ�vߚ�+Um�tԘq�3��6��[8���Mî#���#���%s�I�$G��Ĝ��;]�תx�7NF/즅0�zt�b���'�a ]��A\��ps�i��2֎?pCI�Q�W��}R(.4���ƍ@N���Yw�Z��r�����<0X,��S�3+���lإ�I��u�@����=�'ތ����`�*�P��r��q�vCe��	O�NK?�W܌�j50%<�|P�NP�!�Y�OՇ�n3�u�A�ِ)=&��%m�c��)�����Be�)����"�g3�*Ά��A@x�f�}��?u�W�Z�AM�vM̰���}�bEgg����滏�,f�t��Z��Q:�(N�(��&GR+qf���q�o��?��������W����|=��,�	Y���9���%��!��e[aZ���yM�!Jb�?�P�C؈@���$ɐ���n��e,N��{9�!"%wf͸4��Jey̸�ʌ��2���k��S
Ĭxx��)���l{�q}�;=;ٺE��p�f{%�?��*.g�-b2��W���D-��'[Z�D����]4#���n��ts�L�N@��a/C�8~�B���G���M�_�jt�!��d�8u#�=(�ZD�J�=!u<Nⰽh}A -��">ׂ��r��\�����C��I=D�y�}�:_�����oY%T{/�#����wG&ݙO�O��4MU���߇�6��b��?�[#��q�K��$_N���;b��i���� �r��z7�&�i��d��Xg�]��\`q|aJ���Xq��8��*^ /)�ld��\I9k|a�48�����]`q���~�o&쳕�N�L)o2X�/1��܉��Z��p	N]�xm�H�(��@3�*�'(�l<�i�t ,������P �.mbc�C��-x�*�,�� ՘	I�o@rH��t�((x�p�)�a�\R������}\�n�����E?E��wqh��Õ��PP}�i��d$��[Q���E��<�u�]�`jM)Q1�p�KR��,)�K$bGFC�@���̾���4gx����"�{��e��1���j�1i����>��`&d�Ҏ�v˲m�
<H��A�><u��&a�y+�Ou�Ʈ��7����tL�i�9 x30�J9M4�����
��%3.���K�#����!��6�}C\2�rƮ��!�[:��yB ��|�����I*�gW^쥚��s\M<�;��U@�@"ok��<�~{��\�5��T��a�N,�ԙ�	�N��Nc�4KAB��&����fvP��ݎ�6wXG�@Eۈ+O�-���a�Sa��g[Ҙ�5>�2Lvʛ�H��ui���pd!0I2��^�����suĎpM-�<�Q9�/�e�52����Q
��̷�o�V-��
�F�X5�����-������eq穫�>��׷�Y��(W���YF�Wz�B�4Ԡw����sE&�b�3}z�Y�O��*L�Za$ǗN3�ގ���P���Φ�ja�1��*~#�9��B������
�U�ń;mF#���g�dN��ף�i��<@2�f7�R�쫦�:�ޟ;�6vY��f��$��5�D��r�(��dU���Q_�m9;�b���4ԯ�1�V�E�˩��OX�����%��}�X��<��G/��h�t}늬tA5_�3=�>Q���T
��b�rY vY�Ņ��j!va�.y�/q6�ֹD�{$�v?Yjڈ¤�"kO^n-T��\�F�k'7��<�T`�n�<W���i:���
h�=s��]�d�������=�{�:��ޤ�7�I�t\3�$~��)�#Y���|�xs�z�E�;nœL:��pa�+��,k�&ʴB��J�yx�֛l�P'��.|9�v� l<PӠ.�l�Aة.��'��� �tV�_� ���У̝gö�1<E��%ԃ�΀j���kO!_-�'��D��x�����Ұ��n���B�٣x_�u���Y��ܧf����ԇ�P>��sr��֢1��>�����bv��9pAQ��J�]yI�R����V����c����Al;	4+�����U!�][�0W�A�IF��ܔ[�Qk���?��U���=U=�ƫ<`r(L���(���Y�,#oG�㶁E�Bd0�Y�Z�����������,���\�S���x����j��߹��]7ّ(=�e�Vg烱���J YU��*①n���8�wlWj��QP�&�D���2�2j�S��}ⴇ��j�K�*�S����W�i�0��*��p�&o�ëF�<;e=��?Í��I::���2�h�X�+*|��x�Y`���&B?�f���aj���	2a�!���j7��1�b��$INS�q�Ka��a��<���Gkw�hBsI��R_�e������ �g���"ˍ���D]\�}���?�_*�6^�@�Z�3��"� ײ�f�C4��д�B��[	�xQU�t�Kl�p��s�+b�[�nŁ?9	�a����_��������3d�A� U������'�#I�M�^���u?NZ�?�h���L4�-3�s`�X)��%������j=`�2Ƹ�M�_�I����s�:��k�w[���b�dnf+.�,����ҊsC�9(K~Ks=>f!�;q�]nl�����<��ݣ'���H?>u�	�`2즵.�SR���H@���s��6��
�@O����b�������:p�*~|��M�����T��q��A$䳇@��WX�iҼ*��6'���a�(n�s�Cܮڲ�u���uUVL���˹~�*S�q?���2ÿ���)�"C'ۦ-�6�Ph�N�ٗ�%e)e���(>�ۡy�	�q�%rl�|k;�+�!��TJ5A�оئ�m�6�Y�5_�l�S��Uc>8�d�������6&bS��oQ��W����Ȥ}���lA�i�bxnŻVIŜ�1F�`Qk�Ds�y����EH�a��T����~��9�A�|2я9�6�bq`E�+�AW�^j����C���	��i�̽f3����+,�$S�;�c����XQuw�ŊA��Ƕޓ�&�ݰż��<f�S�O��[�TU���/�~�<Gf�\�EH�5��/�B�zC(��Σ���C����EN�A���O6�,���+Z%h��;��q7��I���|6N�Ma&�z�F���h5�+�	4U<��nqt��{oŐ���.�N���[o�0��g}�H��T ��|K5�	�HU�Gj�\V�h}���v�����+��H�����I�>��
���dL�O��ҟ�� �Zq!� _Tղ��3˷-��Z�P�N�*Q�ͩo��>��4xRe��̳ d��m|ɲ��KȣŚ��0JĿ*>�$8AQ�=Y�c�{�ڷQ�+zK*��/�F�?\#���D��K���\�**g�Y7 ����1�����~ �o-��͓r��JK ��J�]r�W���,�z�I%�#�w��=�H�4�����;�h�����L�YKPu�-�	��fw�C�9�N��qk;���xh�#���ԝ��{z����5�,`i�����իY���q��f�A?hq�ȕ��ރ�D?m o�y�C���ɖ��u�f�����Q,|5y�_��jX�6�2{~�1����0�;����O�~�toql
1�p���(̲+5���"�i}�A�7����+�N2��$�9���Vx�S�k�f�S;68�B9�;P�u4��E���^��I���U�h�X
mͽ�&�ܢ�M-�3ӹ g�te(4� f�E� Z!���2;���`s)�8�W���4�N�\��������V>_��
Y�M����aL�D��9m���н�L�y�h��O�l�m}ԋ�x��xe�Q�<�:�����%�IȘZZ����9]g�H�`�Ea:���(c/�&��|!�?4�J	38#>�[�s~i�w��h.����42c�*�T�6	+s_��}���Q"���6(B�Ju+g�� �i��io�2n�n�X�nN��7]0�~ ��8G�=�t5qfr�D��u��Ԧ���C���
���rS���y�>�DJ�i�F�<����ΐk��p@�nϣ����p��~4P���~<�hц�|�J�ДW�2�n��Z�R�ށ�C���8�?#��z4����Sׂ��a-_����A\���>(=�tSsdw-�S�/~�R����i����@�Ӽt�U�N��*�;6ȶ����{�2>���?�w�O�ѹa�ުw�������6��PL�P�cO�K����[G�4χL<�:�<��+��<��#�5LgT�o6��fW-�᩿�5� Y�Y$��\n�:@�����lp�� �p�Q��@_�\��b�xX��92_7�k.�ߊ>p�P�������Rج��e|��#;��2��l�ݨ#��9m,�P�Q�g�>� ��N�KK)2���ΤA���L:�&w�<��!9������2c.����"�o�R�z�U]�����BPaϡ����u5,C�5ª�%�����}�<��P�Tqzx�$����,�r��}®A9�����.�����˶��R �Q�s��5 ���^���B߳X�&f���<�(+��e@��Z�0E�
���\"{�t������y���5jܹ�f��lt��wI�����K���7FȾ�S�e��in}�n~~ ��؊)<��2�s��{o���obv=�Bv��,5��#1@.	�7��d��x���(��s�2)۸LQH�td"���;TG�d��ɷ�Y�턾?/�P�X6���d�"�Qi�|�vT3Jµxx�:)z�֝gT�Ǌ9���I�A���˙h��t�?�h��~�H��#�r��Rw�3�� �]�{�%�5�Q3t-v��.m�u���OY8L<h+� >0L��˿��I��vtNÞ��n��C������Ht.��B�u�և�зXŽW�xv�G�&�)�u8��5�"g��7�`�X��MY��n�y^���(���QG.����Ȉ�EI����c���U��p�v�Ә"_0�����^a�zy�L%.�:�V����1$��9a#?���<��P<���h��q���������L	j�?z��$E6+���C�G�+L��Z_��,��%�-e讈X����E0�?��LP���h�\V��L�at�*����N�<p#C��̒@? ���+EG#vرd����J�5m��n��BYU|�f��;��t�$+�1�o�c�[���-����k����V�⿰)��'�6��ב��}a�Cs/i�?OhDW�f+Z���5k�=D�Dt�W<���?
H�׿�S�
��;�`U�ǝ�ĺ�?+�k\�}�x�;ZV�\ۜ6�̓������@g����$�m_�p�����y ҅���5���Q�;�qʗ��M?��x���-���9��k�e��Wy�i_?|���Ճv�6� vyc�~v�؍Hd�?Ҷ����>����1����"�yJ���#/Ę�	�d+�)̠o0�7�e���Sh�Q(aG� �*��e~�6w� �,�+�L�B(��������D|&
���h�c��a$� ��^�;��{� �_�;�.�C���� Ԑw;�[Y�Y?�9�
��&��c*N�O�w�t����C�^����A����̌���Ѐ��=
[���Lƺ�*u�����E8D�BA�[����	��L(��ܦzHI��j�w[�$�W��u��ݝ~��3���K_��	��`s�$N�;ď�}cT�����&�C�Gh�����EBׇ�k�A:Xz4A]��+fN-��^�^�,4O=�ڴ����zC���8!�A^h��@���q�v�˟ԋ���V
E�=g�YZ��$|b�f��[�O���"*���e_A+����PqM��G�N��\�a|M�)d����"�mN�2l�����gyfv��em��;���f #�4}��SL�v�����W���U����0���{1�~I�ƣ�Ȣ��8����+�����Ñ+�����3d��w���}��zo� ���qV�~Lr������8�QΔh�ê;��&}TE#m�R�7\�a%��_�e�T�!%=z�jr+�L����<���k�Կ��J�)"vs�c}��5$��\�$�ïA�o�1��R4�%\���$�<��edG�*��l�������N���0���R�3���8���_S��o�����ƗY���J>`"ѥMJ%Bz�^�Y���ϱ�݌-B�>fp�jF\2� �[�8iV�8�a$���3�tcO(;M�S���ҮQ�,%�z���fw�9����l��-@���x��=���D���4���)�z��r�V �5�+0
������6d�i�ߌζ�E*XM[dKS�(�?���ҽ��������=[�nܠ��&���߼�O�4{f~�	�Z���77��9q��ל��P���=27R�B@r�uC'�ŷv,W���S�a�f0���vSڲ�i8����2����E��Oł=���hy�F%%����/�JuPC�`Fr-���9H�%�30��m�M�x8�J�/U���>,�c_JZm5|�ȆؚC�M��z�����p��(�@`�����	�d� �K(Ѻ�`�&t��?�
Ur� FCY6C`�6��qF�*5��jؾ�7�"���nt�Y�O����Rյ�ѱ���<o��z���C��9�s�I>��E�v"1�ڮ� h�9-��7�y�ȁ
ɷ�]='}�H�>MG�jynpf��{��iP3��j��aq�V�7]�	���/�n	���X�/�ȫ�R�]4�n;�w�R�!v�;�XO��܁6�,��
ɡ, 9qCP��=l,�*�[����}�w{r�G���N�uc`o�+%�yS@��I��6��ԭw��~,0s�4��n�}�?5�e1���l������A��Qu��b�9���w���m7N�Y�wPLc✯x���)���u#{����@!L�g��wR��~ۻ�R�� =՞ 7�@=���f����J�e�!�^��w|]��3��o3�.�ި����t�3��Q��n\;u|�8�=�3a[���.:�R��UU���u2����q���q�?*�v�J��9��+��������g���0�!�|��c��׼��?��Y�؁����T�r/�Ρ���w���YX|6oo��]��.�c�m��#*o��N�
�ێ��e��8�n��0\�pn�iN{��%��9��������#}d������޿����9;�x8�d�: �IF|���y�n�@Q�j��ã��"���>�e#,�f��g%�q�g�E�W�.�6!̯	v�4!@?��u־� �B��~[3�kd���s�|;��&_���a���D4���3����;�6=^����d������":�I��٨�`�»�:�c)���= ߖ�ڙX�b�Ԉ��1
u
��Q�E9��?��P6�pG��J�f���J�RoJ��b%i!I���d4�m�<�	\�u��z��r��J4#bAB�/�;m��J��c�0q�י��3��(NJ��b�Yx�@�<7:�4tf�t�l�oP��e�ϥK�V��)2�<����;c��A���x�Ė�������YH[tM{���ta�[��iZA��qd������B��۠=�1�&)�] �W��rH���A�y����vZ�3eN�M��L���ϱ�r�\g�͟���!;��o���~7/�=o33���f!����ޡ�����}h�O�v�į:l�ዖ&�&�Qyak�#Ea�eҷd��z����lJ�����a5j+\�$�S�����|�����f���)����B�D�DjDɒ���>�����,Սd���n̦_/z�G
��z��\?Ref��(] �]���1�(0�\� aY�{uaE6���g��?�UdP��C|�Asv��ȩ����n��Uq��ж�7\4V��m�X`�@�݁s(]+���2��s�hN�ͅ~i��� O\���I���d�n�
�&����ʷ<i}8חH��m���O�#��gݷ1��f�����W����$�m�gq"	VZ%g����-�)
��}��uX��Y��z�,(���S��ipt����@A�4�uY[X�/�f�w*@�
6]�@�
�-��d\ۡ{���M=l��~VL,�r�����/�,�L"�����`�O��~�ݣ͌o���͉�f�̞
g���4�I
=C���r�b��`	_N-��]o�%�0�� d;ȚU�i�qw��"Ӭ��~,i��w�Č���C#}]يh����U>�ˆ��I銑v���ǱZ{쒙fϳ=*E�/�)"Y�g,�Mb�dqZ�J�t���e��:�~Ɏ�źN����tdE�p<�tQ�l��F\:�x��ba)�x!]OP5�k��Q⫐��/'R=��B�Lq��J��Ūs�2]±@�&��pۋ�Ts�:����)!��%��[[��q�V�!O#DȌ���]�)S�y�9�kײ��Y�+�"^^	U1�G��J���$�[��l>A��5c-/Y��VY��vh�p^q�7�M]]��?�.��ĥ*Gp
��z:�=y=`�@;�����+>ĈL��9yƕ�e��F����Z`[o6���
b>����z�_l�� ��;G�����	h)��,�m&9i��J�!�:�	7�4��j��5��TG�!fz�0������i�} �[�k �l��D<*��8�� a�h��,�)-3C&�0{Z!���m�ĭG� �g���zFP?��H}J�tT#���@1��o�M��q����ՇY�u�Q��5��n�:^�*��Q�N�b��3�i7�0���_���GO��^�0h�	S���_�;����h%�q��Ef�Ή��BKI�9�?d}��\|���ФF���k8u����mFS��F"�	�?�rg�E+sߢeS�Q�1k��xW����*ez�����;+W�w�O7P��VgE�S�Rh�E����Τ�7�ƚ�����Ƅ�Cz��k�Lű6�M'P�;����6��6o��5�CnH���A`\����P�N���S�ʰ���X�4G_�N�=��̻u9�ػ~;���Y��.._��V��)��Fq�.(�Q��~����i;�A��ǝ��m�lqZp#���ڻ���8̱�� \:1����Z�g2����b��#�h{|�UQ"�LcQ#������Ӆ�'����\�[�j/�ZTLEJϲ��(��vck`�Q�J&<�PD^��HDy�-%}����=RV�]��o؅oz�\T��E�7ǳ�<��3y�ݢUq��d���g�q���	=�D��hF'�<��/C���]ě�z�}���=?;�bpy�g�G( 	���	�~�i��_|U�=?>q?�:]�l/��]e�r6m5&}�/�k�TI���ӿ�h�z!�'H�dPt�5ɓǰ/d�.�a[�27��������tR�+�U?*'��w�?a�E݊��BV�����J�Ky��+���:mW_mY�. mb.e���D��>��ͨ>#;�#*]!ډr�
��f�q�/��ZXcC�C��D5D��C��A�g���Ǵv��ʑ�^S٩�So`�8���,�:��"(��e��\��Z���,�o�?V��F�n�{��E~H�������_Z�_T\ء�P�N#C�����R/�7��i�ю[�,��[�D��\���*r�u�f���%D�LL��aVD��:^�a/+��#����F�y(n*�d$�QG鷫z����PK�'�S�a�/�(��y������]�f��j�tTB�~O�f`A�+d��/�@3�]�H���Ʌ�������ѿ����h#�u@N�����^_�=	�\��g���e���u7
�۬߆�aQ8Kl^��&�\��F6?������{�Z+,k�����k��I&�1H�d4�E�:�B/n�9h؀�dx6���,4�MJ��b��;bx�.u��i;1����(t��?�ǾLJ]�~@ET����B]s�g��Dc���/�yW�;3FU�.����+�D �<��E��/r;@��	E6��4�$[:7�������A\嚌D"�F�w|�� ў�C�m�@MST�A�xl�eۑ�����O��~!.5Q�s��剨i�y*.��ݳ7����q���ؔ��8+W�����5@Λ���s�!R80�{���6�_t�]�b�UL�5Y�%/)
�) C�%��v�3�"axUe+y���ԩ�[�E�����ƭ��*פ
y�׬���DMd�/�r�_6�D�V]ڿ��!�8͔�:��t/�i	,@�_`�$�6��������->�oQ���C�5ۡ�o)Q���U�0�MW(����f�v�aR��aP���=c*Q��>��.ܚ��4_(�*��߮S������^j�����v��f��sٖZ`��V��_ݚ�y�"�2��]�_�l���� Eo�К-�!(�:��:�����w/��gH���ĵ⮩� U��j��&�N
�Ru�֯������3l@@�C��C�j��r��/�@�#�TN_.0��7��Lk�B�(�:��1��ܴ��˂��s|�r��hW�t{(����_��G�oܖ�Դ��a�}n�B#�x����-b�!�؂����W摣q���!��M&W�&BC*Q{S���)��-�a��s�/�����4�2Yk�6N����`/�D��[z��*�������-�H7!2��_�V�6J���Ɩ�w��F\����~�(���耐��ȑk�{V�G+���:��p<�ʥ�dI���K_
��+-+�/W��f9T��"b��cw��8���j��i��	G7�����%�0�$��{�w�>�}�ȓ��Jۙ���t��7�\��Z��@��]֋)�����~��-�yI����bx����
]t�]�O
�!�ua��ui:}x�4�n/y���D�$!
0[q�#3^��B�;�}!�P�h..�fq�g�1��JaJ��e��1�=�_c�&���qž�Qm5 �D��뒫Sl',�C���eƪЄ��7���|m��K-����p�J��7$=#�3�%�+a%u �T��f
Y�qMu�i5�����{x��g��쵇��?
qC�B�����0v�������)��`׆+�Տ��[$X���9�1�JVqI�j�oy�K�䍄fvc8-r���҅'��1��F�ኴR��[к{l�O�%U�KD'�2��Au�>r6�o�EBh�Ϙ-ݏ����V�:%|f��?�����˘
���~D�k�)�h=�NB��j �Ǥ����s���@67C��%PL��i���8qQ��5�Xds3HE!v���{ʲ	pU�8ȸƖB"�"$(���z����h�`��(�'��֠�}�pIz�Ȟ��M2�G�jr��А�杻߃��ͧ*�}�	�0�C���
)���B��L�*Qca��X��t ��Z�u��N���vB�Қ�������������jG�|6����'~+�״憂AX���Q�O��+� �\����}kF��M̱��l/&ѓJ��Cv4�Պz�f 1h/J��P�lꅪ��9"�F���a�"$�gr����֓�%{���U���A	KO�o!�y��C��O�-�Q)�Z��)8ԝ��T�L�{�~`��u�����ߜ�"�3 ;J~�h�GÀm���J�jW�6��ð�k�@�x��;0�`�]w�ciĄ����W�q��g�j�s�C�8��=�!��[sa���T��lW;1�<�7MS��ޙ��?�*9����Ϸ��w��kJ]nn ��JT��o�Q��W�<����޸�]�q���	���0�#�2�W�3j�3��~�f=�N�^�����Hw�g�*g^h�8����\��{�=x,�$�9� 'd}�M�g��5ZR(���l��.�m���A�`���Wa{ a�����]��'8�u�R7�i!C�2���3t���
ōY��zUc+����#���A� D�Ze��ģȍ���n��E��������)���ʛ� ��.�|a�V��)��X3u7]D;��)6G�%Kܡ_gz��̒��P=���V�<]��b�Q�D��J�O.��!_�b'G=i̘1��p��k3|a��ˈl�5:re��6����҉�[���|��N�B��#A�l�!D���e`�,?�ͱ2��6
�%���XN��{P��W�-��}�9����s:��b9_�5v�o�:$��m1�M�xP�E�9���b$ʺ&fOz_�v�&5�_E.�4Ԃx��S5�$?(u)���י�g{x#N���6���|h�wP$�BK%G9>����O!Qm���E�5��/�l����}3lL� �'���0>i4ʩ&���5���tmTt����]�����O	�T������F�MH{��(+�-�>W���t�x=-�/�>SÜ�D��&�՘Ӽ�2��Zl��܍5��m���u��#�j�z��.�����7&��<�Q-�ys?^�2]͔zPGv��ײӴ�Bn2�l��h�ZH��e �X��wl@�O v$u5�ϙ�4h|����@3��;\�R����FyY�c �H����>!ܑ@�K�}��L%�Y��U3*��_k��8�e���зgW	�;+���)P�Pl�	��_�<�ZnR��.���ecg�x��kՕ�����]&�iT֭X��V莏n�4m���SB"-���8���q����p��S�ŔC &Fy�B���H�6�}V)+�g �T)^������j�0�5y�X�k���6�����5^� /��"t��g<�
+G;��u��8��_��Um��e�;�Q��2����#����@uc���)��u�_��s�g���1����
�%�Q
-?�[^'�s�<��e&����]���|��Jy��H2�8-��|���Q>�OV�|;rk��J=��"����g@�,6���ԡ�'�64'P����Z���:Ǜ�t��d�T1DF0������s8�Ta�XB�鸺�a� vAB��}:�>�9		nh�ko����&�����&'1�Š���O��f@G��o��|�r�����\r'�g��)W=Ta�U�Cu�H�Y���@��^����+��"Tg��������yR��0�s��)���eR}p�(O~@:��8�Q�Ws-ud-Ć�B������֣Ř¢ӏ��dO_$���l�B2p�P'P�O�	�:�3cx�?n��Њ�t��n.�������`xI@]��wl!���W-dDCP:���÷g?5���?C�7���V�5U�׏�/��?f���N�,����hzo�+���U� K�g�k��&�A�1	�BS����N���J�g3�F���l�A��.X�/����$3�CW��R���*�M����*#L\�Rwv�( �BEw
��#�H����&��kh(.��/n��m��!�*��T �XM���"c�H+�mp�Ι)����\��-O��`�|����o� p8�NA�9F&߸�m:!!N�@s�}��b�:w��B�O�N_!�t�5��׆��sǌ�����h?���z���{KP��{�)��x������/�c��ƅ��!��ʠ(m!%��|�3�K���F��v����U�ҏ�����{q?��{��1Q�Y��l7�9�*�̰폶(�h*g�]�#����؄�_M�`�t���*F0����d6�#�Z��s����*��<KT�7��a{8�� ��)�4����b�C�H��_
����M���1�j��}�:"P��7{�ш��P������2�c����w��af����P�L_������<���3��Q�{+�!���Z�6t�(/7訪���|3G��ݱg�� � cNf��L�����u �J�.�������?���a�G����!��L�8TlC����-�3��
�_�UQՍ�%w�/����*�R��2��f�z��{FDK)��w=|}���e�g���m	<HvEa�c��c����b�_L?��聁4��3+J�]���4T�|p?�̟^��b�mT�n�/)s�f�;���mM���Ψ[��i��D?LH�����	o/+4���c�j�=��2F"L�\��pq�0O��q	���Ɛ�E����	���A|䣪F�e;-�24|a~"N�y8� 6���'9���V���#��T��a�h�.C��BC�x|(H`��'��b���4Zx�Y���@x,,1���~��f���|f����E?�?��ƽ��l���P'�_Ɛ�W�&=�fc�� Gj�?��BJl�h���k�(���A���ΣåuY� 6V�_M�
�9����[GU�s���*���=3()�˙�bv��6���z�C�L�֛!�m�h;��w�_�%�u���Ֆa�$j8��ܲj�N\3X&@I����G5��=��k�~���,K?P ��q�"��	+U-x!�ډ;`��gR����aR(��G�5��Jp	0�j�����ՔJMď|6!\��?hG�8���⚝jU�=ᚏx��1�֠�Gϯ=��`�tɒ�Ĕ"O�Y`�&j��e属[��F�zh����X� ?2|ŉRe-�,i�Y�a{2�XRQ����h_�9zN���-��1��2�3�GHE�R�ϒ����^~����IG2��]�BL�ӯ����Z*�V�����hǬC��PG9�؂w�ƒ?~U�Q?]ć�_ŋ"e�%
���Վ�=_L)�svi�Y����v��:���}����?�/i 2�$]\�E�d�����W�g��Mz��z��/	�Lo��a�:x�D�TO8�z|��
@Z��k�i7�]��)��t|���(Z=��xfi���%Y����)�eU҅����TɈ�������^/S&������ LZ���[/ni���7�j� ��ŸB��B(b�=�!�=VU3�	(��V�x��}����i���f����K��&�L�M:��K��}�|��l����O&��fb��������ɟ�n�ڰ��W��f���yh:� 0���l���%�&���"v˚�C .�͛�L��T�N�A�#輡�vFG�eP����Oc��=W�O�\"��wHå��v�I���f́lA:�ۀc��͍F���u�ˢvC�in�EM!��B g�S��t��|�fU���Ѧr�I���I�"o��>!1ʎ��`0�z$��d�M ;��!+͗	����]��5jG�E�jR����&6G>
���]��"'�ҫѴ��Z�.�W�1�JQ͵UqQ��ƛ�s���,Q�"�����G�|k!htW�'4�LK�b��\퀐��33�<IDcJ���8�p0yv��Y�����x'�f`I�"�+�4�Qr�7��y}_�mC��|D��aN9��F�qQ4m���tǗ��#�9�ّo������Z�'�?6��W֍�ؔ���"s�ׇx�e�Sr��,�0	�~�ce;�~�D4q��_hm�朓5�:�7�?�2�ci+��LO`C�̒��S?g,�uӄ�c��¶�i`PR1�ޣɀ�6�4'6$��?����dS���m�J{�5
.l���s�[���暇�Y�{2�|^��D��Ц��>}�U��M��)�/�l@�>�芐k�c���\��&j�;��uo�ЕDy@�J��"�EF�C>L�<��u����Һ�6Sq��v��r����R�g8?Z�������A���.�����ä���g�\�l.�Zpb@�M7����-�ޫLDqi^�$���&u5[�b0
�����%�Ɯ��+캆뿦�6���-� mOƅ+��@���w�ݷ�H�fS��2]����2ŕ���U+:�o@ x)��+�׈��.Y�fd���V��!�-Ã�5�4�x�/��/6���z^�G��{�J���u��r�|6�9á?��+��nƂ�i-]���ք�r;����|=i)����	�'����y#�뎔[�W|$lDaF�: ������V
8��X�.����襂�Ѵ�q�4�4l�`2�DA��)j0�Y$��ic���\��I1�m}M8�"����ؠ�	��L�1���T�m����Th"�ѕc�,�&����^��<Ƶڊ�����j����|�b/&��9�������6��eo3����u@�tRI��M��8���۳�1�ie[O�ܔ0�jo�s���_���/�%�����7%֤<��5o�"F����9}A21��H�?Խ����"�}�˨��&$�(�d��������'�a�q�2�M��Wq������$[�R���z�>�b�B"�Yf�\q�K�rOC�����^_	��ݱ�-�u͒��ba�L��kU���#��1�17~O
nN�<���Q�Y�d���'���6�ԔV�X2[G���A,���"�dZ�}T=�ę;�C�����/yE�1��l~�?�GDs�D2a�������U�E+����}�7{��Ҳ)�
O3�����jv�pn�f��&Q�ZV=�e�N'<�� 6% ԫ~����}}�v"(#}���&��p!.H�������Y�u�f�
��(�W�i,)�D���"L֯��]��ZC���2N��N
4|�����M�HQ~6vPa�sd�'�w���1�Li�C�PIkXY�$f��wIZE�Hl�=�F;���0n;��xmAAy���f��ߙϟ���N���T�O���TK�q�W?��5� o�o�q8мxkҊPo����m`���x��k?�(�G,x��{��>;1Y�ѐ���ضO�baDǇE�-,xk�YT6x�B�N��3���υK�����*� NؙB|o"��ϑ��aa�S�r y�}��۰m�J�G��ct�|[�* �Z8�gC0����������ՈB�(_(��U�G�e�u�"��S�	����%�׉?�QD���$D�R�_j�6A<甙�i�a�?_b���R�j׀�Z�,1��P��n���&��!�*��3�lp�r`
���H��`M}C�x��C)ӑM0�T	������CB"�6�bKi��|��x��(#�?!.�Yo��Jr��K�A?�u���_�L��_6۫�Ժ�Ӱi�a�du^U��U���"kw�Y����V��5�4j�թ�i�?������Wh���[<Zjo[�:;k��Jl��3i���C�/�=���K���A�/�<n�l5i���f:ԋ#$���̆4��_\�k����������!8��G=�5����i���Y@�$EUē{�FO����}��J�+��o����B���p�������[1�� ��zU{n����` �����</��0�?��	�M�BʍZ�|:0)ok�M���y�<<��BF(;ܭ��mCdX�Ȗ"�+�ف�����Յ�n�/3�WS�k�	���ý+\r*V�A��OW��{�����;����\=��cB��-8ޠR��� ����Z=a	��0�s�>�!<.��D=�k	!�S�2��}U<T�/6(z�f��_2�S_l��'���.�/���=�k�Kv�|	-/�C���t���<	&�1%�S����ʷ�b�cކ�-f�+�t��ڽAr�G&{	_��Q�:��l2�6ײ;7a��W	�h\_ L��[�ci���>�ke���.z��C2^y��8�0�S�^�ϻ�c�D��aO��9�_F5GG�k�(��ڐ��E�Q^�d��y?�T�[8�U��oG�5���Ge�O�t�8�M.�͙se͖"u�v�������-[��/n���R�h�f�������Ά�S��X׻�at��̰���0(k������e�lX��(����_��� [ׇ�yFbA�q�'�j�~�5<i���y�y}�@$�NFBuMU�� HE%	�	��*wΑ`� %�.9�#�1�D�q�B�#L�{n���
,�	G�z�@v�y!�����8� �ybTDخ5M��_.���*9���D8q�؈20�#ײ5�0��f���M@ߗJ��cd�7�1����)�ܻ<��F��,U�"B"��=Q�g���t	뫺�k�.XUJ��.N�6���'���k�~#��s�aU��|���]�3W%�'<�B�lOH�@�Ө1���7���V*���w�h8~�}#����Y6 t����U^�E�*B�\v6j�yb��Ǿ �Z���LFDX	�^Y��&����c�4�K[��@?t2����@�B�P�=o��8����`���;�9���Eyr�b�:˳�k��l���h: �����e|��f��2����HP��Q�jG�oW��Q��B���eC��x�Y�=~��KD�Y(����YVl�����cat� �K���m��ζ���b�ko�P�m�%A
���A����jS.Ĝ2~(r�[�N|.�@M3ىBǊ͌�9�B~�:������T�i�uu��AuA./�D��N�2l0�6��^A&��=�J�/��CL7jz���D�x.6�$i2)�x�9p$���J��@0O���r��#h�ǎ*f�I�����"�=�&��ceTݘ���%#?�MP[�����%�g�g��
m�;G%`T���ae��x�jS�"u P�����!YMYťA��Y�4p�D��B�t�2�������X-��V�e�{�S^�Ǒ�v������P���b�{�ї��=S���r�-���'!���r��=�����w��7n��09��X��h%l���! ����/(��(�8� �C�i� =}s�U%
p�n�����e�����+#�r�<�k ӗ11�T��Z-v��t)��Ӹ���R|�z��:V�4O�1���0�1�&���$��CZ	s���#]3���m�y�h����
��DeX�Y,�{`Y����ha=���L6qa���h�0r|fC��׬j� 3}��U����Yt�14��dbx[�tS.3 ���<�:¸#�@=��,]e�n�!��\�V�\�Ϋv�0MW4(b�ݮ��xv?�`,�TW���"v�kԭt�N�N([Ĩ�uY�Y�`��%�0/)O���-W��ݟʗ#���"�SB���_�}� �P�y�f�i�-|M5�Pg�T�����~��d� @h�^�Pp�Y�}�m��dOSӪ�4�o(>�Te]�f�Z׻/ge���@.턤�/�&\�!w|��>��=�a�k�^�
67�b���<��v
M��k' �~�ӱd�sL�]�I~��
Z~�\]�.jp�&�Q;�(U��(J�[�"m��_���/J"':�ۍ�9p(�5�� �c(�p��s�y�f�̾����%Qw��ܺ'�T�cB}FV����#��EHKB����o%W��8���Ǐ�U�o�`ր5�*��$��
�_r��i�Eڹ�* S���G�@.�b�R��Q~`I��M?ǃP��`�|��>X���
�`d�!L���2�Y���`n�[d'_���w�[�dapr�6A'}���
-)G�RCM�����Z���bĸz|+�o4
m�y��ڷ�=��
�jմ�k�U	��ZO�Ԉ��K�TJ��CӓJ�"j\���3��)���f4�yeֲ��h�]r���q���C�O�ἴI�^���~�0s'�5���ƀ����L�-�|��[_kW�v�Xn���%Ak��i��G~N�b=��2�zZ�p�I2�b5a�R�j�s���8����o�M���"��4ORJ[|��qJF���Dcݟ��k��p|- �#*��ny��?�|�cu3�
x٭J��}�E�f��bb���7��'Z�v7��}�j���s�뀏(6Uce��u	H�'��K=+�Q�`=�Eߡ�[D��Yi�SXP�vzI��OW-!����[�c��#�l�n;�n�:Pw`���$;��Ú��c!t�'.u8��_������~!|�[���#
~��@���v6�ޙ�֮:���_k}q�H+�g�A`��u�y�a�M�x�n�X���_����y��� S˂#��7�|�i�Ez�̡����ix��@=@Z:�Qh�FL�\KfF&�x���Q@n�U���ǩn8���>�7���f}��y3U��>X�Ar��=��M2v7V 1cTs)E6��_ c�N �N�$���W���}�OFָ�;ڃ��E���	t<��#t��x���k���u��k��㿴Ů ����'��w:���3�( ����T�Z)���(���X���L��s��E�XN8�扥O� KD��Ⱦ1X7כ�
����}�7)`7��>�U���R?��0���/�8Z�h���*�a5U���;�E~saKe3NT'`��e�U�(�sn-���=�M�m��H�����mj3��w��Sߚ'Y��|.�{����^s;�8tN�<���.i�Ё�Q�|�S�����h��(��?T���!���u �,���Ҝ��ҧ���|<s�xVZ���T���.��ɴ91)v=�v)��-C�o���=)a�iQY�����<�⮱@���{��Ȥ��AP���H�l}d�v�щj}��u�E�P'2�4��` �����;��K*sT�}V_k�K���f��^?J��c�D���t�ﮥ����y��gO���Q��ʇ\�b�4��V�CWa�g�G��b�R��tK�����0�@�&�6J�DX�oR݂�W�t���or��,�;zL�͗�����zI=��(�`C$�v|վ٥�:�3�t����a��}�1d�9$�K��2�5Cz�Id�R��ĠS�Mj�#V��7��X�p:}6d�;�&��f�9��<XS��R8��i��q�H��B��P]��.��#e�n�ԗ�2/�7��C��ү���3�H�]��z�RcE��+7Ts�0��9r��Z�Gh���6.��pJ�C?q}m��t�x��&oq�5J닦�:����g��u"�]�t^�����Y�_C5��ᏹ��[����%���ؼ���y���J[���n�3\��
�*.q=ow��
�e��U�R��!�rS����i����e3T@ל�.��m��y�`�>�0��j���j�ҪQ4�&�]��e��t�<��\g���2F�q�vZ�� ���Vm˂b"����~̌�正w��<�:*����nd�"�\��`7����L���z#�m���t���pM��h[s)jdqX FD�5���������s1] %Kȃ�q_>]�z�J:o��NvH�~��� G�5p���L+তŉ�Z[�׃�����2��@�|(G�"��1�(�� ��p�m����-5���S�_K��4�ǁ��s���*m"K,C/�ux���|:��;�����L�)vZ"�M-��x���
֏S&��3�HQ�rW���V�8�49�}����0_i��.:}��+R�)�#8xu�	vZQ��j��4��� �.8�e	���@6��,?TM�:��A��םF��r�l�L>�'��T)����g,` NU��h2ux0�Y��_Z��*R���3��:�����8�Jîe�F�a�P�u[�x��0PM�?C0�)`<Mf@lB��!���EfFf�=B?�Nde^t�^�w0Py[BW�1dr��l�F��!{�ih�Sm��݆��:S����e�og�<�ݑ`�|�Gߙ���Jɨ�䘏,�v��Ij�5��S��ǰ0���|�מ�c�Q�~h�����i��9���zן��'�Н`H#$��%��6"��������cl�
gO!3���i�[���֊�^�Vt��w���Yxs�{K4�uG_���� �@`v}ns�(��h�UR@r�8�UTN0�%������/��[Z�g-�f��g, �"Ojg�8Hܐވufː�-:��^K�C������e�D���FN@Sh�n⏂l�?������������R#a�(��j�.��� E!����,�-�e����Z�)+�o�OZOJUP��+�?��=��S�r6K�]��Ft���|a��FQ�5����B�}��n;�����a!ŉ�&pk�����뾸T����xڌ�MG�_<��@��f�X0jy�vޤ�P��0�����[,t�3�^`+}�M[��:���8������Ɩ�X�� �3�,�R�8�zlS����#	d��г��#\��E�$���-��?���\v�*=�~RN~�`���_�pc�ȋ�ɢ` �g琷$�Z��r�7
�MS��~����l��C�*9������M��y��+>�q|���\fÝo/r^�I�W P���~�\�@��&��9Z�͆�n�[h�5j<�ӽG��.�B?b�)��I��Va5I�R���J"A���ݟB�-3@�#C�+��������Deګ��i�MN(�`v�#^|; (Y���t�AyyE91�n@�����f�� 7ֶ��Ǘ89�xL�b�X;x�k�K&]L���z�e�zn��S������\���$�_-EjRJ�_&R5�c�Fų�;�2� <��BP�"�4�J�+�q�E|V��31��7�w���8��Z�r�����xv�d�*p�JW���p����r��t���^�#�w@�!�,X���S�;�'7�E+:el�%
��D����W�/~_,����t �^O'Mc�$<Q��*}ZG��=���q��
��|5���^w�1X�G;�9��u���~�w�3��_��l��y��}Bl5�Wbs���fe����"z� �����'�J)��3��@��E?��4J�%��jqX�L��,TO&���e�m��U�����P��rI޳K�E{/ap��F��K�e�;���ǘ����dЧt�y�P9O���z	,n�N�IO�ō5�G�1��\㊉J���o�lTs6CLGy+�M0{ /�]�3@7�d�B��I~��1��������������!0����K�D?�L��������nxQ�4�Þ��B�;P̝\�6'��Q�U��F76Ze�s3А�ل{���o-��������~�٤�z�hp��*�a���z���@!GX�3��N���Q�%~���G]D�j����_vZ�98���b��H�+_�?���I��EYB�`Ƒ�5.�6���.�C.E��:�w�aE�~�z5E��m)�Ś*�_��? �lL�M�ʪi��\�_;��PG�]�ռ/�>D�+�'w�ɹŗ�n�L�[`r�a�h��������Z�� .���8��"x6�-���y{���+�s�q�C�k��F��9��ݼ�Fw�7�?�t��Ѿ�Fڜ��>�Ϥ9��]�?��Z%�L�
$3A�փp�'LݷU�K���
����?�X7��`�������s/AR��BJ����F���G)N��RN�Na�p��U�����bE�P�1~S/j�E)5�������6؝�<�������'�:)��1�V׫%f�)6�vtP���qS���d;�V?�~6~o��C�Q�J�b�R��H+qDo��ȏ߇ș��z�gl#i�9�� ���� e����#[Q*�.�Ty����觤�So� 5�y~,��>n �$�Z�4F����A�97�긇��7� E#vKC6��!���N1s);,`.р��P���غ����UȦ��M�q�%�M�?mY���ì�jh�(ʜ�0��N�G��@�b�NXA mU�����.�s�`u��s@|N�1�� ���
έ��"�/w$�s�N�͐�&��UG�����~r�<�$.cى��56�]�����[�L,�h���<��Wћ�\�<Z���E<����� T&x�V��@W�#'s�-�'ek1�ٺL�`���9QkQ;�N�]�_��j����	����3=�/�����+�� ��U�po3�s������	����JȨòQt"�H9f�o�e<��)� �����9-wB*�n�Bϖ���`��>�2_�}`�s�3�m���/OfK�Ur�.�D��K4�A�ruUO�����%f
:a��iC�8�1��L���)�kT+_Y>�rt۬����Z�I����[��Zy͚ʲ���a�N��͵�9��M��cHI�����i���@>ۣ޻���k�0q�[�,lo@��ȋV���.����%˽�F��*�gx��&J��R�t�C���Vw`�	�dja�y��X2�01�@/�N���|��l�8�֒>D�A6��6ds7���K�2��/K�dɞ�r�ѫ�e��� �±d�����K��ZW?D��M�̽�vÖ�2�o��cb����IpFj/X�Uc>����*[˰
���� :��]�K옲.�Q�>����DYJ�R�x��6�u&��V�<�;c���ya�ȲQ$�x��$/E	��4�┺}�?w�İ�'Pr9�b��CԌ@���RʯA�V����+�����lb�"&0�&�RU�밡���K2�Xң�D��춑^�x(�}��f߇=��껒q Q�vB9Z
��M��hO���ӄ$mLh��,V=�v�&OJu {I�O�E��F��Bˎ77�pDJIcwq̲R���3�fBU+:�x�6!�����y�C�����>�㌴�CՈ�E��)�5��C��^�h� �4I�|K��
 ����1(�-���t��V}��kDvXj�x	_뤹��/(N�C���eB����gWH�X\T洹�0.'�o��������Oε�8?1=�jΈ����kw�1�,�����/V\"��T��9�u��-6B5lj�
�Q���vSphO�[P"�� �HUƿ���ߖd�o��BF�B���8� �~�K��(�t��N�f��С=�ߓK�i	�6��o}A���� �6	�OehR��.Ҡ�s�{��}"1�!�Դ&]���HSԝ�ge~/W1O���|]S#�KI��rG�N<�)iO�g�s�#�H`(�ny���褝kթ��P`�NX\�%W��|�(�ev�#(�6�x�XT���)���j,.�]Z������a��="8�_�GI����z#7�~�(V�9)��Y'��
k#��N�%R9�_��)7K0W2�v<����Mu�������P8e��[^��79If܂��p���UA���e�6�qO��S��K�E߷�_�r��������Y��������V3�q�*��D�5/������D��)ѕaN���"�
�����j��VEyOv��Ŵ��\VFvQC֣�����f��w��U�n#���,)|S,!9�ޔɼ�Q�r��D�w���e8ѮD.qb��X���31�����R����I�̗��X�����8�^(�v��h͂WS�Fv�W�3NU�Ė�l&��*���HweڏJ�/!cLӶBK+X|]P�Q٠ٵT���du�lD�V��d�EDS�m���� ��n����FQ؀�(��	���l����R8��g�8e�1��y-=j-S��4�/�r��F1����Be���,�<���#�������w�箐��
E?@��f$ژ*����JFZ
eS枴��F\�.eJ>���"���e�}θĖ��sL��&�y��45����졎䩘W�CY�:kE�W�;]���8��I��]���d���@L/�0�_(��j9����s5���WS�d@ �]�,7OS����w�>���@E)!�1����X�^I�:)����`�Ag��-�ۘ��j��*�E�Z<l�p��YF���Ț����Y̑@JL��t͞��0B������;�>���^N��tlR��6_�ѼG�),nU��mT��>Y��%Uտ�!����t�_��!����I)������I�;t��0�M!Uu�_!a|�U��!�;Gb�y�@�����Y��u�%��qM�V$�yɀfnk8��� ��q��3ab�".|�D��4�m��t�}u�Y�m4(P�����(|��`���^�4)��=���c�~C�_X[��0�)n�U����zJ�3+ةzlQ�K��%;K�hH�䷄��J=�WG&�"O#S�� y�Pv�{����R�[S6��|���;���( �%T# Զ�FKw]Y�p0��B�+1�4��|�޿�;R�֓>�`�"����Gٜ�B�	8�����b���}7�Vp�7��=�;*�
Xa��1�����0e����s�/d}��=vJ���!�=ͯ,��>S��,T�Ɍ��
]�"��B���7��D�/AF�:gÕ���b��j֢K�����]`����6�љ���w����$� ����wN�\(�`���ۗG�g�h[�t'������x1����'Z9�ؘ���Y��F�b珖9*��J�e/\98���۵��䉼�7�
��|PN��%�.��@���S�v��t����~�op���|s�ɕ���ߺ�#Y# 1�*,�7��s�Q��"}������$B����SN�L�ꡔ%��-�P��ۡ�=�>��
��c���ڻq��W�	�d�=�'�Ƿ�EϢ��
��n@XF9�LU)NT�t��RO�'�p�8r�����(�5�����@�w%�)��o
:���[�Q��0A�Ӈ&h����kD?ږ�{�:�1�8ӏ��!z{�,�V�vWw0U���5m�\�l��/;��G���<�X��Sz^������Ԟ�<�s���C
���P$��0�ɘ'*�����+Ţ4ZE�8xѓ�بf���Nd�>'2�ˏb?f�� ��b�!`@K��I>��x�%"�jW! ����E�ɷz�>p� =����B�H�̠�k� ��|lS�4��L�+,���y�Vg�j����:�*4o����o�\�`���%V���{g�9�U��6�5��X��5������m�s��ׂ�%�%~��[�Gӎp(e!��9�ִ��S.ۨ�9_��g,�|dݔ��P�7�{3P�Y�j�����vW_�ˊ��&�W�85��[��_|���:�������p.y�d䆽���_�1����6�䟬q�����[fq�X|�"6yh�h��{�y���>��Ⱥ���x��:�¯�L Pʵ�e��tJ`���Υ8l~4��V� j%����5�8�z���\y�xE�'�.w��F�C���;|����&�z�S9�%�@�p���;��o�ט�c.&V�=��P�+!WK+�1��}�쩕�;���I�.�����5�#/��2�l���M�#5�j	i �cdj37����}�:|�%�����,�~�
#%�X�E���#hȳ�-����	A�,ǋ�j ��#��TPG���I�P'=�7m���\�?���V�	��#�$CYdj��.�"Vnu����UwQr2{m�����8����;�e�y��ȿ����J���m�󾯮�(B�9f<}�m�eo�Z��7��9l�9��'���_E_J�9
�"�P�X�58M�ڬ��ƲP�S9�������	@�ߚّ��Eub�]m���X\4�O�߉xC�&9R/�A�f� ��|25v��i�hʆv�\^�?l��ˤ�|	���D{�'w��RC���5NWo��â�x�Z	4��ƀ#tG�����h��S�nC���&Tb�a�	�����\� `�������6`�hb�b
��ޓ|ghr��[ƺY�����D���?&CPí�Q��Ll�<�w����]���\{#�2VaYzP��*u,��^�<ec�=�<n0*�+P������0�v��5��Ǫ�Ҙ�@�ĭ�F���ߙ6Ye�m(�r��=�P���7�����E�����o���y0:�*i��L�?O�C�Q��-�kB!x�v�MZ���x�ֹY�D�8��3��m:A�x����q3�[�,��w�GWo��k\|�DI���vEڠ���}�ō�J 3d�X!a����5���%��{o�f,&�_��;g�6N�B����twW�����a/C!���	�
��J�#L���oe���,��{Ff51�Ɂ�~�Wr���Xm�bq>?����Q#rb�OT����'�s�|��j�r��hn#�'2*��[�"QܨQa��:Rە���ώ����!v�����¶���Q?���^���^��N���hK�"��S�0>�[WgfeqF@�wÎ�������~�u���^�\j�Չ�A����>��OM��EDJ)���S�b��BA����a��a��ȗ�`�DԕS�Pa�92��kf��]E�^H? �^2(~�����%;1��#R���_� W����k^�9#^1i<����\��B3�G�ݟ=��$�KO�)� ���{<�����;�vd���Ɯ��8zD�蕳�p:��k�K�o�nu2ƙ\�� q7eMR�]�����4*\��m�Ӯz��_ץ�k{�`��L��L�Jtz�]h?��l�O��xS]+���??���Ƿ(�@�9�]���p�SYE%��'�`��
�Ӌ7*!6����gZ)��h�n��74��L%�o&�۪�S��fj>��"���3r�C7?9�k~(��I�wq���8�L��t��j�_-)���g����Wb2�O�t{6��K����u�]��+֯4R*x��ڨ�1ZV::v���Rk9��Мs|ZX�H����7�Z2C8�rz�0�R(����s���#�*Cլd��}7�en�'�)�b=�g�AW	S��`'|��n }��bk#����Į]̻G����B��Klm#�~n`e��u[4��_Q�,x�i���!�l�ŋ�L�=+�iζ.������X1����w@窴�B����VN��pN��\1�sO����&�
t���)S����Y��Ba�.Yq�\ ����BI�ݝ�7��EM�p�I�E��~"��C��^yM��)]������!����Ŏ?�g斦.[�>����;�hJ،"�xR��9�F��6�bt?Z�Ս
��L7��%�n�� C�M/�[���bF��/�����~j�&�8�\����zP�r����2|��r^�{��F����
 >�3_>6r�V��t�_I5ūp�1S9�E�*��L}B*%`ύ�^;R^,�Dq<i{>�a�8�[�G���1|��`�f�+�4v�Q�R-����
�}���ZUJ����'�5tԾ{5����_T�N^`AE�"��QŢ-Ϊ�ӝz��� I������%�o���G����,8�yֆS,�VS�sk��?�;չ���w>�� ��ݽ�ok-{�Ǜ�=�j>b�d4��E"O+����kTH*h~��������Á.l<�:4����Fow�ѐ!ʐ_��-u% dbe�'�������d�B�P���h�i5$~����O���G�� ;��ia0_�qLe�_�� I@o�ߟgR.g���y�S��Z˼Lq�V0��kmmqAg�w�Zo�a>���(%cW��׳U)l�q�u��YϜ�hr6���7���j�vAv�� Hڞ�c��9�o���=��#�Z�sXB��튈�64�&[q�]1��`�?�Y����r���W��E:��{U��� �ʅг��!y^G���h��F/>�´�i2�n�UJ=��q~0���1�[���-9K���H��C���nה6���m`���� ��"
��V}4WV|7����Bp��� ��C�BImU?�,pwԭAե�˰��k&��4�@K��J&{�zAJ�=��[J6i&K��8\`�OM5 n$�@}�"����6�i'r!����ژ-�c�*�p3��<����Aj5�Eչ�C�~��� �+��t����B�DyF��;��)=���ܘ�@�p'D�`�Z�̯�>�F�6�P·'�'�W+A����A-R㉓%/n����Dx�������x�����Ȗ�;ƪ�oI��q��	ke�f�Lg�����5�4�q�s-�=���pW/X	?`m�#�IhL��$-�^�YN�~��������ih]K@�3<6$��x���N9m��*���ۍ{-f}(�EU�������H9����ã��`i�-b�5D%�+&7���.��P�O[�Ev�`�$yĘg�3g)` YXQ��5���c�<.ꝕ�M�щʛ̄au��):�w��/��(�V���B�.���Z�FN� :6��wݎw��Qb��;f  �&�s/�8%�#~':��T��+�on� 5�e^�lֳ��غ�� >� ~�Rv���ǃ����=	N�|�كv|Dc�&M�7��j�����2oe̙㰟�vȑv�^�$��ǀ;
X��de�QE:�a�ґ��7���\��f	�ڹ��:r!�e'M�.�B��"����P �/tp�cHKA��*+�p�>3ze��QZ�Ѱ4Hs�������m�R5��]�υ�B�)k�eJ,������bj?+7��U��S��(?��4g$Bj��\�\tr%����Q��F�����(���,�k�L���>�����U	�<O)�lT�5u'�^+���n��@�BY/8H�FV�X�4#�9�̿�y�ծ�ΖSz�D��[֋XA+W#����#�bvήI{�g������)�/�nvP�r�����`�w�*u\>�3ܳ��ȏԨ�m�wH��@[Gxs�y��0z�@�$����
�l��-*UW7����jy�4����h˧��G����$Z('�G�8�\7���7�\��#����r#��?:��	��D�t�6��6A)l�t����=�g$~O���
X��5�R��J����}�9`��-�[:���I[�V	M��H��[	=�ϒZ
ƃg��!�e�}Tf�9u�Y�3sE>���PB]_�iਫs�KL�?��ʖ�d�{3\����� A�E-�]���� ԛ��V���v-�r��{%H9X]��ۊ*Xr��P�Ȣ�h:<�Mh�ҟ����X�f�*��ww.5�d�qJ���kL�x����Q	��:a�^j�''^�����F�D~����T��Վ�� Q��".��?�V�p�m�w�vo�V���o�e�Gl����{��{�^݌i�cp��V�=��@�FL��%�٦i���7�#ߺ����<v7d�F����:T�ٶ�t�"�o$YPI����+�y���s.����0ր�M�if�(8�Ó���bS��WR�5�d���\,DLv���9�{�8��|4��D\����RZ,���T�<+�4�ރJ:X�!z�F��϶+��"����R��;�e2V�}֗:�kA�B�\�6�{�-����SH󅥲�'��L���։�n����_�_��6~��Ղ(,j�@C�I �4N�X�N+�)�H��@܅�ad������,���ϊFt�XQr8j���s��V�Kq��V@��CF���\;���ֆ�P�"&U��"PRĈw*����{U��Y��a�a���r�����c�+�6׵	f/m:�aa2i�xT���jL�-A�	�
7f�|a�#(���-7�V�ӡ��>?O�d��W� 6�ф�כL��~��)������� ��C�q~�J\�I�%��,�;ҙmw_<���)x�q��5�S��C9�������9�/��!S2U�i�i�Yv�q�s�{��(ˮ�wT\P���U��?�c-S��Tw@
�<��~��n�t5��gV��erO���F�4��gd�r�x��:t4=�'�ㆩ3�k���9�(TL���}fS�/P+����`(B׻	st^֙�昺��?f�b������������������?�}	�vo5�w֬�R�'.dxG��O��5�2�
x�p����� 2QX�G��Fn��w=l�l:�F"V�~i�mJokb��J��V��V=9v��^;�U�is�Y�9��I��~FL��>��z�*��P�x���8b�p]c�ӱ5`�_���ޢ�#����>KL�����mx�|LjTS$�w�ӸC��~��%c���x'�� ��˃�*�j$������i�i)�щq���8z��5���vU������(��������BwX�ѥ#��Q�Oۼo�����G��$*��@�>�^�������-BS��fz����U���\��X�K��1�.��%����w�"��;�)7J���D��,�\�0i��?�5.L�E�*r4�r��茝��WP�1�|w"c�b��py�S�*$x��� #��7W���c��P�@Ԕp��0��N@#�g����9�ͤ)"A��!�ZB��5���-a����^��Ϫ*)��dz�ݦ��k�q' �hi�;݆�Ǻ.ԑ� �#��o�yJz�0kS��&i.�I�t�@���J�[�����</'��;�.��ɹ�-�UsY2�QB��ˌ�ޙ`w�dgQ� ��:_^�R��;é�y���)�T0��"P&��(U\$���**q/��=5�mf#����զ�X'�=��2��V��uk|�����B��UF���E����Xc��!]�+����K�̯��8�� �"�I<�V�����A�a�AC���$W!!�@�8
^��s�S�ό�l��k�Rd�h��MTi&��B�a8n䡴 ��)NqOH4�h�:{�+�O�Syv,���6�~hԍJ��?�!Q��^�Җu�1���~�Y��9}�����{C�������;�S@��v��-m�T'�����%J����	k�M�`�ɉ�IU�LEM��NWw��/�m�:Z_$�������t��S!���*@�7Bax��q%��z�N�$�hs/�F�"nF��M��.���,±@��5f�k���C�|I`ا�~����JLDE��Mŗ<�Ox����;�0�N���-G���{��Q+����ñ��}��#;�d�P�	����-_�{����8��+Ca4�r5[�	�j>OqB�C�������_&��*��sm�(�Sǀ)T�%�|�ى�9����q���¬"�A��46���K�`V4��;��2N��ji�����5�J?���E�tf|x���RD��H�hC&��E;�݂��
̊�i�d�K�w/\�ېh�dX��I��E�-z�-�xU=,�L�\A�Q�K9H8(XE���I�$�I�t�2�g�Rl����6�@�Ü�Ǖ0�]L�C�f�7F�sW��YƉs���K�E��nMdδ{�������)ZS.�r� � ���Ռc����o.S:��I�ÃvH"C���BV�W^7��f�B5̑6]RU���@���{�.�~/�wEc\��`�!�th^��,���O����l>+�0䒐 �ְ:��odSȅ��(��<z.2b�C��M%���*"�n��It����FX����`St�H���Դ��Yl�
Ƞv@3�U�^?��vg y7T}�&T�h����yމ�v#ލ�B��Of�䷃`�h|�IH�*��DQVk�:³�����k �ڬʆ+�I��"�/����*ɜ��xE�jڃ��V6�&\K�ǑIC�fJ��Vl��2���y8[I�a� ���{6�/��ˋ�u!��7G}��3G���k�~�<��mDc�<�P�V��k?�|����🪷��\�s�a�$3vɡ���k25��몸ƃʃ���W��H�#]�����"�r����;q)�o컪=�mK�VW>l�-*����%x���ח
�Ά�ݭ׵ڤj5�<-��9m;���:��I�������g}�IY��bE�9��R��<�Q8�ʢ��v˿�ܨm_T��!;|�*�M0O]� �1KWwꁊI� ��^�˝�"G��k�¦�!G��v�R�����k��"qnD����3b�2����J#�����c��[s
$>���=�x_�Xg��P��__���$�m�0(mH��� a��<��=�*:x3��ŏ�O%4&d(9
��Xr6��ӳ�n5%�D�m������%��VG�x��e9�`��M\s)����,��o��6�}�걈�N!O`?[� ��-�#7a_�;��Y���B��E7��]�5�jS=�=�J�5 3��i?"�Q�u�Zn�Ӕ`��*��0��H[
(��}b�,��0we�)����h��q��-���OK�ڏ����](G��F�5�H�/�k�ق���璥��ӭ�,�#���8���!a��	���k�ي745M�Q��?Em�9�@�R�Bٌ��*C�S�l^I����c�K��*�᧮�x�G��E,��-D�o�Ļ�?&����_q*<��:�JP���>��K�5Di�o���S0^I� P�V{ʑ§�(,�AՍ�M��NR��v�r,&�S�G`��dچUԲ1����(�L1�qc��^Yz��d��O�O
��P��"���m�XV����'��ວ��w�!�R���Q�s�����EC�:��)[�2�%
�N$�O�^���m�W`��O�So�������>
I��?/�xev�#�?�BZV_���,�N2n�?�g��w8.|�Ӂ,F�b-���[xd��|���00-�eF�7�:/����Kd^���(�������F;!�)�D�F9�з��S�}��@��:�ZA�8N�Q�1s��:q${|��s���"�R�U��j��J��Ѯk���NU�|5���t�~c��^mbY���;Vf��z!�l��������.u�M|�����vT��fy ���+`�W�>�U)�kZ=z�ře+�!�BF��m.#�(:�v-���wz����u����q_����F�Ò0k��QYP��bb?At3ͪ
��sY�1�'�s=�6�fr�-�A�ޢ_�u黁 ��w�q<A�w\S���
+O��gNNJ�	S?�x�Y�]JR�2�ўt�E�vW݀z���5�f��p�e\��"��BL��u$\��:�FG�2��v��ש�H���8=��,r��N�9��g����<�P�G�B�pU�5��b��ݏGA���Kpå�9�6�N+G���'�.blk��G�F�u�n�h �Ŏ%p߄˭#���X��Å�=���<�a��xdh{�Nz�����l:@i�孽���L��6��A���c��5IPSؒ�,�|�

�i��Vm�V!h��/���QW��H��.���Ҏ�_�hB_u�ּiu�z�oNv!Js�J��\�	"bw�{	���4xߋ4J]聚������4�=$"T肭���{�6�}�ն�����t�,!��X���_6f�q�q���t����@m�К��9�@�ՓɣN�zy�x�$�O���|%�@ɋ"�_��U��˲�
�n�D6S��*ͣd��*�T�?�q�.�#�`0I�ϩ����M�"��a	^�8�Ԏ�A(�.���S|�@���M=�
�]�s���@�p�@����p�Y������8ґ�<�:Y�aQ�5���m��`û����R'��i���نhŮ��Ur�e#�(� $=�Ϭ��N��8wĊyӶ~nt�"ɈfV������

��g�ŋ��d�ޑ5�<8������	82�%:��̰xa�QE�yk�>[�|�H?/��x�5��M�1��a&?�����2�m`?�~�L��*�.� ��:Tn�3ھ�����ވ�Y?��y�;{W��Hn���8� �Q��P���`�Qpo>&{�<����s��Ƃ3�/͞ъ��zV�cQ���d�����T*фIjkګ-/��+Q�|k%w'&A ��]�ޘR�i�7gP�UI
R%�Pvj�Eq9{���)����B��{��:Kݭ�:5��*�ǐ�	6��!5ճ�	�˞o�~�+�1����Г�� ��
�,AtW�L:��I)D 	M���^2�-AK���IP0E?Zr��1��"i>
N���Srڙw<5v��W�,
�"�D�	���{�\�v�Xn��q��C����qŬ-ާП0�	{0'wF�����<$[�~1}�5���GX��m�.b�ٜ�Kw�os�pS��DG�,Q˒�Ź���R~�5aW��HF(M���$'�0
M�?@S}���@	��д	F��1#��SGG�+c�F�m����7A���/�m��,i����G.F�B3���9=s��g�^��k�O(�K���>����۹�ny���:yz8�o|	�.��cښ_X�·�9�5�r�֚�@_�� ˪%]�B:5��0�,᳢*�ʻ O�}��,8\5+���Z��5c��L1�Q�zջj���A*�R}<�J9��������3��?��/��rCe������5OW<[��;�l�ڇ^IН #���V�K��e6��7ᇂ���<�>-�la�JϽ�̦�:����`p��`�7:I{Q��:�u�VP'��a���R0pe�1\s�%~/h� �j���՞7�� J���\�ɐ�_" %z�]���<�N�?��O�x��3*}/|�>�nY�"��n���rHX"�]r�8�!i���#����54��Jp��8�Yn���������\�'�4L�='Q�	�K]�r����(� 8�z��:Q���EEu	��"��ߧ�*"��|,��������%�ϼ�T=C�}7Q��J9��89�y
��\���*��ŵ�7+j#��ǌ6NaF�>f�kޥ��#9�O��|H'��E����g=+��	�t���q<#7
��Ѵ���� ������¥�ٰ�+�v�&���5'��`w�/O�E(<5;��U�깾eY��������6�P���nFI��|K�CH���|JK�oήټ+��������\��踌 ݃ � �|��:Y^䓑�CZ'D�
��ȳ�Ӱ�>Ơ�?VM?�|Ͷ5�#�x��Xe���W�����v/�|"H�P�B׫r�_�t��WW�L5n��;Mk�܏�F��/&��fZfJ'��c/L!�f�̹�q��6�/[���O��`g�ƫCIz�4���>�;�[^��i���q}�
�n'K�P�,$��Ja�9���ha�c���q&틤�����[�M���#�6y�uׂ�g�ݛ��HǾ{�w1=���_ϸ�fqͩ݃�y��_��u!f������)�e�q�:U�.0Ʊ�)�h\k b��ӢH��uǳ�b���5��	��-�*�x�	��
YνE�gXΨF��V�����f���9y4S�o��Hk��lq��n]���]��>\���<�4ՠ���k��vWI���h>q�)nU��W�z�,�Ԗ����;	����*��-���'�c#�Y�JJ^�2fL�=B��Kj�5�
e}�M#Y.)���4���@E�վ>9Q�dB����ak�ꤔA-�	�1,��a��A8MȽ��󋖃B���Ae$��Ûmv��b�j^{�`{/G���<��J�w�;k��E�E��0�J8����xr$�����΂�әɦװ�DtY��˿�X�E���"��A�O��lj����MϷ�P�����eT�v���^�v�|�:^�d��0��$i����������#n�雒u�u�΄���꒠�S`\r��$'�P�.vlz�V�]�ޣ��86��F1'R���MC�;`+��%:._���U��aa�p�LC 5�N�A���!Pu>����(e6W��%��I�껴�@���,�-�Gѥ�Į���j����(���A����Q �U&��~�.0�Ȝ�Y"�3|^L�	�Ɣk���r2��>D�U�ݸ��T<�%2���%��E��[p���9�{S`Fi��P��¾.��H���/��ۣ�̰�0y��{�b޺Vީ��8 �%?Q��p9�f|�17lf���oޮ��P.�)��V,93�9��sb��!��⸣(5*j��?V�n���c�pAE���|
�x7QV�Y�*D��N,��~�"0�T,�����Q��r�n�A�e��]ޅ���P����99�y��^7}�o���L���g�~8	�I�r�:��ѓ�+k�"����NPA�e+��
Gg�J��d�$�q��p;�S�G|;�RE�.�l6�$u?]����;����ZV�"<!�I{7
��`N�٧Tx�`�n������MRA�8�����P(������<�I�58�6�\���uf
J�(�h��aE�'z��6?R�z�B̄QK�c���N�L*��Ď�Z.s@\��J�GNZ��6JC��V²�_o��=�J }�o���R��D��S�;�������m���O�ԙ�3VlGHq�}���+ί���>=���;�r_Nv��%J�g�лJ=�f�����G�����~���#`S���_(D��!���=��r�#v����P���x:BƽB|����
��" d@���Gq��x�ٯ��q��6;iA�sR���Ɔӣ:� 	}�R�ˤ�4�<{\}�Y[��9G���۳?wU�
��/95g�$�B-
���Jßu����aN�� ���ħKoeA<�i:����i[���0��*|�?r�7�����`5c!�,�Z΄9�NTv������S�9�g����"&��l��Gp��N�Z��D�)�ᔔ~�M����p����]s9X�|������	�Fa2H8�����8����WCf���1"��o�\��h*'�G�ZE�?dC����x�䯪��������&m2�|�2�a$i��L�_���W������,vm�%HV�λ��ǿĕ�A�v�᳴b�h�\X-kv�P�@ 	���SY�c�E�U
����0,�lm�ҕ|l��a9�Z��) ��f�[����.u��n�6pL�i
��g�{H�w�
G�����a����݈3Rt�Tw�AT>�e�k���y�>WX���\�����*D��a��U)���0�m���[�󔐟��/���$�u�[�8��u�H=�Lz3��"���i�m���f�T�:q�����yO�#Hl`(Ӭl��-�_�Ɂ�g�՘��sJ�ϥ��G�S�@��N��!� ۙ��y%"�ⱗ��{4������LЄ��GdD������ɷ^�-�Xkm��;�5�#c��-��ߝ�M|�o��8����h��E'��3�Ö��?��!5��D4E=�(ؼ[0���d���	���G<�m�6Ѩo;������"g,�Mؚ�£�_$�Si�z][q��ZP��Я*�xf������
���ך��$��v���^f�L3��zXr�Jr��5�Pr{(���z-/�k�a�dz8��<dڌ)^�CgH���@���Xn�.4��C6�u������}_/tʴ�e�)�/6��2�k���j�j��H�S�(��  �3�9p���\\�x��;?��!�}pd�n�zN��ȭvZ�&����ᣀ�h^�V�g���!��B?��3X��eYΌϕ���.~��k7r{��x��X+��~��¡E�= �Aֿ}��p��SB��!���.X�AX��S�:Ɋ�&�}��pJ��p���믍�u�p?�+��
��S���<a�F�To��$)�~��IcN�T3�^?�F?�(�_�^���{62C;]ܫ��[3��UH�X����b�Gh]�~r	�& �f~/3R��U�nnu'��cm�#=l��I��&���CKs��R��Ԡ#�
�-��թ[⮽c`ܱI6vR(6��[p�vRN����B��.D��P��n���
J�,�Z��Z|�zP��(���g��%G|�Ֆ
W���߻���5��aǄ�%i�2�6�(�6��
<�[�^���TK���j*c�ct��֫`-���W�i���ٚY��Ѱ����1���S����Lb�;�z<<�v�6hVl�Om�D��T|��
G;"˽A]�6Q��8`�a
X�j���($b:ncM��Vs+���273ɮwa���U�&�R4_hk�?}IH7���D�L�8�\P�\������-x�#� ����f�o�+o��m�l7��@9�zc��X��+�WS�>�a�L����a;ē{��0� ��_���a;hׇ�Ru9ew� Q��3��~G�ja��r�B4N�S;&��ƵR��8O�~�d'��K����䉔�������F��K1�p7���]&f��B��~�7�l�oPp[�%�fT$�A�%YaT�z6��M�p���c�.�yW�^�J��V{5\D��`q����K�l7eY��E褏.�;��L/R�T��U�ĴՏ�͓��	_�X9���$M۫&���	l��(j1F���|����C�}��{
׻�)ԙ³�@8�es(�$��Q�w�j���y�ƕ����ak�$9؛?*��G�P��E��O�p��K���2���U'r�F�ê@F�g ���0"F � �Gp���i�Ж���J����s��������=AW9�)�|WD�:�@pZ�Zi�^=@�� �_8�@�g��g�L �����&���u:�����6dl�^�zG.Z�4�agI塚##��{�Hq«z��|�Is�l�M���&��@�)��<�Ѵ�h��jz?6_9xB�����̻�JL����@�_K'6o�l��P^���獷��������t*<W��$ ��fŽ�fB����Ǒ��t�C~�}'�p��m8�8��̗�d�Cӫ�\��L�� ��{�����T��A��^_w9�%tYBU˺1<��\ki�,g�z�F�+-K�q"�:��+���y�t֢aY6���6[���-x�X2�gLV����0Pk��Dq�R�(�q�~�+Y�S���z�F��G*p�\VGN�f�l�m�ɿ�a=U%x�7�ޕ�:N��8���P�D����9 9�W��y;�L=��Y6�e?���*���B`��?5��f	����o��k�:��ƕ��Gܫ�9���X���/��P�P�~#wί��H8b3z�c!bs?��)�V�+��v���{�i\>ۛ��e�(md�v�=��g-�U�A$W���{�Q W\�g[,��5�zĘ���2Bѥ�Pw�����U�T�r�sSgŗ�Z$+�� ���Ns����Il�������I2m�n:ل��bȽG6�vȎg��֙��}� �����-A*|�M5�(��E��ꚞ/\P�_T[
�U��
Å&eAT��}B�3�bD�R�D��w5F��� ?�)� �4��;�*tĪ�o��Q�RK3P�ynu���M�|���Ty�^�i�t��OW���~	����!�s,ET}�Z]�)�3��c�?�0����������&=���6s�1%��]���~x�#�أ�H�f��ye�`���P�T3M>g�h��h�z������� �><��v�v�%F*cM����N�U�2W܆-�}�ƽ�/�$x� '��q,�&Y�ǩYr�g�����_��Oݫ��6�w��#�eo�T��8�$�	��Xn��爸�$�g�)�t!',x }!�
4'\y|��lmD���7�0��v�sĭx�	u 
����S\��BUK�U�×�g������^eO��=�|��NzrԿ��h�5��be �z���lI�)��'Lų�l�li�-'q_	.X�ea��jk�sO�����&��-^[��̄'�7u_n����V��i��)���;�VϺ%���j�{$���Q#\��u^Ӥs����T�S����Zx����"����_�j��-3��f��� Ȳ�L�vQbD�}&֛@��+0�=s޻�Z'����`�ݔ�yW���ڲ͡2n+��
�RY9����0����g@?Y�U����o�Yq��~�U�ND'D�i��?�.�I D����'K5�C��~��?���U�Q@ԉ0+dȻ '���/���I4t����a������U!�+��c_d"$5��-7D�
8d�%�\�J� ��_Z������E/��(�8��J�w)ōq��~z��� sd��w4��(9ؠXT�=�zm��1~e��^5�33aP�
����64� W5L�����}8��I��'s��dz�?��X�E��J�����0�P'2�up$p���i��=���T��Q��m�|g�,O{��{�Y*��D �Y��+B;A�ӏc{H�#'A��@���.�X��8�:��\x�C=Pf�0�X����'ft #��hA3=��A�ԅH���K9X1&��>�7�=sӝ����:�D��:�`&�L� lg�q^h.!q��yc^����:���@�W;UΩ�=�sW���i���4�J��`�# ��FYuG	���jK!���%��H�89��t��?�D(4a��ɽH�r Ic�A��"q�7�0��O1�Z] ~p ��5���qki�b|}���{�?�\n���rt�o���]����	�lR�+���T��t�cA�xg��:m��~
ĭ1F�<w�?׿�T��tԋ�W5�}4��� Q��<%QF�[�&�����@��5���N�?v0��C.J?ͤc��N�%�L��]���s q8E��/%R��.�L��z�p���x~�bV�|�����R��
^Ο�׵�����"?'c]�"��EzM{ߥk�g�����X9=�\�]|�)��j����whk�Wb9a����w�C��_|��T�Hli��L��WC|:=2���*�v���u�ϣ��r9��LL>"�٘�u�W�*�M�r!���K�.�l(-�3#���}���S�$f��$������枸�?��uaw�9R6Az��\/�[c7��=��K|��C�z�{F�l�����SR�)C$�qBz��*H��X���ڊ���p�y.-:f��}oul^�N�Rټo���N���V��!��Vd.�ު�r�I���I�'�?<?�L�
�'��$f�:��}������)���}AIhi'�D���{�JSC �z^D�����8v���H��L�W]v�0��4v;	�piӄ�1o�| F��H(}kB���@�G6P�����}����7+�Z�	������3��i�6�N���3K��f�5�,�_���N{܃y?̰ir�{Wb�s�>���08QJ�[U�P(�w�ا|���5��`�V�o�?�z�`sR9꠴3W?Hi�8��H6Z�|�oU`��;��{?����Gh�p+:Q����l��z~�������3U�BB�zbK��h+K��.ɞzG��UA��� 6��}�\���+�Q���5@B����pL���<+]�W�7y�ٹ���2�L��S����]�s���u���E�Q��;]��PHKT)r���e�h��a��OֿF��!<�����l�a(H�\Z,c�*�x����9�a�tߘi{�.�9N�\�O�.��891
?��u=�Q=8��|*vH]�Ix* ˪1�o Cg�׉��v]��M���T�|}Є�
}�aho����`i�����nRX�
Ʌ2�����
EB�pZ�'7w�Am3��)҄�m�D�������iY7�.
#gd[e��D��li��ѷ{��,�rk�}OH���I&yxx�QJ�Ќ��%��F���P��ݛP�J�]�W��^�a�y��b�������о����FX�R��YU�����s*�~�H�26ښ��2�@;I(�p���\�?����Jy���g�N�=P�Bꙧ���Az�A�d��_m��]1�����Ի_w��[`*!YdP`��J� d�r����DA�gYӚ�>}�c�G�R�� �+����Jb�8���/'lK�mcʢ�Fv�_ؽq�L:f��5�������+�ʣ}��J�a�BJӖ��ZΖ�L�i� ���|�����Iu��@�|ۆY�+{ k��ަ[}���W�h`���^�Э��"��eԏ��K\��f>�<����k6t����7c>�N�SN���^9%5�[_�Y��xu�	'<�#M��zY3蔮S�)��+�vF�>�H�2S[H?:�N��Tך%��	J��_q���^+<�H"H���1k���.�N��T�=S3��'�t��h��m7Y�ŵ�W��X̦�L������)��Œ�C ޏ�B։@z�~0j�2��	�b�xA����1Чz���:Wg�~�:P���*nm�H��A�P?�z�-ԩ z�"�ߍ���O�r��kY�Խ���7.�	i�(�����hp��*����aH )�U 6I�cg�+a����.s�Y�~YF�s����I]�a!Ԉ��g�K�=M����HX��(�[�[A���,/�����D���R4)d��s��O�(�Yf�W��7�MQ�ԥQ*Ƶ��O7�\��hg����D��o-;]G�[+_uN���9���:3T�zd�ЦG�����௽��a�yWY
nTϪ��}To%�݌0FD�%>1!�b�%�n
Q�V[#D����i6<[1�:\S����Z`�i;�EY\���P���S3�7`��Ps�M��̫ԗtM�z���TX<�k��ٽ�K���`�����Xq'���׾��D��ǣ�u�0����F�=�G��~�����#�cƓx���u���ӫ���:]
k���!��H����"�2���Ƚ亙/��}`���CZ A��q|(0������	U:U�0.��}20lZV�AD��h��U�t���p%��s����F�j]���r%��W��]U��B��C�~�K���Ҏ�ю�ɑ���&3� ��tD���̪N���\�iH��k��;��¿���&��>�s��3�[�EOi@v�����; ����.�y��";*�,�YW�����r��3B�D�|��9���������aPA�je�uR�p���9:�Y8�%ll��O��3��X�K�w�3��J?<��_�'S��6�e'���KJ�'�+6#^�6��k���/l?�3+MQ@�V�P��'���%H_v�y(J��f ~���tZ�����1�E��a�����G:jgzYB���� \:Z��"��ǎ+�M�ǻq��J.(�^��{�v_��y:�޽��t(<�gY����'B�����o\�]�7
�S�#��ԉ�rpT�� ����G���<�����[��35(Qg	����<TߨL�M��L��p �SKhڗr������E�B��&⢪O0��vA~��q=/��*b5�<O�"�L���2�v
�z`u�-���Z�M�"��-!O�6KfTt�u%&�퉳�xhN�7j��~{}�r��RR��aPS�� ��]+��R�q��_Nk����;R*�<W��X5�����8�P{ �3_��B*G���zJ>���}*��i�39���vȈ��V)ܧ�)�^_8A|ا�xͱ�ĬDl�$��6ւ�ĥ�\��ǲ��k_��H��OQ�(�$p�{Q���VW+�$ZEi�o��}9v`[��X�e��<�%�������إ��sȰ�����3O�+��_8���j�Y���fS�]�&تu��pP���-©�\a%v�a�� ��1(uXegZw݇�G7A2���"�-z�q�$^���exm����y	��`��ֱR�l-���>�T}��is$��<7����6�	NX�>@gd~�,�WT���2FXX:�/!2�W�Mi����r�8F$�
��ؔt���:4D��F������*��Rv����ޥ���4�
KY.���]P�@Y;����T�{#%��Q�5�Gtף��#�`}�ַ�!$_�"DuA1���9��®�gF�c�3단�[�B+���Q8��Ƨ`<B3�됹�΀���P���Ӝ�����I��X ��7�6�@�`t��G���n��Y��ӈ��]��i�o�H5�NnA���f;����e�u�/�6�m�|<�v��
��Z?���~��#mO?�I���]��?y���I�M'W0IdO*�S8�����Y=?x��tcջ���0�	MIh:vi�b]�p��vs��<�[y��K�g����x���Z�eD翑1V+�c��������8C�����Gh@�v'����J٠-�G";x��9����>���޵�Ԭ�6�]{>�w�ݯ��dr�r��4�qv��>?	��Zi�~���\�M����`�"�Ib���u�l#��$��<~�VSyUkQ:����>�����m�EK��ۡx��	o�w.��u
��~_�����ϯ1O(MƴQyg����G�f��+#������P�L�ݕ�U"�j-��E"!��^������U
'��R�Ⅸdɥ@�3D=f������񓒆<�5Jf�(Oi��pɺm��PΧ��;���ԇWo���Wu"B�������B��Љ癊v��qL��\>0��Z<9��G�|Ĉ<5K�sS�P�
���+��|p��.I�1��J{u�_m�Z���z׳*q�y���l�c�2����Ҡ:���k��)w-�<�kB��X���+�Y�߬�d�s��i�`�����M�D� �D����:m��Y=�����5��(M�*_�0I&��S�G�؏j���$�hI�"� Dg�NS�0Lb*�x\F�~�~��o �*N�Q�6��|e��צ��j�r���䕠N���W3������K~-K���{�~����5D�zP��3޸�*���9�_���S-%0�LZ��3	���ek[�*��X �q���E3�
>H.� RW���Ԗ�3 7^Z���Q쏢ؑh�m�F�F��c�x�x�U����E<�QV ���7�MA=[qgP'~?��OF��l�=-'Z�!ċ��.�ٹ��rG�L'�J���C�����22Vj�I�*�4�v28Ms�z1���h|�'�%�o��@P���̣�p�(1v4�y�$��u1N<"��h������]P;� ���y
H?�Ig�%jƚ��V���J�EY�eG�k	ʥq]Q�CY-��a�G��^.�hu�>E�*�� ׿���L(����ӵ�pB.��ej��dr��ݭZ�|�=,A��	�x�z�Ԯ�ɣm��E��+�J���q;������n���iJ|5*�\<�~@���%����J϶�qC3���	��]�T�����{b�z1�HN��(��;���}$�"�B���"ͦ!sD�M˓�\�=� 6�#*7������F�s. ���G�)�t�%d{t��^QC?����cY��r�Y��V��H�'�T>t������ܲ���쭍T��m����7I�ψ�Y��FH��!$p�F�������H�BJȼ�@����xH���nL]�Hc[CκGYp�i���N�<���/����b(Ȧ�ǐ�OG����)�թe\ѐ����%Z}S��Z,�`�K(:��vi�ݰ�j*F�Q�[�)kj���'������}��F�c�O<
AW�q��%�;,V�|���� �я|��?T�.� c(���H+�.ĻD��+d΋11�ѥ��w�̕I�y��5��32kC���g���iqfY�o�;m�Q�X|���z��=�V�D��k<�c�<Nњ��.ȃ@j��j@Ԇ�-�qj^�~=^��ˣ�6��3��g�<ܝ�*��߈��1�*�p��q�-�o��C������":T� �z�r�]*��k�>�F{Hč�2>>�¿YInAtL�a�w��pR_�7�E�tvl�A|�H<M�sA���˗���r�g�(��X����	s�	�)��H��HZ�1D1b���3i�#N><c�����r��p���d�>��V��8o��A��8=�++vu߁��9����rϘ-��N��'w.��ԝ���t��LT׋Zmu�pk�S���jX�&�Q��8��^eo)m��4�n?�m���>Ci���W�ҧ��3��82�%j?�`�r>^M�t�s|��a��J�Oe`U�_$l�qF�6Lצ��D�l���x�E'o�h@��)k8-��[��aA5��	@�W�� �5�8L�BWe�!M��rE�c��b���~�f��m$��4�y,LңôQ��/�o��fp�"�F��V�:��������@Nמ���	9�
�k��߭�`�h�_K3���}5�?Ɓ���ϙaW���q�cХ�G�ၖ++B@�ꊀl�a�| ���nD��K�ō6���d����N��Vʯ�#��v�꭯9�� �!��{����V!Y����C@ Sd�cFh�U�b���o�2��~�{��,��L�.#�`v,�z
��[�Aܭ�l�T�4q*(����FW��B�/(\���aw?+��)I���btn0�sY4[ۓ�(���� ��ko䉀���vhPB	?���O���`W5����AăT��Lw)���n���T�d�� �z��s���E6t`�_t`BT�
5݉���K!���ڬ� "�	�X�'�(�uҦ�*sN���������7´��
S����аupE����T�� ����R�A���oMEik���vS�o#p�3]J�ǐ�\���g����C��e��ؠ:6�L��Ý�|w�zYS���n<��4�0�CF�J@������R�-V�,�{�F�����d�VZ��hJ�]E��2�(�c
*�Z�`�w��� JSң�&�z�vd�V�@j,����ʅ�X���#.hP#^_��]M���`�5���!�楾<}MDWs��UbE"�0Ӱvt�iO��@z��`ryK���,�?>�C�v��+��� ��a���=x:.s�c��6���N����<���D�aM}~�Z1���D`���0<
�΄k�.���B 4w��?�$LA�5`6�a|��UCƾ���,�?�:M�]����r��0 �����|��naUFOЛ�o�a� �Z� ������y6{��`w-�x�u�f�����)k� �HC���	b��3p�-����<��C�3dD�[wqic\�Dzr�ԍ3$	{�`��nP�}����?x��]EA~�u��{x�N��K��s����J0�s_)��o0�&GE�[�����=�T�2��>��!����EVz��Z)�7�m�T���	]�H�T$gs2t����v��z2�N2ʐ7�3}�!݆$�>��n�D���;�]�_��Y\�>A��1�DdM�-{+�Q(F�&g?��,l����F1Ij4�p�Iv�M7�
zK���Q.�t��?*�f�"�EC'jŌp0t���d�`��_��L���<E~�>��x�@�@�݀XG�.`�5�N{�gDi^	��P��F�'���`wJ���&�)}g��b�ǹ�Y�Fq���ԙB�A�L��z���aQ��]u:`ڬY]ȥp��^k��@���u���R:Con7� ':R��*�&��B�_UI�l�ﻞ�<^˭vH<�|������b���a�!��]�xW�� pv�%���ì�moŀc䎒)��՟��1�_{3��c-�.K.߃XW� C��Z�Z�&&)O���?�"[�m}��w���ܨyV���t%��S���u��!eA�V��o\�H�R�P�+��ߥ�c섃����{��u��7*���nE=G�^���U!��z��;�QЯ��r�Х�N
�b��^K�E�w���|Қp����[���c~���߂����=U�S�KG���N��	�!�Ϲ���(���dr����K���a�C6v��������KՕ���9-Q�U��9��R�IԶ'>(A�ͫ�,v�� h�P���++E����%�HT8��;���f�wv&��_�#jrx_�����ϋ�x���a�]�'*�{��:o�} �V{'��=�8���t��eo��o�tF��a!*��+��Azz|r�(_B5X^$O�b|��g$u18��i|�\�(q�1�1��1򸃬�Q������d)$VT����5�G�b4}�Ȝ�s]��$ʻ���«�<1ߩT���E*wa^���Gz��%�83��g�up!Q{۵{?<r�2�f,D�B�H�Zx7̚I����Ay�w���Q�Tgd-%̏����]�Q��Ħg|��G7s�!$�5M�/�[�t���)T��Ao����ӧ,�`�z��!R�0	Db¼�������GV�!E*̲1�JqZ�����z���D쥵�\�A�XaA��*�>�^YHqfc�`����>+��C�y+��[ǧ�Gk�K0xn��S�
u�6l,� ��B�ry��蜅+���'��e����1QWp���<ܝ��ix���M�l�F<��2��w���4bn|��<�Wq�p�{�_�����/f��
�U]4p	Ƞ���d�3�D����֟�^��yd�fv�B��(C1[�L|��"��C����_�JmR��ɦhO�����%���+�-�3�C�"#��o����?ML�;'���}�F�ׅ7�l�����`X�	M_�/*6�<��*��̎7_ n@���FҐ۝�<��6�U »��j�<"H`��_����0{����ٸC�2g��ߞ Ip��a2�laq�&��tR�qei5'����1�|koK��1U�4�ǂ,�6˭(��m7ӷD�7��{iTMg��A����<B;[\#KP��B��ъ�چ� s'�hO%۳��z�A@��g �Us�zz)l� �	q�AA z\�d�PCC<��3��d=�������C���Ǹ����y���8����t������`��l��Q����� ��S�k��B��M���7���ʣ���jK?E ~s2��1 ��s�P@Up�5�8Q}�6���k��e�y�����{�m���f�?R.��h�q��8����-n��jZ�HP���8�������=��������W��!���o�= E(������&�;d2�H#zgSCG��S1�L�B�d�9�M�� ܰ!Q�l��t/_sBC���x�|�
�N1ˇ ��D	��ˇ����������&`[ܻ*~�Z���S��T��	O�p_o�TSI	��\d
2�,�p�$�A�'l'B�?~k��焼K�]�sЯQQz>�N)	~���h�L�$�[����F\�4{ml�����o{���FN���i��f��ǐ�gin�s�'��O��?�§�-�w�
��� �;5���P*g)Q#��XeP��DeA��T��w�AL�)�L��j�;�Kz���.�Z�|�o%�FIi���<�0��v}��È���bCo4���	;瀞Ϡϭv'�E�b_I�Vj��(���?o�KP�#IdA�������^neM-0 ���O���GAP�9Pf��u������/�g���D_�׭4c��.�\-��'ο �H7�4�Xk�D�@�LqNr�8���|�Vm[��'�[�*c���}�V3�0귩�ծ��3���Q�b�=cd��T�N�\	0��(��Z#�at��E���ɗ.�r��4kw�H)e,!�%��ņ��7���B0��x_R=��b���C`du��A��%���K?���D}f���d�t����66�1��@��e��M����wk�,xX��|�(���hu��'�k_���H�>?%Vkؑέme6���]�YxJ�7W��������y�����]k)^	�4�Ԩ̏��;?.,;� ���!���]e|�U���-S��Q;]���k/�e�Ж�=#¸c�3�@�������	1yU�-°�1C����4�[�zOD����it�9���l���'%��;PPz�|����LѪ�Ia2��e���|��`���;Z�N]�`t�퓌�+>�R�y۳��o̖>p��[�fd�F��a���4�i�l�:���Eyk�nYVI����s/�!�A�Mp;Ȧ��u�e���C�.�w�J�bBh�n`סw1������ۦ�ޖ����o���35����+�U�?��/0��-���t�D�HAk������	?jj3N���.�˞��l'q��H��񔒖��#�G%�%t�S=j�dT�\1+Йh�>�sq4�)��SƇ�m���x*�U@}z��d�q�[�K�l��r\��?���:�],w�H�:���>B�o�a^���@��d<+�P2����Y+�梓B������?�e��-�R%P���#x�/��H\.Mҙ���7wz��s��� s�r��1�)G�s�Ax���,&�'ć�f�kCh㷶iگ��tn�l��';�T_�㢶m�
��Oj%7�mz��H�o�(cl���~UV�����F�dg��m�`�Bߤ�i*�;���[_8\�KS[�>���1�P��������H�q�9��'����.�(�`��q%���W���Ē�^jR@?J��jOE����鶝�B��Vr� �b -r���rq���g�B[�����둰U�`��0�|�v�45t֚����� ��#���+�1�#�sxg�nꭈ�#��4�}����EĆf���˼tn(J8J����<�b�i���Жpaݒ�~w/���J�lJr��D�<�<�U鈆���p�s_K8�{�+x���6���%4���]��<��Ӎ.rg�4}�_E�?�7���ϼ���2؃���'^��\#��g��I6Բ	XK���і�S*_���1�a܃�<����~��iΆ9_iR��]�M�NXV�P~p�K.q�)��J�������Li�3��q�G�N��]	�e|�%ੴ����J�$͚��[�Lnp1����D�W_﹐��u½ߒV�n������$�˃�"�*j*M�kR�i�Ӛ֟�bf����9����t���]N,HN�d�Sd�*��8N�h|��F�!9#+�.�/�4��
#�C���K�+�X�����&�<l]2�z3���κ��� ;��"s��p�3-�D��N�!����j���`�+4-���3��9$ֹD2Mz_�)�Ȯ�S>���iT�X7���3��)w�k�cq��ž�D�41�8����o�j��+�����b�Z�n_��̎�Ƕ�������T*Zr+��������-o�r$�$�~+�FT�Z7����|ɾz��x}�R/]�u����XUm����O���5٩�+�j� �Ƿ���g`G�'�8�M�+�i)L����6�!��Ȁ��P� }q�t#uf�<����ܔ�* +(~LQ�W��\�mltr`�ԯ'VHN�Y!�>+u-I�<uS+���Kގ��P7��U|�)�nH!�^�j=�����l֚_��|LpԹ$6����dr�wt�"�V�"�0Y�ʉ��J���~���`?	Cܤ�{z�}�����\���uKl�VQ[�?��ӓ��nN�N�������zrD��I���ضT��tݞ3|��9��p������Y�1�)u_*o���$�v�Q��Z�\�5���B�@ ��}C�jjɵ�q���y@�|��n�7���m�JU����<�5i0�;T<�1Pl�R��+sg|���d��!�E��ǘd������2d*����DHJ�1_����	��L#����d_Ѧ&�-`_�rV	[ƛvvc�[4}k�0�Ί��s�Z�e��_h�xw��]y������������gꪯ�����]����P��oҴ��H�`�DW�Ih���T�B�s�S�y�����%�����A����] ��
��hd-�`�V���Ƚ%�׻�$.W7������{M6('%�O��;f�t���.�2K�bq��Ll�n��}�}��N F((��kw,;���(�N��!^�����ի���m�[H�����~��q��I9��p֣5��2�&���t��t�_!�ܺC�����9���BE �J�/��ђƊ��.��iw4�vxÄne��)�7�>@�ڿ��l'�T������>�Bd#I�%õ�M�`�h��Hw��r<ꋰF]��A� w��轓9p�h�4}�>�L�Z��������;�H�M�u��a�ɳDOr���Wq�F@��?�q;�gaX���a���qQp�}D�8�G�uN2%�q�Y�>�~� �bx��?z]o�����@L�Al��Q}r��v%������v��j��I��&�s�Et�������?<���z:a�9��4�J\�oGU&��e��?K���4���oL�	��|���_��m�������1������4y��vځ������sU�l��{.�Nr��C ����l_�E�xHO��g���>��(a���Q`�	蒥J#
��2��9��!D�7@�g�Ӫ���Q��÷�9J�#�g����n�CX{R��y�r�uS��n�K�b�]}!��
w��Z�w��R.�7ٗ{P�-y�DXE(��w���Ŀ�J(瑷�����5�۩��V�ROA��z��o�Ρ����`���V$�g��/�XhhuWt2���m�{W'�N7�Z6s�[��S��L�N{ń����8��Y�������N�*�܂���ѷ�zR����1�N(K��,T�����z�
[m�	53*;ӵ�7W#tDI�p(�D�� �uu����ܕ3�qe;�)�M�~�,X������X6�2d(Ō����qy�[v��7��w�'�����I����l�'#�|������>�����=�1��Di��}
�n&9�@_w!�]�j�÷���ۘ�V����_��\�P�˰\�}Nİ�W��/�Y�4���,ڻ�9z(E��	�1b�M�Q��Keuaty>�ɂ~m�j�$��d�@q���ˌ��.0_J?S{����`Wr&E����(�@^����^����j1$����۽�k/H*'�F����ʰ��+��.�`� JA�� `n)�Nм�q���r
��{=�i��Wgi��I��-��M��qC7K�\����4*��@�N���	#�^'R0i����1YI��
�_�\M�R���cSW����Q~Xһ&[�ax޶�r@]��~ّ@���$n�Q���Z��\��q`n���C�����Sΰ#���jlX�C�Q�~���.��qN���a+p	ޤD)� }�Ԫ@�Xv���S_�y�*��|:2�-������FRT�c6S�mF��}��k��_P���f����t����V%�%�H���;�#l���q�4E	�g���;t��P>��L+�Rk������9Fq�����w�
��!��8`I�kq�g`1����h[c4��ZP��#�Yy��҉�\�����7�Q�J��*�t;7�(}$Ջ@۲��xy������C8�?9p�^���ܵ'{�m$������&��Lp]�Q=�������By9��xå�^���;�[��zZ��ں��y�h�~;���J$Y����
tHV���MQ��ߌ���e#0�&`��#�'�1$��Ā6t"G��AJqO�]a>�F/i���H�)�mz}G��
�2��ȣ����11�H�F�(숯s�����}>L�|��`y��< ��~y(�gъ������?�m(��D��Ӫ.��Sc�t�{��4�Z��������P�nˌ"	'���8{��+?�1�����M[%�������csC����=+����9�$����H��Z|���Y�w�����vy���̡j'���5U�oy�L4��آ4�z(�s�1������FϏ&4	W��2('_D���T�ji{)�Ny�����>-Ϳᦍ��C�0���tm�An����(Z0�}��IIw%��!HK"pF����S�iy����	Q�S�����tD�{�)-T�`�tDUz����vV,���:���p�Q�����b�[��u}��'mY2U���F�[�c�Y�<k��&��%Pظ��t&�Xz��4_f����-��ڬ�����aL}�v�;v}��?��R5���Y	S���,j	����n�W�m
��p��1 ��؁*Rv��T���׽��}o;��&&�`��a�w���u<c-w
�Z�C�*���5���."��멹�;0%�İ4�~������!�M^17������ٯ��3n�Ur�rar����.���<h������k���
nǹ�3�h��p�IE,Ő�t�x[�vd2����܇��Cm��a���T S��G����i�n�yr��G�m,�ߟ>>"��Ə���mޝ_���O�Q'�wEJ�}�nrp=[d�ٟ��YFUI<�
����=f�E���P)mͲf���qN����~x3�}E�~��5׎n�m�}S��E�\���ֆ�b��- ���R�oo?d���JE9��;L�4濢�8WD0���;ڏ�1�*�����e���>j�A����n�fTU���V/w#@p[��B�\���_��3��	#�VMS��3;	N<�%�~������gIT��0A�h��UD���6����Fpf�uJ�\U��緩��� j����П� ����g6�s���4M7=(l���h^����tW}zd(0��M�J(�酿�[���*��d���Xۅ�8��1#+?v��tf@���݌M�ٳ|�Ro,�v�ǺuLbĕ���_���4�����
C��~���T���|f�_�L�wF�r��~��j�Z&�t��TU�S\��� �?���-�:6�+�H�����!�5��r����N�H��Ɩ�AҏQW��E�@�r�`��M+�fG�b�۶\��S�i���W���L���ծ��`��&kd�Ӝ'����̸x���D'���6�<tS�� ���>ɪS�!�W��?��Ç�Ԓ*eu�a�'i�E  �Υ�� ^�
\e���n�2i���nr�����N� _�����#`�Ck(Ё��QT|J���<8_��[�}3���M�xZǜ^���x'���D�����o�.ܿV>��KvGR�#�ñ�37�M��v.�H-��3:u��|�!�����Ҫ��	(~e�n<��Mx�����)4`Q(
)����Nȡ�o7X�$@Ŕ�����q���~�S>t��5���1�w�����<���5�K��џ�`�����]���H�h��r=ҕu�KEXa���۵��X�6q�4�d-r��L�sL��ly`b�Xh%��)�4&5��b��[� 쟊�dƮXM�$��C�[��SJ08Aߙ��'���d�^��;\.ȑ.�=� ߓ��� �ĕ�Z&���v�.��_h�q���6 I�C�s	��$��R{���}�<�M+N�n�Ύ��T���D��g���w���#�>NDm��)��*��B����rt����t!�������$�MI Cx��F�s��}Ɗ�`~��R >tAi����)�t��H�s�D�zA���\����F�v�$����'vJg����	�)} �*�T�����d~Bv�k��j��r�a6}X�vOd�螩n8t\��%Bx^�ߴ>�L�C9P�j5@��>"�aA�5�M���'����L0 �e+3�A+�	�N[yؘ\;�pv���K���n4LS�p>�o����(}9�9��<f��j�s����-F�e�D0�Z�4)t�L����*�?�]} ��=�.q�\0o7P��%�����W別�:����ʫ��3��!s��|���J�Xd8j��c;,��;�����N���>w�m����?�Ar�1�t�:���D4�I#"wR?$3�1��&�`�k��B�]���S��= �/7�K����0� � �Q�M���i|s�w�A�2��v:Բ��VRq�&,Pn�X�,������#�X�C�(���LN�:83�O9J8�%zz.eb@��w����<} <~���͇�����7�%���{9������ϪheF�l�9l�8`��V�s��/T��;��!V&�6e�8�P	�W(R��w?��s�2}8���-�N�
N�$�T�ar��������/�ւy��5�#�V���8�iS堽)���aW����c]�`��N��*�Mp�ڽ��ss��b0�+3�::���jq��PE�	:��Y{��Ix13��	=x&�W,D����{�eg!��*5{�FId)*�T�|��R(��&�qkN5���̤<U�[����~hR�r~�D��X@���<�*���+g��5�)����ܟ�~��L�� ��[W��k������2��9�U�Wr��#��F`��O񷘸�m1�^/����h!��Q�>�D�5�qv��Gڹ�/�J7�!3CMO��#r���,���{$�G�r?���K[W�Q�̱�<���9�<+�q�_/�ѳ��}9�ҽ�NQ�ШBS� ����9�j�&�7��]"��=ao�{מּ��G���T�C>���pR�AA����5m֕Y���~��wyjrxy�a�n���/�q<o26���O�A�v"XQ�e���p��,��,�V���P^���y��I��}7{���2q8Z��n\8��b�>FR���p;�Ȯ�@*s%?([��=<�D��M���d�o��1�$�i
���0�������Q�L��ʖ����̂���MȝT�5���r;\��Gq%l�m���g��Oo�	�����z�7dM&��c���騫�||����S;�\�!4��g�D�t����P[	��*#�>���9IF��a	�zb�Ӱ��PT���;z�R=�^9u�G���쯘H88�LfX�� M1��V>@!���]�T�b9�~�v��ou�`w+�"�卡P0�.��ABtk��]�4�5����س6���-7Gz�_�.�C��e��1�Tr@�ud�)�Ѧ�*[�_\ ��)Ж���;�>?uS��~i�eS���Z�nsұ�b����s�7͓*C���y���hI�ZU8��+#���:�(S��gD��y;aI�[?9�1\�*�Uu��-�� �1��e���9�PHE�U��VFh/��╈J}8r+�{����������ʤ(i�%�v��j6��ϣv/���¤�!E|�乃�Eʃƴ<�^Mk��2Ǚ,`��z$�3
*�[���R?����ō���q�_�GS�!��ҳA���$�K�S(EA��Hmɗ����
V	�\�W��.H�����^���Z���tqi��Sr �_�6�V�:_���OJs�