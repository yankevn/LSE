��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2X~�*���O���k�<Ζ�?
J��I���iR��eϴ�J�Ij�Je�V�e��JB^ �9�E�|�h,����� �������c���k�zbr���A�5b���J�f�"UP��"� ^$wW�1�t�Ў��	�/G>�ڇ�[mȺ��j���K�_���)ϕ��4�����k-�mVs/��͆Cw�$U؇�/4dY���J�=������ ��e[M����
㌞c��|?vNqs	U�{)�i?Է���;�Q�-��r����r4�J�k�R�O9~��	����\X�M��^!I�Z׺y��A�R�^)c��=�X ��`�R��YZSO��U��}?�5J�*9;�˱UyT)�4<C�P1��-ʨS��^*���Dl#����󛦵��qD�s��$6Ϩ�@�;��pY&���ǖtm���>���w5*�|
{�P�dKݱܪ:���ń���4����)�\�ޤHy"D���t2�m�I/?{���z�+�� y��h+4�Ў��" ��E~7����-����<�a�ӱ`��kh�I<l�c�w���G����z�Ƃ�>r� �f=u9��p�Vh��2Ã��^C�T
otZ�6k[qŸGhtV�g.�9X�P��Zj��A��5�^Tp���J�k��XLr}�}�w�^i¶P��G>>fˁ=u(��� ]W�2���s6�U����ĝ7�#�5�f��W��G�h��¶[4��#d����Z$�;���<��gNKy�̡�-��,�Z�?�I�߹ʩm{�PQS����c)x�h�߯x��1㺿2R�z�+(s$�ZAo�~�du)d
�c!��6���
#J3�M�u���cϖ�.�|t��=� (e�mVȓ���H�P����	��R���������5F��g:�$亖��w�gUQ�ɠf-E�a����[�10�2J���¹���8pv1��6L��]`r����'3���S�D�U�n�4~QPїVF��Y���T�8 �q���²����������Pm(�?�J�z���R�}��!x�/{�*�lxw0���!^���M5/�&�����/�i��ay�L�����`�s�bi���A��QAd(zބ��N򰽣��M �z�X��c4/;}�?��X��y�)G�)8������`rG���_�ԇ�VH�8�}��]�DUd�ݪ��z�q��#���rs ��={�)���n�q��ښ���V�;#��h�`��xU�T�z�f�a(�����q�B�����E����;��Q�� K)�.�Nqvϯʶ�V;�h
B���`3j`�=h^��jϠ(a�hl�5�,
���GP�[�2��Z�O�����+�a������V��	�>�%��|{"'�1ֱe�!Bó�s�*j��11�xjL9×C_��ڊg �{��Z��鈹P%6�d��b�C�N��F�ȴ��[��_1�Z�?��BH�7��2�V5@��5��0��0 �IWp����*���s�&��yv�c�h'��繊x@3&L�"���,�ʼ��UmA��Z\���짊��5�>�}N�^����Z�����Y_�v�/T�M��}9�"���ՙ�/�bg�	G&�O<�9ΟI{.J��1#n�F��y;Q��5��[��$���i?o�kP���\`z�2���Bn�^|�o�ߦ��vE���-�2Ф�7���Ċs֑x��l�EBv�()Z
��� G�&����4~�+&~�Q�(0��QlqVǇUV��]�	IR:����luaG������P�q��Bߜ�;��36p�o&sJ��#�<�Zt��]�����T�%��K���斓�Oq@����8y}�y� �9�A��˗�*�#P�5�@�t&��.�E不@ׯW�/���Ry3�5A�2�����~j�-?�I^��Ť;��Mnz6�J�V%�Ek��O�Ψ��O,�EO�v��Cr�͸�:�|w���W7�o}�$��譌�Ī4a��ƛ\y�Jc�- �D����T4�n��,,����Q^�}H��N��z�Բ��@��l�b�5ǃ���s���es%U�_�����݀�	�`���C]�`%�p��E-p�:�JE���]�Y�8Ĵ8�蝝��1d��7v:�`K���`ty��	g0=�%7���O]N�Q��#b�R �ye��-_N�
�5}4s�&"��D�(Ie����8$ܟ
�~���aO%��z�=�4R�8�C�uи�Q�7�P�\�G�����j�Ge#��}q��̼bx�#�?>*������ �g�v9�R>���`����I.m)�+��#L"/+ǣ�T��v�E��N��5詴�`�5V�������4���)Kf��<����φD��i��c���!  �(�j/�QT�� �)U8|�=�
��C~�wI����E�ſ�	Ӟ��
v tn�s��C
U,OF��<�BO�`QMbRP(Mޏ �B���kF�9H|?L��a��EH)�+-+\O�B��
�4WP��U]z��lI�s2A��#
�{���ãlI=��k֠���ֆ+� �Y�$�Z,���A?̡�6��jH����Ow�/x���Qկ��"؈ZzH�-���ֹk0(�
c'ݤ��&�<yX�����[A��}�琺��r�In�3H��j��Q��J���[�Q�7J�A��?�Ι�iS��U~�Ԫ��q��N�2����|�Y�~�Le5��b�����*D"seZZ!>4؄�)_��wG`dys4W�r��9��$B���,Ȗ�+��I�*-��}�a����4�^��*�/��1�;���@{Gh����n`����o`��P-)T���r��9[���Y�1m���%tp�Gjw�C�*b�1pB�Or��AAS��7񍂉���O�ό0<������DMj2�:�BW��F�ӗ����&GGM�5,~�����
�(R���"HЧ�(�;	,o:m7��8]���E���*��,��o>�]J�b9�0z���۸����!,�Ū)��X���ήR���b�w�?[��+J�̍� m־�&����K]��$�zǍJp�]��IK�?��6閫T�l䎜���#��� ���&�2C��=���A���n����X��EF�wp��Y��ƽ�氙��=�)!�H�l�Uai������%#ƓB��k���i�i(�\�̂���UX�E�9Y�z���j���>�0�����3���0C�d��GCˉc9d�����#N&���+��	��Nͯu/'^`=��U�m�h�x|<"mеI�߱0nAQ����ߚ��r�Z��](��сN.�c-^��M�*)�@�B�HT0o O�p|�W����`ӔT/���&f��e��+��]��%�"�e�UQ��6�k���E�=��M��ꭜ�����n��-@-����өL���Tspͤͧ�4[^x���;t���Dl*�n�`nJ�%֨������x& �]���h�����X��E_
�E��MFOʺQIG@�h��ޠ�#[�-������0���Rk�4c܎��7���ks^�ͽ���<k����0�0@t'Ov4�@4,f�ux� `%�y�J�S��\������Շ�z' �"����:���7Ch.K�mĴJX�o��&�����Sg �l�*���SN�T3�՗#X�!�>p��i� vI-M�Kk�kf)���\e-��?����9}���� z�(eܱ�m��㐘��V��A�d�o`�;��֗�P�>�D����Ǵ�?�vI��I�t��"GA��e ��#��<0>�2�v-�d	4%��d%ȱm�+f��2AK2d�
�@!��zK��ړ֩�[͈CN4�HH��D�ƛZf��*�O��r.�Q�E�_�__�s0�r�\tZ�My�OjuKa��X���/G�\c6)���YpOVpDxۀ3"��� ���Gy����^����f\�2A��J��:,����� #�LwT�_�?��M�ɜA���-�r��"T�[��?�(���8�����1�:��Z�>�~��_:r���~��8����0�Cmm.�.$����J�p�A����Z%�#̧C@�鏓�m�\��8J�'�"p��S��{�|����Ƨ����ƕLd�_n~�B�_&�WƆ�ak�lj<���+��G�󚢄J���?����s�MuG�KxNN�X��Ƞ�D�(��5����g��`"��1���i20�ppt�"�_��n�Z?nS�����Eɲ�5�	��<�ـ�h哔U���=���+M,5ip��򷇗��]�C��_���y7	'���1ƌC��q���:8ub`B� ��d �����1:��T��O���f^���ƻ|���� *���8
�[��ћTϚ�O�O��Šڬ���S܅9�߮`ʀd����A���f�]`�6KT��:>�M���$�~H�F}!�〢����0�^��O�����I#����B4�jwᙡ�ה��g��O(�08�J6Z������X���\!����1��uEI��ޗ���!�0kL@��c�?̝2���^�|ϕ`��F�Q.R�(�w���W<��� t�S�H>���@�+Z��Qm���[�^��������}�. ��[w�� �(��RJ¢QY��"+{v����lZ*��z9յ��N!�#Ѹѣ��+3�|���qqӔtړ�z[��C�&�Z���G����SG)���l�2@�OhJ��z�Q��[W������-3���=& I�s��m2h}$�3��ۋ84�b������VBmk��g�5�^oI(51KO �ږ�[�;T �a.|B�����_E�����H�`�oe���g�����|/fҤ_슐�7N��U  �*�
��/"٩q�&�ӭ���9fB�WH<��L�6���Q���Eq�E�ǊL�o7c:aF�	�h� ���('�XHUP����O������G7���#��[��Of� C`�3눃��"�?�G���]?������t��9#�@�$ɽf����뗊^mX��t��`���3��f��å`�|���IC���Ke@ �g=,:|]�����]��p�@��m�C$B��'v1�F{LJ�.��)��zD���9�}�
Ş{yZ���w�9��tt�C���c��}����Hv��2��t|Ymq��#H���Y���4���Fߨ���l��@w;�:�_��t0���k5H�%�{�UQ��-e']d�}m� �D�Dw����]��%���'�F��c�����d��I�;Y(�9���Z�
�A�h��r�b�`�Z��]�Nq��`�.����s5.��#�PA$cW���4N9��so[�B{�m����BB�=��]wv��B��/:�Mᜟ3��;N�^[��2�sGo��'D��3X�/WDR^�Y��ܽ²��v���౟��s��\f\���f�lK	L�G�Q��&}�l�����=��B�D<L)�gP�@�0�{c���	xd��g�#����<D�+3A�����w�H{Z���)�v���~s*���<5��w���W�� �ab�1ژ}Qц~h��p���+GT/�ݫ;���[7��\��Q2���˔��o�#o��uI�Œ��Ǫ��s>�V��w���J���b������A �nWF�ߑH׳��O�`�w�iM&B��	y���@�P���,����%�����3��g��Wf�+�5x�,-����*���b�k����oɴm'CNޤ I�'��߇7f�9=SI'"��Y(nc�l+2��wAٚ����6�`��~!,�ٲ�]�������+� K�3OÝ#3KX칼�o���]_#�:��ލ��\�W���ܷ�(��e���j�t�h�w�U��}9Rg���i��ʇD�+�4��CEHW�%tf�V&Z��@}�}!��ұ`D#�bc�G��F&���]�}ӿ���ж׍���������ϻ"y+D�Ӏ�2g�^�Ⱦ����D��9I��6pR�?~�6M��0/1֓������^�LA���tZq0#�|!��#��-4�:0�͑c���h�S�C#��S��"���W��?��9�8�\��v��%��WWU�H����9 ��:�>�&�'ٙ��;����\�B���{�[/,X�����<(K�mm����~]�VWBp�!�"�i}Z���kVs?y ` Y��I�Ŵ��Xl�&^� C�s���O�e0*���Aק���I��{J0y��J�:�Ԍ�FWX�/P<?����e���ӱ��g[%��<�w��C�vT����8H[o�+�Ƴ�>�e��������n}Vf[��8�~7B��<���N��^+��Y&�:O/�L�i����@]�JE,2�\X|�x�f��H́����`	���0tX[c#� �f�����Lz�� =y�5��I�]՞��.d�:������zƭ@�|��)���(FE�L]���\�J�~X3h�P�fz��_����(��0��en��+�F&���}��r8=����h�w<)��J�N���E��SuM���gJh�����iK7�o��
��8G~�S�
�oU'�5�����x�Sy�)J#�\\��H�Й�	�XY>��8a;r�2BP�����R$K2�~]UTdЦ1��b��L7Do��f��X��ԷZn�@τd�@U%�)Q|Tb=��R�j�Sx�i���r5��:����&Z��

<h�<�~WO6���9�5 �F�x�e[^�ŀ��3�tp���g����<cL��YU�A�k��Aə�.�K�?/�*ҝ��rh����D�o�R�>�.�	�
��p����{��/$���g0�s��Բ��2w�α@MV���4�a���q�	��$XM8�B]i�#�	?;�7  �U� ��2�0��d������ gtgY������I�FR�{�ʯ��'<�	��l�HcV$t�DIWo�v���{�Pw��?MF\0M�\r��d���H':����(:��lQ���Qz��3�GlY����3]�U�YNk�����L����:�	�J�h�'�*��pf-;��ɳ����jD&ō�!��������O�558�$�3�t����Ȁo�ߩQ��IUu�|
��|�w�����4�@L��+�*2@q����\�5�2�<[�������$Oå�n��s�
��+87��#�"@SM�O���Z$��;> 1H��ծy��#�?���g[����at��uܷ+C9o�i���kezAV=��K@//��w����)��Y���z[Ɖ8XѐR3SMߐ��������CC��+D��QN��U�ݫV,@"VR0[Ⱥ���������Y����Ŀ�j<�� �X�G���;�-z���|��d～�X�R}6n��N�����I��R��q���l$t�CIn�%lcۆ�m>Ć} 1�"N\k�K���Tއ�Tlt�ߝ�[29|�BP��`�/��/��u�|>�H
c��� �Ȕ����}�^q�_��b�H��+�*OG2�a����&���&�Y�Z�FNna0mv7g�6��V��ڊ�Pʟ���$Ww5�P�2&�e��Ìe����k�����S�@�%i�2���=����'4�^N����#Y���!u<��$�(���v5���SeV�bPO�V~����G�$��t���e�9�)�#���2ԵY_�;�eab�� ��G��G�����@��0SN��3�}"޿����x��D.��_��f��������n?[��4���q[ZX~f$��*5y*w}$&�� G[������re:z�FB%g�����Gֹ�!�Lǐ�%�����r�� _���o��#�Q����I1� ,����I�&�5G�f-�.�=���n�l�sg�i��������x�
����k	��MM��v�s�:<�^�X����	�\�o�]#��7�����F��g^;�Q��j��XVL��E�:��gªM\.��ln5��Q�i��m���	}���m�;��u��{.x�d�j�7�g�׃���
R䎷h2�(S@6Ft��E��q��li��.����d5?���#����0?0�mx��R�ϑ���|��,�l�]^�V�U@&	MHj�&�B8(�r>�g}]aiF�G�:�P�eW�H3��o\��gL���J�S��n��?����9�7��_������Ǟ��8���DsB�E�]��2xS:��F�Ι����Ro�Rꩽ?�9����� ��i�(�!V	5�EZժ�h$�X��t݁^ ۳ճ׵����M� 6�Y�txS��{mDʙ6���9�,U����>o��٢�j��϶2�"j���n��r��Z�J��f�#��C�'�!j2g6
'�6��Oق��z���}������eΦ�}���#�a���r�MR)N�o�*�Aw�-ؽ���	�,}��FsA�C�F{;v�?�B�Ϳ�|�-��Aɪ�TM�d��
Z�J��=(;���*����
�	jp4^�����`I:���r"GCؒ;�˾��������nA�Ԏǒ7��u]�q�87?�T0n��h�{�U��/�k�hHrX���~aD�����~�t=��83�$�f6!��&�s6���t[2�A�đ<#�у�H�M�s��8MK�txv%�KC��-R�t{Ƴ~`�$(�����0t���JP�_�R7��B��Sݠ�a�>��@%QJ�.�޹3�J�@�e��9�w��FO��x��6�T���	�4&��'+)�)}��_F���$T<�
�\�
8Ӧ��X�Q�n͠i/ì��F������
��oTI5�$���P�����ET#0MN��:��	�k����s���W�p��`����L���!�&���1�+\�F�i�;nN-��Aq�Bd�e��D�2�5y�K�h���a7r0G��F%����C�X�d ���p��E���8��5���K�߲�]����u�#\��0�;�}i���,�p� 끓�Nrh"@�LO�g�vɬZ�6�g×;��cO�j����V��m��d@#k�Xa����A;�@�z��&��;ШJR=[f��R�^���6c���q_�"h���@r�/.L�V��������4�3����������l��~EL���i�>�Vm@Dg�
�n�Oo��?bk��V�Op?��پȞ�[���g0�AM��4��O��%r�ʀ�"W��E��ɧk�0�!c��n�e�B�R�-�j0�$BU�}{	�8�P@805
����0����s���`*;�dJ�1p/h������|����vC�dr�WN�C��u�34Mnt'V���D^4�������U1��0S��	=v��E��4�Z~\�N���q�J1Wd��K�}�Tr�ُ���t�eu��3GL���a��7l������j��� �W�دT��+`J�t/�I_] �G�$�r3׊����]���H��w~�}��m-��^�
�>�Q6����MFq������m;����ъh�I �:[C���@����O��֧^��K�hJ�t��ʵ�N����+%���i�A$fN���߂��9đB�Zl��{�* ����kb��j�3��AT�m�s�<Y_��X�#^�~�-d{���e�ݿ����to<#;1gh|��ڭAE>xvCFz�D��Z�>�N��1ּ��X�R9)^\��w9��ި�1�,��Q�m�w�U�1Ad���;ڷ��o#���&_G� �'���a���vdd���.@�N�E�JtBT�x����XH�Og�i������#ȇY�	�"�����u`��5*h|7t����[m9r�uj��}�A�au<���7�i����JP�![2��-�U�L��=���(
W^,��Y!f��:�X�,˒�l�_{��[m vo�LM�a���<"�&mJ�2ļ�j����DQ���K��|��'�J���������XS��|^&���y���_������/�9��ƃ>�%�գmbU]�A�0�5Թ�)ͼM���f7z}�זz��v��F��ر��;�-y���b�w�m���;Ec�v�cAճ����פm9PM�Of�k�0h|���e�B��S�q��������a}��s�,Ga4��.-8p��Xh�6�JRw>���&h�&JdmR��}�_�^�(J٤�@�e{F6��l��,�Q+W�ċ�� ��s�
o�b_
Ҿ�i�$/ ;������ ��8�������CN_�i�{d��5n�����1�Y��Ai�DЭі�b�e��m��z�ل�� �� �c��U[�k��
>i4��0�V�tcvδIR^���oYϗ�����;��oof��V�@������EBO���܁�έ������~ۄ�8yR�A��k��ߴ+��79��\�ðC�p�����Or^�����Ą�~�������aNc�U��7��Qd�rkƯ����j:[���a�W�M�l�M�YW��X��-�:��H��~���vHo���}f�(��+�W�ب�ɴ�P����(�7L%pV���ey=�RE����Ϯ��g֔COb.m��m%F}u�`��L����
C��_;���`O � �jh����?�0S����ҭ�����p��ܧ<�Y�����o��HD䱺9���)"��*Zca����]^�c�쑍��D�jh��sW��aބT��E�����:}����@�܊���'���9�t ]��w�s�X]u�uջ�� #FP����3�%o6��.XC!���cfc��W[�4���I���~�l���U^�=�� <f����^)����M��x-�{�W�����l�fD�x��m���ʁ�i׮��v��KfOhZ@LMk��+=	ey~�R��p	�^����uz�Q�H�[��%�\[���
�U�a��V�F��Ȕ)���9Qq	�?Ŏ��g�<&���ٮ���y��2���[�-���%�?1rg�-�c�NR~"�4K%�M��-�G�?�ߟF�X..�^}���x\�٪�)>(���-���B�ӼW�{���o��uao|��11k�U�ޭ��4GP��]��+8�{�'e��Ma_IlD��䔸���`�v��yIof4~��^�B0.qs�8���	kv1\�z���	8�X��Z������w3��'m4���ǖk̉�Gy���^�� ���
:_
엤%ޣ��߹��T��\S��c��Z pj�)�3�~Ѩt0-�%�=��{�#!mA��Y�P�?���$�D��.U�q���qI�sDȗn�QE9�ԣK����;�g����&7yԐ�9 �� ��т_�Ƹ�e�wFp�<�� 4߮�����T����|Ҭ��*(�s�tˤ[Aǖ��g4l�ٝ$��Z;��$�-$rp���s�G�����@~0��?D��4��^�?���]��x�[L9�*��o�y�*��	ޭC�.T�`�_��O�Vry��a�������ߘ�q�(|��e53W8�k31K�����@k�Bl��h��3��=�2���r��D	���[\�";l0aZ�2�$ S7Ԛ�F ��Zq��k硫������֝���5��� 
ޙxh�cԂrg��ߠ����o:�]�����D�W}DlW���>���*|tL9�$���9�b��'�JPQ�E���7HL��s*�W���aAx.Y���!��G\HK��k�7qXA��`�l_�AU�nA�T⼏��.<�����DM$/NSSYXX�j݀D�lD}�V�P���wJ+�ްؤb� \�-�-�<4z=AS�O"��F�@w�|A���"����9�d
�1h���8���g��ό��������.,%������.�ܺZ��;��9�Q7��y�mc�0��HuV[,6��p���������="��KX��Zi��bh�)�ӓ��}��L�0�6��(�o���6��QIִ�=o@"�[GZ�J	�w�y���:�t'������*�4DQ9�F ���D�g��4�^|~>���� �ʁ:v�����.xw_|��sE&W'����9��ۤx=!���w������jCʠS���'t��G�W��fuA\��e�-9���;a����5���<��*eW�'X��;!UE�Mp�roQ+��DW��_Wb��&�"C�QS7#.6̓Sz�F}��{M���
,�����BU��p7�l���9���9_��Wк��B����G2?"�Z���rd� GG�&+X��,N�b����=��
�������~�s�;E�Ѩ�\�?�̻ �e�%��]�fPɑ\A
,��d�#XK�j�,�� �l͜(N�0˒đ¥�FbYc;�r���6��.��P˂^�*��ƌ?ͣ�_�ݙ7��b���t\~��\E���oM�9k5�����]0c:�v"<�Aq��s�fĉ<��$��X���apM��c�=����5/v��Q�T���.�|U�1&���!"!k��UF[��W���� hL˳��鋭ᕗ��8A������b�����	��AN3�;5��}�봥bX���)+�ۏ6!KL3NOrL�zI�'�!��9�Q��R�5L��圖��D�>�����҃Pg����2k�����#�{G��&�lj]�B�XR���EF��9�s�:�x���4C���4�T���x����̆��?�[}1�C�[���F(�Q��W5���nu��!�����.�Rh;<�$��Z0�YI�c`��z!��:[ܗ�=J/��I��ȷ�4�X��z�z�����Ww-��;�����b�-�{}�m�D�F��}G"�v,�2�ƙ�?�����C�b��J+5T������g�ؓՄ����B�'S�������ޣ�:��5�5(�1��=R���32!Z]��e6��3W	$���+'W$�Jz�8���Z�F�c�ӡ�tk���j��7���tv������y2D����1�G�Hh	�FL�{%Ť��Ӽ�4�f���YI���5��c�=Ø��� o��+�d�er��\T*��t1��Ajf�S7N�G4.r�Z�6���~4pMR��P��h��2����3b���<y8e�z�[��z�ll�+_�<��1�0��M�)j��7j�/%I��1�WC����h��[�CާKM��
y��\�4^���V�sh|��i`I1�β��撼���v��ݺp���}?�٘��V��7&3�� �^��f2k'Bxɔ�S"IЬ��¤�xo�u:F���J�V(/HEU��J��,�?���I��I��������p�Q��HG%N!L4߁����e���c3�jA�w({N)�$�t�0��9Z��d��1��>!_,	��qoɜo���B�!k�G�~�R�Bkv�#*����7��w��t}��P�a��d ��I8P+y�nxĬ�e�^sæ�'T�t�@%_��F�9�w�l�ھ�G3�9�玏�����#�'B�?��aXM1)�����e!2�v�sV�|hӪ���:�~�3�2�' u�.q��jǬ�����y�aO�رN������W��\uX�y�+�y���/ei���`Us<*�X���.�M����w! �G%TpQ�Pf�۱��8=MY�_7�lq5w��P���?�w�8'ݲ�����!��ڃ;�(��i4Ű�(.��� �-�g3��~�5� �鳥��_�������<���+;��>��� [��߅�B,�ď��=�E3=�7ƹ��	�[�3���Ϥ-Q`Μ�1÷�s�=���g�eD�T�+f�]@P�g��!�*����@��i<)���̎��@U�|-"t����{�����!��y$���4���ީJ�*��XV�|w��B���	��*u�K���������Ԍ��&#7�O�����\�WN�{��Ő�ø�n9D�|��+�H�]!�f
�U��r+>��4o����`V��?��ٽ֋���Grr���@� S�L0bk���kВ���y���̛�ӻ56�pwLԱ �5� ��	��ܩN��pW��3�U�H�w�]��}��h�X�/��FޅӀ?����X�k)����9�������H�������M[��9���f$�Ջ?�������Li�V���U�/c���m�ds��5A���3ݯ��n�mNF��d�c�Eh�_e���F�5lPD�0�fy��1
U�;ہ9�)�i��F��ł@�R���mm���;$�����Fqw���-sF,�,?����v��*�ftz�k��}���掇�`N,m��!.-�_�Y��9�� ��������Y �R��7�����/��5��CI�^�7�{���6z���Gm��}�ߟ��d�TΝ:��ʣ���J�"M�L��Ĥ�"ֶ:f'�:q���M�-�fo���X]��}��)���Y��z_�hy~��6�r�S����^)C�&>uHܝ���b��	=�17�V�2��Aȼ��;��&�_�u����,�X�u]-D��c�;OL�N�]��^!���N(C��.rb�K�E��:�`v�\�����B���	��U�h����_����A��,��w�!9p\F��c�y9�	Q�O��܎.�Ж� !e�)�_�vjt�1F��ͻ�VOoAJ�m^�~;��>��8�&�pp�S­����Z�����X�d$kp��t�T��'-y���,vY�Gކ�����G�X ��l��9���ŭQ��W�B)�@�n�A�u�G�ǣ���X��^�9E�k��ȉDS���E�&��7�ʣ�論��*�G����mI�͹|��#�q@s�IA�H�	z�R�#�*72f�Ďf�֢v5b�� �Z�iI�6�!%�I=ؾtR�A��`���E�H��� U��i�ف��n�)�.RS�������c7���6XD���X����Ki�u�������V<B�N��`0�)M �&}��z��k������B��Ҹ�!��f�tx���s�J�o� ˴^�I���[x��H���8^��QL�2A,�%�d-��/d�FA�n��6��^ׁʭ^�S��ZJO���Y�;2��@���?	a*"��7�}����SΘӹélf͌�%��7QJB��=��4L�&Z������yK�2�5y.y�f|9��=�D�$��4!������_8QYl�_V^d�D�R��4�_F�/Ŏ����v�nC���kLn*���ݛU� �����V
�d�iy��v�-,��nD�zF%cZ�=T���Jvr��[uq����R~2�l'�Vj�DЀ�>��V���&�>��-�Y�_*�v8�F*\�q���IkGq�\7^�Au��w���*b��%/��V�'J�ե��ۢ}�Y5#.�u��Prh�����R�E�SY#S���sMAD��$��ߔ�r�k,�2�	BS���AĀH�_����)�s��><��_����b'2��|?���2Wݹ�ev�l��~�K-)}/EA��k��\z�\N���E�kS�URԀ"w_�+�gD�w�F߯Ncd?��w�h[r>8��;\wv2(+Mc���Q��^�j����9f{W�tNb�}�D�<i�b
�0�wPX6�����/���W�� ��q��e-���L�H�4f���I��S�Qi���D��/����)�����7��ltg�U���M�{�B�~U����=k��� ְ��yh 5��ǻ�p���>pɋ#���U�o��^��S9�
d�#Z�2�f�ˑ��~$GB.jB>A��6��ҐId�P�q�u��W���'n��}w��^��t��K�M�hY0���`J5��� ���h��	�vЦ7%��-Ʉ�^�bLI(p�*�0�d_	�A�Z[�\�!3�1�0irZ!+���嗤}�5�w;t��0�.�<���/���!�S�=_0*:W�X\��ns<aL��*'�P�����Ҙ~��m�*hk1F�m�_pg����h���T���q��xo	�+���cT�%���{�S\�:�s�*ea췙 F<��n!��6m�#��$�u�Ύ#�׻&	mִ<̴���"=�h42c""}�,O-��=͂�����T�{p$t����
R+�^.2�F��\�
�E�Ͽ��΋�S��p��N~}9��%tGW�Pe��b�ل��ur�v��F�i�=�w���qT�߾��	�=�t���,!ݐ��y�?�\�s��J�]�8%��!�O�O$+�A:³0|8O�d����V#��&�Q�Vɛ�/hƽ7o��<� �D0��e΍c�3�]Ԛ�+�}p\����ƌ�u����ȓŴ���Wz�3�����S�S	cg#B8��Gb�T��-���R&V�P�E=���)8��Ҹ}Q�����p*�`� pcP�)Fܼ����5��ƔFTQX��/�h���!�f�_�H�n��V�3�6��D@�f�8dH�il@}�7�e��Fܜ//��rK�����^/�ڧ�������E�n�lmO�4p-�P�3Ƅk?��z��ǰ�־�1�ӍFk�h��3�6��z�k���m[�ʛkt� ܖ����5M=/�(�ҵ�@PC��%���ɛ�>4.Z��M6��bˌ>z�>W���u�)x����.c$��牂n��Ԟ-�\��/১��IR��-���q�4��������g�Rr�^�����mu\���y*����p���9p{��� �����v��X�RT��NCR��g�@x�*��t��0�Ҏ<0!�O�b�Gi���}n�ی��K����l�îWE"�'�����'Jγ_��g�d��6l�>�]�.��8���ˀl�\L�i|q��ӓ���9Ⱥ�M*?�8�X����^`��#UOm̞n3N��L�l�<�"���3��gi�����(g޽A�ix)�)+��gxt���%�ѥ�H�(����|oa�Q��l���ycgVW�P��Aurq��x��{�4���j�/76@����WH���dU3�#��'���PN�{���x��&��iCm���W�7ûz�u~����_2��+"��dJ�Ѹ3,#eϤ�*��ekCi��H��;Lڝ���kM�ʍܪVtr��Y̅�ʑ֕Z��6����������Q����u��B���Ņ{���g��Vw�U#�QZ�8�[?�6G0����
X�&IW����<�G+ �_7����usa2�7ؙ;}�\
�3��;3�[g _yl9#~W��&��(�p4ϧ�\T����l
�->8]����01m�C��0�7��7��c�:�[G4�Ǳ�NQ���{���GK;�aa�:<��	�7:]Ĉ_�NN��iȗJ�)�A�6C"�F3	`�/́B�Fb	t��.;�:2��b���ĩ-���d}Tq���)��W��l��ؼR�%�X��&$���7�{��F��{��A0i����A?� غqe ��	p�1�iȦSK��+�z��/�F}-CVVw��]iq��n��+&8�I^���A�Ǳа&>(���p[m�^���P����H�G��3�0���� Ji��?SQVAh�K�ID^�O�۸���p1��8�F���A�c��I��%Q[�9��9�ԃ�e��Y�����%dӃ��>��Duy�匓�s��^%R<������$�������1�������@��� ��B���-��u'[���-��p���[4]���W���ﾾL�v�[;[�ϊj�wc$�|�j�2�6�y����|n�S�����Ǟ:u��.�]�y�����N�L��6n����	�#��1�_KLZ��~���3X�aΝ�	─ �
�@!Gf��pj+RWmkƜ�#�[��rL9�nS�4�DO�*���7�ld�(h��m���9�BD��ᠢ��G6�05p8��իN�_BiIlq,��Yc�����-�9� ��T����$,/x����I�wC��e��%1[�-Ͳ�e�nOQ�� �kD(�G�7NVG����;k���wP��{��Pc3���ݲ��$t`�98�t��x|K�oI��uo��^G�>�b2�d�;mZ�i�q��K/"c嬂A3�J��*?'����i�hCn�mI�����DA����`j�f�9��&X�;�B��]��\ȟ2��N�43���9�nN
����Ik��7�~�-ྥhs�q���pŨZA�Qxh�P�b�S3�Tj���3��O��Y�ϝ���*��YEС;�Jh�D
���V�A�swę��w���8C�pu�r/F��*�yS:.����>�;L2��m������S��CzHH����d�-2y7�q�ǀ��M�6|N��?������~���h)�Ƞ���k K
z�.6>�߃ ���3\<�������s� և�X�l��޹�$� |�]R��&wW? @���i���
7�~�O����S��d��%����Ba���b]���GR�cV��_o�o��n+��^ .�0�y8��x�wO�0a��	�
���4P��Z�0�UOs��i4��*�fӚf�Ӡ|�pāt��n���E�F]�����P�.ߣ>*#�K+���"-qk�:u��ӡ��,el_����t��P���wc��J���o=�6�� #�#F������<����t�-�|&-�V~&�T'����F[��c��sqe�����䪥��mӳN(�>�����DM��۾9:-����7��-��ŋ�>��'�� iX1y�ԫ���U���fJm�+��E�Յw�ױwƑ�0��
�K��U�b���/dC��ң<�җ��7���h\� �>G+f���6%:3�����4�'�������9�P�Ҹ񄟆d^S4+�L���	� �@��[S�<��w��[�wfkӪ9m=_ �h��5���:{��T����%N먺'���RB�ʳ�n�M����A�o�ů+-]�IbQ��B��d��</AD�-7��f$J�1�=������
<��R�T^��W)�Y@���M
=h}3�)������#�x�.o$�ח}pW�_��R�1_���%�7K��g�R��J������������Mh�\[f�lkb�l��E7.Y�y���U�m�o���NoJ��.˵��jV��d��Nmj_�L�>k��E���#��dU���00���#.�F��!4�J�}W������:݊d���\��t�C1� �vh0� ����2��+� u���b���/&�Ɛ]�4'Hh���PS��� �?���x�X�;?�mJ,v@��+(T3�]��:p��!O��Cp�N�)��y�aN9�kH�.�������z��=��g�U̲��蚀�${]��ͥi��M-�%�2R���$E�%/�H�~�9�wr	�c���@�9��������"�U��ӑCʟ��r�����\nWXN8�0��h�cg��CXM��-PQb�Yw���9V��c0�Qv����Q�񏬞˓ԡ*���g\��OA>���v���QL�u
�w��VO^����lӁ)�������!}.��84�8l$ر�?�ָT�6�k����Z� xzhD��6P��)�LMZ�3W���Й���J�����a�̼�rT�/A�Q]�]����hW1r$���~yA?��k��ԗ�zwz�1t7"�Yqw��ˎ���G�Oܽ����=E׭��E�P�T��<������E��̸Y
Xn��/f|.�j�F;z��@�Vr�i�^�=���-vEpۥ�FNd��8��)#p_x�^h��3=
��@��s�I�NyX���<�9���icON�%��2'�E���5�x�v2�ܗcޢfk�-�m|�P�@㛷K��+)���8��#/a������npʒ������+vl�Ô7]���(̺͗�T�14��%f�U�:�s��j4�+{��V�F)*^9��0�����$׋��D;�������1ϴ)N� t\� �TDoh�^�6	��M����7
��~ž�pn�����L¥�'
c�@؟H$���e憼�t�k��5~�}$�ߐ';�2U�>��k?=:I��׎}E���4��:+*���~_��e�v�u��O��I'	�<�\��W�F{w��S*#(�*IK5��:�:.f�2;���Q�J*O
�Ӊ��<��;�g]���H�|��ǅR�m�h����H�Q%�X�B��b�K�/��Z<Xl9x�TÌ����ۈp���"�n�wf�*�%��9�+�~�S����W�:׎Fԭb� �Ȍ"2Vhw�?�Sm'�|r[�Q��,/�h�{,Z�.+䘡lL���\N�?{�t�hi[fH1BeU_~��/`�'�x�KGsf�X'�aa@�v}�%)�^�<�����3��|��$��i�h�"x�2zL�m�jl��.�!��M�8�Ӗk�4$p��nk�����ǣ��k�ՐP�އ�/R�Ы�Jz��7C���Ż���g�����%d��h$@OWQD[\�y$����v���":њW�EL���	=�Y���ɛX���d|�!��n�A�7��9^�܏�g�/jdQԶ���V��횪��������E�v*$U�;7��gp�ܕ�5+����yܮ��0�۬��\���B�e��i�����,U������0���O�w9&�"�1t�qWZ���N�FJ.�.�^s(��țXrv�i��ǋ�2�7��;�L�:f�ljT�c7�|5��ۤ�4��h����U�f3w��~�4!����,7��H��W��I�y9*>�9�w��Kl�-4��_Rh)�pz�!��NC�o��M��
E�
5�o@S�ݹ<�e�.(Q���*�(��L�Qqm����3����c5��聦,Y+�
�`�5��A���e�ᩲ.��}/u���+�M0"+��u�O�����6�����l��W�A�Y�5����Ʉ��Ds��Y�.X�=�x�O=b\>�YM�;_D �F܄'���J+����	��0��"�K �|6`|+k��Ѻmn��Fʪ��z\����yWO������2:�vUM\�e��*��g&���$;+�������&V��,�G[C ~"�r �� �:�t-kU���e<a��V ���x�%t�����?>�UQ�e�=��CDT�B8��2��ۺ���==�}�	j����%� ͦϛ�����D��Eq��D�4��O���k𥦗`��1'BG����AC���� f�0�|	��}�z�|p=��a
Q�FO&��F�Y7�?	3��ݧ޼��oC� m����U�J�c�V�f�YL�B����I?���| �;K�-�w�xdDv�6�C�)�����y_^���͢���J���A_e~��.͵�G�����t��Χ ,��,�.J�&·�JhT�+�T�Mbɼ`S���;�<֐��F{ԽE&�\$���M��Oj=��̓'fr��S)�����=��PKo�@��j�sr�Ɲ��CP���A��fm�h��4oD���ݓY�M:�*�/rk�x�Mb�r�/zK�k����U�X6ʛ�u:��mJN�)w���q��S�BL�)3�|�n_X�����p̖O<�ђ]��Y�\gڳ�m�ռs� s���>�M�8�t�C̠P@����W 37LU�\���{�M:�����y$$���B��1 ��W�q����چv����ԏ��. +%}X��ZL���y<�wg�;j�Ѩgd��fq�!�lc�ǟ�C�^�6]ݍ�zp+WBH�\ x�_�*�K�qz�Y��'����6�WZ�^��$�@0����4قoO�������0BR6�)'Չ�uMz��;���NŸ��_B�'�Ȍh4ְX����!^C�8�A�g�ƷϨm�u�Q�H�F �9H[�'}"��E�qy,�����������G��$��]�?���CD�r�7j��X��1+������Km�$;�4i5s�^K/�{�c�sk�H����R
M��c��Y���*V�
��":
v�2��4��d��c�Z�ֈ���[�H�����{�������/����H������P��k�A����(�
wQ�2CT�HHjW��d���!�)y�_�U�+5���緶�m�Q,�{+�|�ӚR�&X6b�O��ft�E}Ҩ����1���bX\���^E�@�_�}ݗf�{�N)���h,5|ɷ�������f��g��$2=��i�����ӑX���[��V�����X��[~RLG�k�rzs��[����{�	�u4��P+�D�)oMd�xO1�s{���p�����H�gE1���,����Z�iT�w`�d���K����8�A��j������f�N��0���C���ǉE������Ѽ��X���b����y	 ���x9G���sT��T��	Tk-�/���;�r��+�L�壙w��[%��%����ut/��Vxc԰�I�P���_ֈ��B��ʴaj�+�:��sb	g��w&o"w����M.^�P^�4a+�K�^I7��[*��B=�({RhT��uLwD���k�Ά}
���QE��d�"auF�F�w�����=-��|v�m�b�O0�F�}r��B8T% �f�^�G�v]��`��hlKC���Deg�ʻ�3:�I3X"o�L}xq���oDV���W��sU=�a�e��~��L�׽�4��Oӟ�5t����h�b��q^9�$`	�m���TN����S���mpQ��1�*�^�	[�}������T󩉁��/E���ejH�Ԡ����9��U�\H�%�b^�.���j4�U�� ���]�P��d-�[f�%/$|�a��4�Vm�$�B��"T��Qu�<�2�G3��Ŧ��B��Jı7̝P��`1%aAw�~�bcn#�5��M�$���2�5�'��Vt�u��"��3�X�Ǌ���-����y���vЏ�Ė��/V���3i7����`_< =� �`����Ndh�Ɛ`��P��hn�S��m�>�a�IP��K9�Z�'�b��dP����|�Aq��i�d�n��s'y��c}�_i^�,F������x�)�r �N��n�[(��:�[QI�l���^��4�,'�b����z���'M��{�_����u��7_?Q�&�J��oR�O[�z\R_�Ro��4S�E������0�c��b��{���3�k�&��w2�h���k��2�[���~f
�4)�8RL�Cf�I"��h�E�B���B	�%�QZ�{�\=9�-]EWSQ"
h�#�B�T�n/q������a�Y��reoPKLiV�r1�{��S3+�[I�ݦf�{ٰ��\�����5°'��<o���]��%�2��[^K�	Z�s�O�Au�x�_K5�jo.=]����%��aR[�JI.�0�V�?|lmD�/z�|��ྭN$%��'�L�ȼ�\G5g	Ad-p(�קG�,2�:2����1#4�ni���J�']�4h�႓C��{����o�I�r���&���L��-j�e/^Ѿ�T3>]9K섺ӊ�%�R�*�(�l'T,�	isw~�j-.���%p�xy�`Z���5'L��)����N�jU��`a�Q�R^<�s&D'�9��J�yz�Sv��<���3�~N(w�49t@��g�G?��y�B�Bn""W��tg��6(�Y����Q�<���lP�:�����8�Ǯ$@1���Qk���I^��6K��<�<��]1:y~�Ͼ����+����H�D��p36��<�Kڶc�c.���䕟��ML�H�n�(�֘�k���$��d��`#��e���bݕ��EZ/�u�p��	�7�(l<�TT���FZ��Μ^HFȽ:3Ws�ȋ�uQ�����CB$z�ϡ���D�n4��=3�V�n�5�B8�����j�@e8���y�YX`i��I��a1��}�:�����������xX9b��d���h��Zi����.�T�{H��׽�Q���'Ki<�����f����!�^��Rk�1y9�FWz��9,0[�v����E����5=q)��k�����%���գj��r���X7X*<dv��U{��5!����x�����G��DOq-��eʿu.�s�IoK`�IA�b�U�-��n� �r��L��=������u�VX�5�~��w��զ%˫�A�.~cc���pwea6$����i�w?Ph�I3U�*��)��tއ�~e�o����/C}yV<?>�{w,)�5f�r)8��"BIN�u}���K��pW$�A@콓��[���d5�?]�(8��lr����p8nVKM�|�h�����-�-�X]�uJ�:�B��֗쐊Ѭ�+z�Jgw�뀨�Y�����W�'��"*���e�_�P�t�G�Rl>8�:�� �W٭/�΋����f'�� � ��&\0��hg�Ξ͋�»�
��N��(yԹ�(��Ћ��#��0N�-j犩��TD[Ғ�������Z�|L+�M�	E�G�*<�C���l*Z(�Gb�(��Yb���56�/���;Q_�I\�� UO��Z��2���ŖSʂ$%j!&њ���;	$�D~q�l�Q�痍��1H�.�ϫ?cY ]]���U�A*�/:{�\v�&1ON��N�1��0���>���/c��h�TLT��X�NC���O۝�t����X��v}��(&���Cy+,dr��I�M��]�������z����I"�h���c�_��k�@[o����c�mi��̛�G���}O^3���g�;Fe�jfÎ���Ä��*�v�z��U�l��[�������]͎�!��Ux
A���!��0��lC�w��{�������ه($������c�H=w���ڨP0��\6���/������ ��cF!P}���< �sd1�9߇�jF�g1�IV��o�-)�I�RA��U�]�����0�?X�ͭ3�����t˰ !���4�0u5Vx	��U@|��
��{�w�w�}3e�f�GU"�U�鄻�0��w:���l.�c��)6β8d�UP� �4���?��(�x�*��	��U�q��<� �F�RU�N�hp�7�f}���g:�EϘ�a�OuݣEh\��"h��/�@)%Ӎ�i�t<�Nϻ�L;!�0��Y�y6LJ�<赱��H�Ouf,�l(&��kֺ�Ֆ�H�QJMT���w%�a��x�O�J��`Q6�}H&|���i0	�=����Cݦ4�I�ڄ}T��Dcv����:��[?}�D��=@1�U�)��'f�vR>4�y-�}��X��(�J�����k��MB���B����%����9�F�o�jQ���(p��Mv�����79P��50_�R�uc���x�.��|T�%����PM��A��Vˑ���Z'׺|��r�
l$��jc���0�,�����|H���$I(!�˻��1��N���J͏���aV���6F����n��Ԉ�T v��#��70(ϊ;ḿo��� ŦaG%�7�<߫i��3M�i&`V�a\�ت�^I����2ӯ���������K
���A���͑Eq��D=Թ�8ۣ�0
	��T��~&�bTz�1���?�!(;K5�ج���#�eu���ɝM}r�gv�AZj-@�	ZNXN���n	z��ի��E���%�_s0I��/r�n�$駐<B|��	sjC�}��E�4I�1F#��e��n���ē����w�>�Ya���>��,�쨩�;�yA?l�'B��M�g��n��#t5͓�F��<-�����5��� 9Zb��L� g9jqx_��,���WL�	a�\k����A�IRz)��8\������������C��M~R�㯯e�so$�,ޡECs#�^4αI�	P�`ǎ	*����C ��Y2�F��x��L4��!�@�Ke�@�y��G�T,P��WL?�:����;�\je�~�g�<���%��ԇ7N��M��M(��,Y�`I[P[<��Bahm��Q*}��)���_0�Ot�x��&7�sGR��B�r/�Z�.J��\'S�%�uYv��ۮԡ\҇�Ym2�\�G�dR\m$���!��Lc�Y�ujT9r�b��[v���qǟ%a�/)��'�D�O��i!��,%�<N���dC�/��`��	Or�v����$�#1����K��X���#Lr��vDL���J⢧�(bK����M��&�pX�l�8r����7O�P���V��0��GN@y:IPi
��0��e(�AZ@绘�d�qA��4�
8d��	1ш�j���a�ӐP�3�eԝ,��H��,�PXp��8��ۛ�TMsI�)����%��0�&h��j��\6b��}I�\, e�i0����q����h�@E����+�+�R�����:P��*c�g��6wƞ�;|.�@�m|�$|]��ѶNd���T	~N�2	�K:�?"�χ�M�%�4˟��M�Ru��6��r��U� �2���
�a9oR�h�$�H��O�DcB�W�~��v��٠��q�����z谶��{U_�}�*��e�x���/�j6�ڛ!	-L*,��5�N3��r~����7�IlR����@.�=J7��*@��{nͩiw��iՓ���}�"A��΃�լ�h}\
�l��N%K0X}^χR���z�����_q�S�����ᾮ���d���xM[�R�ʹc	ߢW1twg��r�5GE�Zh5	��\T�6=:LlW��h7ՏC%b�+�q�|�VgӾ+��z���C�Ns���v�=:V_ٹ!��I���_Y.��6�r�v/�S�K&XU��e�=��%ʸ|�OxN]�i&n��1M>79�C8e��ר�$8S�w��~����̕<�}�k�r���hី���zK�e��ҁ�oO��ʦC.�fc6���c�yTI޸d��n�����^�g�Z�W$��l1i���P{��PN!��~�i�
�z���j��˴����f���?j��+3:�kPTb.��Nn�"�<T�#l=��=����cj�〡�9wl�e����2��@�T��BxO�B2��['���іl9)����#�ɸ�LP��Qx7V�(n��rW��	$f=����-E��\8)�*��'��3��	�]�EC NYIRiF�{A1�Ў����{�JS�>^U�- �;W�$ĊDr
_��A���-�{x2�.�]j���s2#�Z��p��p��4Ћ��]
wx]������X�n�t����VH2��ZE����.�O'�1�����Ui�#Q��OX��C`�)�Z%��(�&yT�g7���H_���>��c�X=o"� ���%����T^����)UG�J��vF]3C��Ɖ>B�[Ď���Տ�/N_�k$	Eg���3S �'2
�DZj����{�OIB���WR7����jxuv���j�DV�46M�l��>q��K�!�Ǥ�Oi���q؟��X�u� �ZJ�-knM��� �3���H�~! 2���V+��n�� WWr?�j��0���,�m�#�<�~�ɾ���%q"�+�%�>���O$~]C�b�WŸ�11��Ww�Փ����X�9̼޵�xbB�	���'�O�A4$B�<��p������#�QA�e����ʈ�9b'�،m~(5lT�����c�ӹoa��(]c��_I䍲g�'���C4��&�G����� 0m��1���f��1�|����k���S�ˏx-�s�tz��st�R�=�؍�iϸ)8�	�B�mЛ�����k�&�B��8��Z���[���f���r������)<�� u�֥��8Hre�Q#G�Ltu���!��&C�Sqɐ%���ί�A��a��!���E�o�D��T@r����0�kE�[�b��:���a�Z��!�Ŧxz1<]ipp��uX�*$�B��^���-���U���1p�_�n���6��PB��^Lh�ҙ�����˯�sy��Emw����,��,��!�e��y/�-�;�w�蕤��jǀΞ�%�\���U�5b%�	����V��EK�*dw+Y�IY��B���hÏ|�l�՜���7��h�������j��h�NBZ�|q5�NVe����,�{FtHɩJ1����<�FRm<e(�i��r�ZՆ�*��T���*�#�4�cG����<�����V!4^�1�P�V8�с�6#�����L��lQ"
yq��\L�ystQґW�����Q4歶��?F�E5(��^T�Γ���Rr��4��]i1J�6�x�$�
}R�T]�l2U�O/@��D�B��~�*�O�?+,B�,�0���p��G��&�"�u�-^�������C��8��*e�١E����X�󢣞I�%#����}��P�*;�/�����ڌ�����3�đPШ���G'��vI�����+Tv�+���K9l���ɞ����w����ĕ~%i({��Z9�X!��H8e[�$0�ʧ�X(�o�Vi�,G��pZ�{z�Lj^��Kgʵ�OؤxF��6B�r���qamm�c)I���6�,�m!�L�K暃-h��-�".�Y�D��I���+���<������ي;��?�m0��V�x���&�"�x\פ
>���/�¦ǔU�����IN�"�عujKOC����E�2&�����R��B�ɳd�"L�<wC;�&&@�,Z����wUxR�Pe�<�������3�:��В$TI�=�~Fa�'��R��?*�����F����6y�%u;�Wn��%pd�K��E	�/}=�V��KL�#�2���s	&< JT�����8�9r���]�I���$��뙰@�T�)!-}�/�����1�r>')�ɝR�Sbф�2D�p�'�` �?Ĥ����`�{�\�WV?������������C3n��E�?Co�Y|�Rb��#�?\"I���d��0�f��������FH�Ul�1)���˗}ٌm�%3P����!:T�}�4%�ٵ� ����@���P ]N%-���s�~�5A �I(���(�ˎ�t�=���7%�Ր�Ž\~-s���t9�Ob%|�5vK�֣�K�Ab�;Ϊ�+���9h�`6I$v��ˢb1-�z3Z�?���J�Bt
�.�� ���]�K2@P��1�D������^����$�2����X!��8��4� �O�R�H������L��Q�%�g�n*��p�a�?��SY�B�x5�1R���\ߖ�t~�&����{���[���]�Vv� �O�� ��|���s�ۍ�����6y�C�K�8�P�(4�E�΅��'=a���~�ЩN�M����tsK��w
K�:����ZU
���s�z@���=a��g�B�#*iV�yǜ�Oz^�8�s�����`�A�=>�7���r��*J{�|�M(�#�V���
mR��[g{���y�(B�q(�5��ML���tr�7�
H�֒�>����i<�s��m\yq�t������]�{�eCf������-ef.P�%�w.�#�	A���8�M�(��Va�`�.���\#R31��N��V�gJgi�x?t;�i������U1����*hm�s��"
_a���z�	ve�h)�dU,�sr�?��}R �B�>��)�K�_�����P+�d�n�#\tf��7br���ߝ��񶄺��R�&�j�Y~H���$�s!˧�c��Lh& �[i�9��v"ʲ�X��yc�8~qf���/̺E@�N�CXl&���?����$3�<�J%��
�cAB�tr.d���!��K8�#��/5's�NB ~L�O�-����Y��o'K밃X�h��dI�@��q�/Z��9�l�Ì��)���`�Ұi5�L9� ^}h��'롡��U9��%`-��Sgv~,�}����e�L��A����8��~����0x�Ha��3��8���aȚbS��|��{٭[l�l�L��J�n�OPFD.kaD��4�h�`�.>��4vC�#[�dt�>�.����rƤ�*Uc�6~dv�_�･��<#����%�K!/��w�gΉ�Y[a �C~b�VDF�Bl�۹�67M�S-{I�q)��%�5ߤ��Q�Ѝ �|Uh�y]mV|5@��� �:�f�+���1�"�ơwz�
h���8�t��0f��È#�sR��e6���%�E�B�'m����6M���P���G���[�G��)B���пR3�i�}��`����ikk3)N#�s_#��rc-����Jd�Ňq�B9;T�(:Th��Q5�,Vk���f�T)IgY��X�wd�r0*%��z=m�ޭ�';�v=k=<�\O��a��AX�,�^h?>�+p��ߓ/�=.~��pn����(�>���~uI�R�
/�I��O��u���+��i�p��1����o"��)�jQ� ^�^�P��r*���[�WP�&�^.��d��8o�$����V=��s"۫�>gOrT�~�CZ6:t�u�߇�"���GĿuԑc���i����I�:��bJՇ�����v��ax�������%�Gc7�f������pM�Ц�L7��>L�c�w��.�}�����ڌ�c��҄�45.��\F�z��A��O�`�W��ꅩ��j��h�2(MQ]�S~ϵ���_�F��Ll5�uAH82�$��Ԍ"���4�$�!Â�:q�XB�F��$���M����4qC�?��/�#���P�7E�~��t5]s� ��li�ϖeM��X~��
G��8)�k�J����Vd5I�t.?��ε��fA?�>D�7�X߅�)_A����RF��鎤���!V��D����
]��6
(��^Z�7e�s�V��a��[T��u�5��߉^Y�}�g=�;�`�}7w��f�F�(p䳚�Ӵ���v#�U�����
�:ؘF%l-� j����b�q	���2?�ʎҹ}�J�H99^��r���i�/9�i�2
X0�PݹT��AƔ�{�� Fʜ�&���0�=	�����O���/�T�ғ9z)yŻ�{z��"���M_�~�:�Ђ$��I�j�I����5_8&��u�s�3oՖ"T�K����aB�j��-j�ؽ��-����*�I��c�C���IƐ�&
��"�|�!�iȻ^}Qt���*L�J��R�k."ƾdSXvjY+� ޗ��ʭ0�͜E�`�f�o���~�����+E�B�$�� �����k|��.�T}gm;��͐v`�r���FE\E��^N�cX�3-
Qս��]�V�_�Lr�Ԑxԗ�A�>����<ΑS|�����=i��#�lzΰ���������;2&����������x�{���z�)8�1�3��ʛ֐įI�[��x���Ε�.���pd�ذb����{�v��gz�����.o�Ɠ���Еl�%I�24�_S`G�6z�^gq�Yǧ���kߚE��Wg�q��#�j/������~��E��UW�k�	I*:g�Xa0���ϧ������^�3O���
� ��.F������Ù-�<,��P���2
��uJ���ۇƁ���ܚEu+���͂ /�fZ6�����J¤hp�c��Ka�����c.��Q�9L�B�]u>}IBx=��A)�q�hs02o%����=��:��^
A@L��MÜ2շ�Ú��Gk�Y�SqIT�c�v ��`��x�!E� �P�p
��l��Y��Y8��b���D&������^};Q�R��9q	��3�OQ��K�lM�*������q��6|������F>&nīV(Ld�&<��E�m��ډl��c��3�42�J�;2oPA����s��`�2g,":��U2C�i1�P�F��2����㬦��h�l�u�]����[���~Y�.&�1*Al�F�id'S�W}Q:����$�\��Z2��&�l�p"An߮
�B� a;4��U.V//C�V�(��V���CpU����P6���XG��ڃ-�s��KjP�a"M(�f!�&������]v@��~��ť� ��%��J�-��|�F��Z�M*N��������L���S�,��#= X�F�WwC��*��S_�_�F�aW��C�u���D��5�CDιH�.ϱE�J���w��nӲC{���5ZĘ�F2�\�J�a�Ʌ����!�ۅZ�8�9C�r�jx��q%7����U_�Ig����MҀ9z1|�~=���C��L��[�划�<�����Y���~�ލ�7��24���IK�Z5C��ԨS�Nc\�,	w��E^�9����_��C��I6�� �L�S���Q���Y)v\�v����l6$�a`���������7R��{#��Vޅq<\I1N�pm��þC�����.�ځc�Jm����p�G��ӻUAW��b��p�ET��t�5��p�dϞ�`�4�����C?�������
k�{���f�v�GƤ}�)@��<�L13��pa��!	����ڎ8�u�<��e�]�����?C����֡��eִk��`,�������f�� ���3⫁Yo:DyB�P�l�)9���QW�
�spc�(����١<f|�e������!�mR�����v!U�6W
�{�z�Po��K����T�#�]���ՠ�Wc@�Uo�H�iG��V���w�@g�'QX~�U]I�~�� ��\f��M��v�?�kAFJ_����Nӟ�����3daג�ݭ��3l̇4��J�⢰�W��f*�ǭ�ج��ghɇ�{���O*�)�>�	~����isJ�,�@"��cʉ���L �(hq�"�����8�'�56���$j."���F�"�Z�ZN�0( N���~�r�����ZbWO[�7������y�N�B=�D�5U+K&��7�+Eİk�Up���./7�<>���Ӿ����*�T�V��!n[b��*�l�t��Hk�q�~����d&,���*���	cg�;f���)ݕ�A�;b~��zVH��Yo����;��{�趧�W�8���:��{�r��*��u�fJ��gH���㾃�{do�@���|I�'ڪC,R�e�w~%	��]������ �`*F�}0+��@�5y�mmT�Ls2��ch҇�2������!��7}I�	�>����OYP���ȉ�Z,P
�.<z��oC�큄F++�0|��.�X�#9M�l�1*oS0푛�k��t?���7a���f����+@$��w�Ng�[r����V��`��]�9�^����?ÈV��2��Pn�Z ��
��U���8ˁz�P���-J���T���ň%C��w2D>�UǉC f���5��uا?��D��^����C�"��M�>T�Y��(������}��W��Hm�MD�֭L�}̽?�)��)N�..�����$9Y\�w`�΀�bA����*-}���k��쎮�����">��:��n6-�<����Fb�'�B#.6�D�L��2&#F���p>��mx���Ǣ<��?.�`C�]�D��B��܈�vTw'�C��Lt�>[��u�s����������{t3�q�D3���˩E���Ҍ��+��4EѰ��{c]��t<�o_�2�R�Ľa
�������l߹�����s��;x�6�gͼڷ ��f��0�c��M�����yc��������5D��2��%h-��>9���M�{���Z�M��s�l�I]����4&w�����Ĭ���Ъs7u:��M��i��C|��Ķ(�19k>d�4��A9�~��|�w�}}M_Bh��$�#��~��Id��_	��6mý��¥	��~$K��w��3�uۛ�ξ�S$%����gh�"�&�oyV��iʗ�M�E�#C�� �P}M��s��@^P�#��p����k���M=P�Ձ:��ʂn�I�+ �42l`r�ih�̕�m�v�;?in�����wcv��K�~�aC=�CW�f�Qc��ĳ]~H�knO��a��e�A���-��Sz��j�����;0\�:�8��p��,�=�J�z`Ӄ@�m��g\�mϧ�U�9��Т"��-�l��@.'�%ܦ�������:"R'P�Z��[M�P`�d� ����残��	���u8]���Z�ŤUa�� 5��Yp�m64�_��y���eT��I��9qD�#�K�MBb�Su/�X����9��+�ٱ�Nۍr�"�1�-��Co�HGj�K��DM��>W��:��P$
�L`acp:�n��5�>�/*�k�p���f5o�"&��,�,P8���X��Ӭ�H}(-��	>65{r?�0�@�G���A�64C:��⩣�A[��6���=��T�.r�oab�.����۩<·��U/�F7v�[���xkQ���;oI������q�S,Of	ASV�,=Vّ�J=�CŻ��xl��F��9
�.hx�� F��T��Ě:������Ǚ��+=�7�v�K�"��v��90t h#������3�6���\q�X�}��H��R{��K�`�-"�^4tРY�=u�$K�9�^��l�>��8B��J��(	�O��-)��MZ�\�@�1ÜGC]M���Mڡ��TL���2�*�&�A�#��wX�����q�}��z�+��Tp'��\r�2W;R�}t�^��2$����r�����.	_x�_)ԩ8��j�"I��o�Q�5�`�$�gEkќ��_�#�4}�9�����Ǫ�A��g��8=�8� +m���wl��r ��+�E�lw��0�3?޵_�\ހ|գ���}���<X�λ}���ɲGχ+* j���h��ęIDn?Gm$nE3wr8&�!��(<���$�bk�G�5z�@����`��_J]�ˡIf���A����i��A�3L 2'�$��������������]9��~-}��V}.
�hoC!�c/ԇ,^�z*6���5_ �K��l�y�T�C�$_�����9u�d�k���x�5��5�#jc��T>�8�%�(QPzA��=m9Xxp����Ω0��S��DW�������WQ����V{���(f�\�m*3��8&T�ި(v"��)�sp��|�LF�b�8#B{}�U.`n�_���B���2��J�4绮����te���Լ}��8����/K�.9���=-#9k�
�JL�E	����r�.�/�����E9�zw���ve��eAf����49�&n/�Y��g�y�m�e�HBo�Χ���CAB��b�%'p��;��~��e����-�i7�Æ