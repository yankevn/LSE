��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�U�|�=lc�9lee�fj0�e�19�͌��G�G�r㕦&U��\�L�G&�
3�ߏ�"��@w�������7	gapl43�%G�Kh|o��akW~J�,>J�ٍ�RG|�\�R�Z+��Fu��^t].O ����!��FD��u�ߴ��Oo#�+��*��r�C���"�����.>߯[.�p�8��΅9��_-&�b! �B9m�R��jr��V�Y�)�>�G��p�2���l�p��3ܪ��d�"s��}���V���H`ħ�Ç�+�y$`jq6c*QIq�:�0�.���Lz$&1�h�1fu��4	f�e�% ��]3`�%ޥ���:D����\��W��,�ՋnM0yWn�>�Q���|����I���I���l�@���aXǧ0��vQX{��ل��u���k<@�t�şwL�ҝ=Pg3���C?�ǯ��s��ɝ"5�I{�����|���u����n-����g`Ta\��@�=�yw�	n@D&)���3p�1�XINʠG�;�ܖ��̈��N fh��#Jj��nbF5�1�Y�'S t���Z��1��A�Z8:N�{�z�����2���#��6V����8R46��t�?�q������Qy�)F|�PML�͝�2﷩~$� [p��M��.8��W-��_��p�wy�� �ߥ�{dA����ۚo��4��N�	�AN��W�@�O�~"�^R��z!�.�V�¥� ������6g�u��ٍQ�p���|�qp��e׶�J�E��#��G��d�@���1��X��k�Խ6���K���N�D�/�:=t7�.��ߗ��6g�k�˙@��Cް�׿����N%-4�W���u�ο�̊�I���/��u�Q���AqM|��l&�Ȕ���M�nW�(SH=������3��1�����"*�ӫ|�V+_-��&�]�=T"�$*��m
k�.���Fzٔ��L��� �/ð H�P�MN�N]�\��PbS��O�N^`㏥8�I��S�*q1QPA5��U�[��5�v�B������!e�
������}u���p�|��:��#S��:}!�m��E��4�F?��>]w��is���Ƿ��n���[U��;��0dH$�3:`��7ۜ����>����%S]��V=~��r\����.0�ʎ�ՔS�Ͷ_s�w�(\��f]zW�m}�Ę�ur����< ���ѐ�;���9�5OĬ�5��g�a��I�s#£h�ބ�f<�[���S�j�Qa�E���tD�{�(l��yB"*\)�g�~�����j�_nz�ῖ������}(2�9�G��?��/�1����auo�U��LH�
��!I�A�Hc���jm��/�6:�(rc(\��N�$��	R����m1ۢMo�rjH�Ĥ�/9+Գ�`q��/HK!.�Ny ގ�q�X��T��{D.�Z���(��J���4?���x�ȸ�v���WZ�t ��]!��,��S?z3�m�c�,_��f/U���_��>�DU��?r|ړD4p�ބ��I��H%/obk9�N��0�Ǭ����,~��0Eu�.�O�!�����uTr�zVbUK�ž����Y�����z�-;��B2yU�� Щ}2]mZ�W���?Wn~@����-�hGn;�*n�Ӥm�V�nZV��W�$��1�no��"e�GZ�O{Ǵ߲b��)���`��nz�(I^�]�����%�x��J�C`�z ���HS*�د#|�߯px�)B k�����
�$�Z&o΢_/�EҀ�) r�[�E�5��RV*`b�3�����uq��ʮwa n���-�ZsTI��L �A�iXe��%K4��'���ĉoX����w�&���}����`��\��.>���|��y�W7G �Zoga�F��R qΜ���h���H���#�2����u�!�;끄_�M���fGb,��E�%݋���2�~�^���k�#@��a2���$�tP��h>'��7TCch�;���QؔE�݃Ԙ�/A��L.$�	�!*l��uX���Z&�:1���B�h��0��n���y��W��w��,��3ݹY���}qM-͙�v�c�(M��G�hagf�9��dWm$���ߨspv.��F[&2nQA��'�>���񢴾"t���,�"�T2�����f�|{��o|n�sZ@������r�w����v}q���5:��	:V�b�ex��<�ʖ����iJ�����z�H
\Z���P<Ѡ�Nϓع����M����؃iɤe��xm�XS-i3�cja�8Y��!1��*��h��]l�;�B6�'�{Q�����kQ�EL����'\�ſ�ARЄ]���������nr�w���N�}�fw��f�<:���k=p�t%�#�T�G����D��k�c�m�I���h��T�-�g�����Bp��o�yor �>Ʃ��ۋh.j=@��\N�/�f���S�A�;�1dE�p|�{����>��@4�(3�ʳ+f��V���'p&s�e2���Ă��A���..��aM�+��J�<���	!δ�Xd�i�_�'3!����&�U+�&fO��7�@4�Ә)�h/&1M����1|ߒd`��՝{�cK(�ی�8r���,����G�Q6	�=���	2Ӳ~��Sβio�(��Pg}!@��靰���3���M� o�6O�$A�(.8ԏ�u|E{��÷�Ԩ����vu�@l0
��3I��*���B��&L�*d^~���/(�U�x[���>�o�Zf3��ǝ҃P���잱G$7��۫ ?eU;��}���He���G`�6m�԰(�.]`�R��P�_��޾�7[2�no�<��9�E�@9���"@�	'�4ƈ��cl�WX��b�[1�@�T�d��/��T�74�O�Wr�|�8��f{�~B�Q��!����l�A�n��k�i(0��.O�d��0��r>��_�;s\��s&���[~҂s�#��)du���Mk�_���L~>^抵�'b�!v!�d`�_�h	;��� !U���^&�x���H�����&B�e`�	N7	�.-��W?�`� *�8�8Q�D������n:��+V��
dś�&S#�=H�f�?݄�s~׶|·MXwT�>�4}�;�|D y^�	�ҵ�%��m�O��g��\6� ��p��k�I��p?(���(Mh�{\$G�!R�V3\C�?K�[�LVZeO\���O��b׸E�g�?9�oL���F��,�̡l"ʀ�&�*b��JC�d����WY�.(K��^6�ƭF���m�.N��|���b������Ȼ0��	>=����!�]2�5����D��Q�`��<�ZV�'�~G�Mt�8U6$k��3�m�A-��8���3�K�ڻ
���p��S��/G��oJNc��@��(R�u����i�?9ފ�D�	ɤ1N��:� �\��X�����.ʳd���t�g�D�>S!�"��H2�^�)e27�ҕ�v���zC:��$9F^��H�x���z�Aʗ�%�+��ܒ�����~�!o�,l	$�8��M2�F��lSO��a����Y�|����}�Kt�z�uP^Y� �ݤBL@��vM;�D�^����b|�v�?{���T�]~�`�	Kӵ;�K�c~/F�`Ƨ��������T`����'��jK{�J��i�+1M$�k��4���c'h'	V� �E�"�W�K�߯��y���U��ʐ	��s�J[��>>��߉�X��܆��"�B�[�ǯ̏Rj��%7�6E�����n�Ek�6���A� �@�%�f��`f��kͮ'_���FI	n�Eu[�d�2�����s��_U[h'wz�<L<&�k7���bgͱD�g�k�Wy�o���a�����~���sa��f�����}_�FN^;C��G�pI��B���d�k~�"�TT��%���X�VL��m>�eB=<�W�^*���x��cգ"�+����B����ܜEh��s&�ҿ���$jջ�0�ߠ�O���;�������NV(]�Ru6��9��R�8��ƽ��h���8��d�`.�h��s���h]�4�%��kx���'z���7�a��d%�Fja��ba��܇�P��c�u��5����~a25���]*%�ƞ7���?��4^�}�I�=U釅/F�-��-;��d�]x�y��Ԍ�M��T|%�EmR��[I�*����J�U�j�b�l�Gz����q�<�L��9�Z9��i���D�/9����:�o�#�	�C3����J�>;v ����#{]t�3f�����r�]��[���,�t.i:�*�����Q��W�Wn��ܮ���Phbǥ��΀�K�� B��|,d0��G\���_��~�-�g���.�C�*x�#�u1���EQN�:_�*`vi�̑!�j/�l�.��O@���uy_��$�*uh��g\�1���kN�������4Z!XJ'��7�O25�Ѕf~<����4�j���b ]�zL��t���1�rK�/�F�,��B~��gd���Is��s�$�jIS�����{6=�4�U�����~�UY9����yw+�7�YZ�;יaM(�F�m�22*�V��7V#a�0��;v;0�`�v�*7��ت��B����J�"8H�D-J����
81����l�B���ʴ�`��nZV�$.�Cch�Yv�ӑי���n�٥L�T��W�M
�~5ş�1�$ߙ�4�+gp � '���(�ha���N��[=�$E�]Q�f�6��h��J5�φD�
12x ��B@�,�u{�[��a?�6:,�L4��<f�tUjk����N0?�S	�+w����J˄�-��+H��k�^,��~����S�}�.����yI�/� X�-Y�&�oI���~�\�� ^]�䆾v��T*߮�ieaۏd?����G��s��|��4O�s����\	�ݱ�����b	#��Z��o{6B� ��Hn�x�����(<�tG��R��`D�v�z