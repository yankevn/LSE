��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�7�Kۺ~�۪�����b���B�8D"խ~�����:_�����԰w�|'w,
ؐ�on�(�(��c��q���@��������Xj��Sog�a��[<<���a(>z�=vs���i�
B�Y�i7UO�5/-}H�c�U^�b�� �� t �3�\��pW��+�F����e���uс�7��;�����􏿑ܗ�Ȩ+Z��Z����C���=}�:���|��IECM��5��R*;��x`,������;&<@VG�� 2�36"�S�܆�'��s[%4WT���±r�� 6P�����s�~��(�>�5�N�wTe�4y���)�Ũ�Bx���ζD=�z��!�Ǆ+���U���{ft���i�Y�B{K�G�Ru{�s�#u*���E����@ɦ={�*4��.O��, ���k�B��p|DvZ�j5j�����t<���>�k�!�cH�����@�s�_J��m��YF�d�":��t�vBâ��7{{ΐ^�/��p��D�Ep�[��F�V���ie�5<r*}c�5��^������|.�=w�ݬ�t�Z���={LECZ�$�Gr�Y_�s��VF��͂A�w�Y.Sy�鉛�a��҃S1�Y�ӗ��PV-f�����SE�M�V�W����=��{ϰh��7�8��}��V�`�s>8`|��~�����݇�O���j�${䌖Tq��]���RtF@녩B8�c!#T��)��vb:�?������ۻ��>�W�A��E�I66��x�S��[O
�	��\�𡮣wo�/��Ao�ݢ������tm�N��B�;	$��}����l� Ԃ�<��C�����ɃܷӴ���Y�ⶥ��l��ά��y�ݮr�nu(�A�-�Ș�(�	��}�	:���f�ƭ��b�mD�*���#Q_�A�E�ddLX����<��1���#-ev�#��*I%p�?�Y/��Fe���q�)�� j����@���/� $��ď"��®�=Γ.X>(�M��8�g)�,�6�EAu��=�+�W>u%��7#�{�q����VSʕ��G�����ﯱŊ��;Rԉ?+3�vɟc�����XTHh���v��\DM�ªs-Ǣ3��u��f��XUl�b�x2"[��T����<ȩv��R��Y]9M�h?1N��v�����[)�ױA�@e�2A�s�1�y�'z���4��TBAg�xg��wXg�<�@S��t1��U�,�a.�=�_��o'(3�R������ЭXX{�X�U2,@�ɰEUhj����6i�ƃ�CA*lE���r��l��0C���|��$��~9Aѯ�����o<������0t�6�l=�9����.PS��(�ܹT��
RR\�ԭ����PP)��6F6��B��X�zIx�ՠ����,{J�� &%{{x��Z�њKmlG-CKDj�,�`��c�+�wl�X��(���܌�+({�S(�E6�V� �l�s���̮Y�vN��V�p9���'��� Ѿ�vu=��*œ³������<*ar8��Z'\��W9��5�K�
a���Q�ב��1�d�߹�܅9>��a����EԀ�+�ȓ��׶����:=_�}�ѡ&�@IC�G�)�v��9���)����]}��.`���=��_���u�U�+��Jl{c�\M�$�����O�`���8��=zP��"�<w��V��{l���jlzG�3gM�6��y�	�
}��D�q���n�V��E*�;�s��9Lo=k0�ȉ��b���R���ݞ�?�侦y;�.q�aI)LV��"�;�'o���5K���\/�q~%�r�U��c�3�)�=�:��4��6C�d�c��H3M�[C"��Y�~
c���9�D���
���;G�b䳆�7�UE��~i�H����SN6̼�AM�~d1���K�l��l�|ݹ��Y}�*ɕ,t�Q�ɞ��aA�ʲ��_aG�����!��œ�Ӎ2����L8\�8����뮔�U(_����{����1�]'b�=ԥPy kfؠ��,~Q�-�W�CN�[e�;D"�k�T�С�<_K�0�}`��@�^!��+\��G��v �(�GD�g���9�~�	6����N�B�/��[|�5�DU�$���$B}!��)�i!ei��|J\��3K��RH�B~��a�C���v}i"!E�Y��}9w��E�F!��^7�<����Y�e�
� ����(8߶���3�-F��@�]T�P��{u/H���`)�|;4_��^�`�Dr&C���aJ��"��VG6��1�d2��?L�m!�~g(l�>�k���	��ʃ,�����ޞ�B�h<iFݵ�`��⹶�q��4vŀ0U#p���U�!�AF��/zn��v�`�w� ��3y�¹F�������Sh�-0_/[��s�ں��l:�5���зo֡���	��D&�31���	0��l��YV���`�������9;��Ϗ)=u��ڶ��e�����Ya��v4�Q� �\dp��Q*�Ǆ%��Sr�|�ì�|)��Xi2��TICCy(����)�pb
�8�8�,��)vaJ?<_?�˓32'4�rJ�X����5��!���z$�T����m�Li9Xi[a#M?N��N��	|�2O������Prf�@�� �jo��e�h+^J#��
��[X��b������m#Dğ\F��x�n���$} z6*���%?-��Mj3���~���֍��Do[�g��_`@��6�TN�`�(������^
���!p߀����\��U o�~mguI�0�|]J��P�KhSL�xl�i��`�2
�Dg<�R�O�ʬ� :�F���S{��lY�]F*�L��~��O'���+�N�j~v�x�'�w^R�v�ޮj��M�{�'@aAe�
��ϩu�0�vs{��2<)x��6��F��з� }
�]�-~��[u�����lQ6�L5��-����Bw�jR>��E��g������QV�����"�4��iM�l�==����k�˺�k܏)�%?��=����7� �A�����6��$l��n��#6�i8��p�[����Y��:���+�����R����y�OBT��S��M�g���� g>��������"<|p�(8��?���"��$�r8���~�F�_ob��]���4΢[\�H�^)�&�-���k��=)��%���e�~�8��[-�K�{�8׬1�*J����ء��2a?��D�É���C8{�t�����5EnA8�!8�G�P����A5>�15�����=�o@%�	��*t����U�$z�nX�7�v"w�����y����HzL�(�S�W��&�,����iQBͿi��
�ʥ}��n~����^�U�߿ɮn����l��5�y��\��l�r�-2D�"�<|P\E�`�g��@ɫ�I�FYu��)r�9G��TeR�����PXX,B�p�3��B��[8���FݨˬX����>mH�K�aƍ��t�uV�eЬȭ ��6�d�uI0�`�I|>����*�$�J�+WA���]���a�+f�=e��M���ť����MQnd
��k�c� �a����B=u�i*CM?��r��bu䎘�$�bt���ȴ��xp�zǫ���m�a)A�{������x���v#������m�\�54������@/�.�� �({�����$5�UPw�-��c����w/�Y �h4������s{t27�Z���׬tĒ0�!m9��e����!��%t�T�̨bx@��~DA�^2���fyP,$ �s��VE#���J�1���u"M[!%osT���<þyg��q-_��D�os\�.�A��a��S�ⱊ�J�>M����_
�n�禍��\*G��B�<��l��W�J"��q�|e��w���4��)�����i 6ֈOݍG�*Hm֖L��߇����{m:^N���PR���dU&��͠������v�iso�sP��CW����%�?%�n��l��UEf��炾+���uuF�{�W��@��4�G&���%)�0C�%��;�`&,����%��µ6{����Lnd]�žh-VlJEvjc�6����+��_�/E.]�t�8�����C��12�)�r���e�/�~
5���h�_�߇@���D����iՑ!��֧��X�k�n�l[� �?F�Ԗn�����j�Y�M|�+�.A��3��)���p�9l��t(����V�I�ފ��祂z�xEA�d���X�߇Q�lQs9z��	�R2*����-g�1)癵��g.��$��~��m�e@#�����9�]�������ug��)�Aҵ�T�^����o��|CĀ��J������lm�ƒ��d-
�ὲ@���uǎ"mᦨ���y����{�<5 6A�|ƒB������s`����H�Iq&�௬�Wf��`^�V�&E�Io� ��g&��&Iȡ�G��P]�v%lX�V��¦wJ������I�I�Rv��G���I1�<���(�B1�n���T���C|m)�:�L����Q>}T� ����Ĥ'c|׷Z��0��j'�9'����⺀g�3~[�)��X�-�_�|��Z�#|�Jȳ :�p�5�(�Y