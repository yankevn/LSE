��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S����)1�
�f?y��pI袞��f����M�Do�1�����4<��y*җ%��J(�h4m��z=�)c'����>���o��.�d�k�$z���W��''�������r�g����Я�0��5Jl��k�ȇ)�S��
���H��A��H��T�L6��v��l�Y�H��I���/�d��W#��xZ��+���UV��s|Ly�J�¸���$EQ�����bn�O���¤6wl�":�sa~��pؽ��',��'�^����s�;��4���
�N:��p\?�U��e=w�
垟ڟ�ߦ<m�b���S?�	�4��E8��.R�,k��L��_B9nI{ 閎�"8׸D��:�6�^�k���K]����^�2R�E���K�4��U���q(Zq��ȗrU�F���A���5ǕZ���;ҟ@�[1^�;����hi��2B`D��|Q��E�$H"#$.-��\r��sЗk��i��(�gȁ�+RZ���;��Jñ��]FZg;2Uy���haQ������&��c;�_���JPq���-fj�8iI8(+[���?Y�}��^�Ǒ3T�:�����:s�P8�Oϣ��v`\��K�����?����e�!���s쿕���P��E������%\�k�
'SwslR�N��V����������CL�d��N/��w!��E:B~a�s� C'��6Y���u��I���I���Fq,�b�d�Έ��]Z��"ا�%�c�#�C2D��qMk���J��}LG�%����,^��� K��_�gO%��z�$��k'�X���*�r�h�����M&Y3��n�w�� �ڌ�E���b늚��D�U,ݼDmg2 ��l��5������G,���;M�b2#��R�g�XP�̙_l�� Oݩ��πE�k_G�ev&�JŘ�d,U����i�%z���G7"������	S�5$�to��Ź�/v���dDyK4��N'0�[�(r'd�I:%��^%��!jI	�� �i�x$x����=@&p�����2B1*�%����k5��#��9��s������"y������*�U�8$C���W3�(��k�8%H����6j �~E�l���g���Vy��O͙�V<�XO�|����?�N�2��)�h1��a�鷧���J���/Gt��Ã8���I�p$g�;�����pl�}���ƏMY ���1��q��I2>� Ym���d����>��ce[ӚŮ5 ���^���Yӏ��}o,K�X�U���}�j�dZ_r_��;�{��A���8����kw'�-�CӲ��iS�&�%r�fzˏSv	�W��K��~`J1�(��И������$�_�ZrJ4�ۡ�zeհ���i��~���wږ���Y9��g;����"�cH�S�Jm�	W~ak�C63s�X�J<�4�q���r	���N�.�Ӭ���&�8��#����Z��	K�
a���Z�Q����:4Y���]�j���x|_��9��/�)�V7+�~�a��iM�f��>v��Nb�M9��=8W��D���qz*(�gb�ІV�}AE0�}pF�����Z����/ʒ�H���� ��
7�e&s�̊$��U�#Gc�LwIH�X���hLк��O����������x�l^�+�퐀bZqy��\��pǠf&�93'��k�Yǈ=��u��)y���Q��8Y�_֮�{$9��@r�S�\�:�X�R��L]���x�����^����w�Q�g���h�wv*��YJb�j
v�ڕM"�0�3t;ڎ�}*g�v��`��@�tb��Ѱ�<��x�yU}#댅�Eش�S�b*I�o�L;�Y��j�b���(����/��h֔t��E|m	���-�e�4��m��I/17�-v3��:З�.�:��,�{�J��-m�R���u��9V��oU/]^2�^ ;�"���_�Heg��������B�����3�M�w�E�u@�@����\L2#t3�{m-���a�Pzl��������X\j�'@=�c[TT�H9�Pn�>�Q{����z�������v!r�1C��ƱN����6[��㕲]�p�mV_](����ݽ@Ι�vr,�H�E1����m6�yJ5�ܴ�t7փ��So-W<SBtzK�|Չl�oR���B6�O��E&�K)�6����&@��s*KWW�9�/H�_|� �C���k��!_��<��݅�=��"[f�9��!�3��w|t��;�Y�iG�O:��� tQƑL��/���?՛��(��	��RQ=�E�;hS��{ѣ.~R����i�.����2^��Zm3M퐡���T
ߪ�)d�`L�4�C;#��Kc�1�׽m�6^�W��m�Sl��� @_\E�l�E����=��o�wy~�㑋�p�x�!3�U`lQ(f�������#/;����Kpb��B9#o/�2j��|V�XL��u������}`�To]ɸL�!�y��b�xm�QQ��H]hQ]�����D����"^�n"ɦ˳��i�3���J�T�\3�l���E�N��I�p�\Xw/-�4�Z�h�1�{�t	�NЭo��
w��aM��bC�Kc�����ѳx��x�~����[�׍�-��,a���������;�9l5��M���5�Xjf2~U�T����,�Rt|�q>�S-s�J�S������/�hŞ��H��U�NtU2E�,n�o�������p�zx�;���;�CK�_l��$��2�лG�~+�3�ԉs#δ��s��^���I�!G��/��h������6�RCE"u���	��$��,��ji�&���򿷺�d��%�TLP!33��[�3Mpx�К�W�=�ۀD1ףY���G�}� ��G#�]d��d��)=E��r�[�]��24�zƦ��g���a�4�C�B�!ڱ�8�^=mªX�9/��S��� �}�j�%_t���`st�e)8���n����������/����LޚZu�����t�����
�,X|�{����_/�Θ��e��f�G���dETg�VT�קr�j�i]�-�
���`����J�{�8�,iKٍdk:G�y/����^�f����W�|��H����U��cL]�Uw;�0�]l���$�˫����k,�%�H���}�u7���;F
r��������w~=5�G(��QM����&`C;�-	-����H��Ńb������������m^���+�K����t=�RG�nA�%���VuҰ��P�+Fkv�f���`S9p�2UsO�P�~���nQ{&^D��������42%��Ɗo������1����O�x�N�#D�q0�k��ꯘu�ɮU�������&��$V�3-
ʙ'�|���5�_���\��Ci L��ism�Ln�1܅;�賽�auB�v$�Bnrnd���Lfꩌ���J�����R��L+I��c��Z�GE(�U���,��ȏ n	��ds[q=�#��|�X��.���*��I��K)���|�;��1�B!�#��,�%<݉�k[sژ?Ȭ&����`}b�-"M���hO7i՗�ZHW�(�����Z�ش,���
A�%.�Sݎ��P��Qf�<W��Bz��a&WW��׈8	|6�y��b��}6��:��W@�k�p�E�v�u!�񕾭h��K��[h~���Z����A���JL�_�<?Lu�xc��+9S��m����}	{mU�@d�Xy-DF���7}5Q�L�T ����,B8g��aNk���O[�K����[)0s�Y�L��*�y�fK\�X�<���N�'R;Iȃ�2~�ԏ�~�y	���E�B�_:��l5��`1Q�E�ߤ��/�A�W����	���	���D����HOr>�k��|�ɵ�-ʥwKsL���v�p���et%�1ܙ���V=��o���}�?HJQ a�X��@��6,^�1w
4�'JR#Y>��4� P�7�~�Oi�Ӎ!�L���w��Yhu.�aS�ܺ�}|��pHƈ&F��Vt���,e��|iGϓ�s��3���b���pi,굵_0[x�Ǎ����W^�!񺡁��h+�.��^��Hs�\��58��"8��l#3�f���(�<	��z+�g����S׋!q$���
�6�!��P��ՋC��.(2�w+ˍ�m�I'/y��<ۻ�}��V���Q@5$��t���gł�����ͫ�UD�A1w![�w�A'�ZG�|3��������غ�W"�S,X��i����0��I��W�΅������ˣ6�?3N���D��bol��.6*��t"Ӎ(�F���r����봾,��d��-��o��6�@_�= G�R=ъ�f��*;ؚ]Yp��	M�X��G���}�k3� F/���&���atJ�m��2��H�k~b	 �Ur��G.$�l��rĚ�����1K`J�Z+��~��`�g�2>�	:��sx2S��۔Nd��])sS6�����GB)W)����f����d��i_�ŏ��)]��=R1�{��S�����F	�����	�WY�俩v�����.)\�Ÿ2����_�y�=�g*g潜�`G�I�c{`R�� "�na�5�˦�v=Wr��w��3�X�!�	�kұ0�"��1[�va�4�! ��9$�˽.� QYb�V
�xzl���Bp��|�Q���)��� l?�x��f�˾˗�����V�W|0,5@ޡ����f�w�Q��;^�P<���a�P�R*����QM\�}�����.�T)h��b녅�����N@�~�q9���_�BWxfuxC
~�R�}/�.][�����N�o۫�ᇔ[���Rb�/"r>�u��!�����I���Ĳ�m fa��{0���@Q�<��}�	��!t�����L'�j���ʆ���s'���_��3�W��ͪ�e��#	���r
��m��28�{���@����
E�]��t�m�J,�5.�Zw0W(��;e�j��u���V��m���Pi���3��p(�ۉ��A����U`��b|浪����;!�ڙĕM9��>���|94���- ������r0���%Z�o��]!t��.cYԣ�	H��6�*���H���`�E�����H�_�>\X�,��R���?=��w���	<�V#� 6z$���3���{�d
����`d��=��WcFШ��/
Ӧ�[#�v98�N�ީ��<<���dsDMn�?ƒ��\�9��h`rZW���(���&���S��$�,����o)]�&���v#�uz�ز���`pVՕ�Ȼ�;52�UT����x��i�	n�g��j��%�-D�;g>�q��x�L��M��<&�>����2y#����G�Ň0%ߪ�a�����S͐gG�h�����r�������[Lr�2Q�I���3��*?m;k�.���� Q���H{*j%�u�*4�����v+xk%gR�.sG�5��*��H��l�Ւ�äD��*�#p�.��j"�P��r�ѧ��x�_����ba���l�5\O~~_�i�>�R��Kp,�}�*�L��\/(�{5�1F��s͐�ơ�8-�R�^KM��;�s�K����"��.���vR?�,��ً!�C]��r��S*��ط�����y'���?��u>��N�"H���x�p����_~�\���[H�h����~�E�S�����.��^��'��a���B�[��e^��徝�Se�`[:9!���ЎGO2Z_z)���=�I瓣��)�hY�����O(�����!�0sѳ�ﶆ	2��tk�JvFc��ޝ�3��O2�����n��c~����7�&�7Y�jP�aKn�|�0w����F����ܒ�4P���H]�x!q�P�܋��������[�M�"�����E�9� ?�o��FZD,��˝����es6�ü?�tS�?���Ͳ�7�!�?��x��m��E��>��j�A�G� �o|<��HK�$����LC�ҁ8�F:�gub��|����w�|����R���8E���єA�����,�l�W��扲uQl$�/���-�SZɁ�����w�_��3]H�������I���j)�%�z�t����A<�����=~�}��_�g;��ࣥµJD�}Fat�d���T�r�����|���@l�li���H�%S�4	������3ק�H&�Ntar�?��W��7�s�+��gC�-D������g�J/�����%~�N!����'�����hD�H�S��z����;��b���m���)��u�ˁ	�uV��͏���|$��%�t�J� �iI�ܖ	|�|�R+uѮ��
��y�����2�����<c�[�a|���^�J�����H�SLle�����P�̫�E�Eպ��L�Z�@O�>�*�lw[�1L�9՛�Q�3�P�*L������)��]�� /�&�J��P]BJ�ղ�NC��5�X��e�@;��~硌�T(H�?��p'�6N������FBb�fD*�Y�2M�_Y}�
�M�����GOA(7¥�ʵt�����դ�*�{rvh������sH?jO7����"t`SqQ�� �.�!�4�jv )������]��tU㫃P��G�;���^^�o�k[�����䀌��.�J!$���&0Z�7c#�B���$so�b�L�!��<&�M1�=E��8R|wQ����j�U���n?`X�'�z��$��~F�/�W�R�2��[[ �~+�ܝ9�����n�
�hTu�uL22�븍��|���*���#��S��=�Y����o�R����yJ����̟0�ݏq��