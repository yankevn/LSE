��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#�������xڢB�߉�u�=���=t��K?��W
�"dm^ 
�a������^��7�[������^xf}�!�0�U�'#��sǫG�Vꪇ�|\��&��$a֐�m�ЁAHogķ@MzL�ʏ����iM5��N{��M�h�xȈ��1c�'����]����戄V�E���(�b�y �Z[�]�@[_�k�TNI����TC�	�HK;��F��\O�V��>{z���[�1��*�M�t�ޝ;,3�)�zZ�i���U3�m�#�^�0p�G���K&.l��]v��bN��<{��>@*�_��Z�}$�*�0�Y؎K��;J||�[.�Ԗ���B�,dH��u�TQ8IzK�k0�u60[y`ǔٱ�)V=$kn��Yt#\�o�bJD`"|�*���(
� ߁�D�卵YJ"m�T�`e$�� ��$͞�M�j�"o�"C���D����{��ႄ�ly��?<����:��e�VV6J��h<��z��!����b�K)E���b�.�V;%�n����%�
��2B�N���.Q����Zpzz�΢*w V��X��v�*A �V�����n ހ8��;��gP�Vb��v�嚨�?�F��v2���(��]#q����#�֬k4��YU� ��	�gd΃�\���>?�D>��[uo��A�B`��<d0v��M;�ډ,�l�@�~�@�G@�z3o���ag�U�S�[�� �l�Z�i�! *�x`���Vl��zCm!�o���p��f�|����D�)�!��ea���fQu��}!Z	�EJk{�_y���0d1�W����Զ�� ��M������V~�8hwJ\#Q�l��բ���}��/��z�ZR�Fpp|:___iC�.�SDq���d kPo&�	���5�C���e#��h� �@g�S�˫Hr��,�H���M�	��zJF�H&&6,b<0�qG���x:����v��O}�2�o%�ώ�/I�>گ�2�gK�%�T4�{a�g���P�
��WY)���!)<��1�_���?�$*�#��Y:ʌ�������NH�%�C�5�I�v<��oѩ�`�\�"C�C�_w�P��Q��'�rl�=0��aej���# ���1�f37���-���?��e/�bt��hZA�ٴ�\ZW��R%hw#p�eΒk_r]���`���W�P{(�����1�}�Jz$~DB_ŗ��{7��;�~��7@����ާ�OF�/f�3t�~���ޔ����~�:�fj}���+mfG����������;�.Β��z���`y�xo�^�(g��:�!�w�
?x>�_�w*�	E�2�
	�L�>�.C���FY����pľ�QK��0�}���	+},;@�$L�K��͚����τ�
=������α튫�(
�]�oݎ
���\oR:㤦
��B"G���!��k��֭�`�2�;��F��}A���r舰�;�9Z=�����I+�؉*`�I�����R��֦�X!=�l�%,/�Z�����~���g(�['�Y�V ow"���@/��+�k�{�ԐP���l��,U�#�
O�LQ}�>����Ez���N�t�%���]*��k����C�E<sǝ���lT2O܌���é�U�zSW��������?��u���u�m�,�����T��f��.ʱ��[��7v�<��:�i�<��6���GH~�-.�п��$���P&s,?t�� mA��]�J�R=5B'`�Id]�3l���8gci���	��͙��x~�Dy*X��62��H��kL,mH�\P��{�ac�|Z܈��nO:Lp�+�סE��8t�I�4UM�bP_PR���}^Y0�U�IY��ʭ3E��H���G�X6~kn�}Ғ�d���OZ�ȗk��k�]�dVEu̇%�rցӣ�Q뵓�j��QC�=|�uLsT��f���qtrU6A��_U����.,��j}��4;�[*�+�������ܲ8���ײ8����b�*r��4޵@A�Y��� aa�E�/������91Gt���9&��X���f��V�#.���n�D�ϔ�b-�{��v4L]�¼^]�y�$o�-D�m]�����L�C�أ��m d��=g�������A�]�{w%�}�"�
Z��������9�={��n��G	�]ەY��zc���``l ��%Z�x��Z�ȧ�R���{�af�D�sLLL�Z"���wINaKB�L�d�e��O��8��.M�����V��s�B�-���r�&Zs�C�w�h�xv�8���.z��HF�h
k��}�;H����m��tL!2s�d�ܹ1O
6s�A�?�A�㛒'��p�����ȶ��N��Ŷ�ڢR�W{m�ĳJH<���d����B�i��9?v����#!�%����m���g��6�o����8s Wڵ�������6O@z��f�g��k�� OS� ��`�ogf�^!���"c����C��̋^��L4�5},������utx��l�����l��ϔ�`���q��`��3~�}ԑI�UC�7�\�T���?ˈ<spc�)��'X^�KE�H@ˍM�� ��{&�>q�Vs����4�6i�����XB�m�����ǂ�8A����iy�������<�1$�ܸ�Pb{�2�Y-�c`�&����J�^K�'0�B�������,�X)��,�j���88����fYS�G|���Z��1^O�oڈ���ӄ�o5�u�s�_y�Z����ū5φ�!��N�ƃ�d4_��'+�j��=�>�J��n���ɏ@��q+�;�{A	����`V(��B1����T���Yg��k$X]Rj=4�5��8F�*�F�8�bs	P��ȗ+uz@��]b��d��W=��aؔ�k��{����+�6�����{1�v]�㋌��!��>j/�U��.��/_A�A���n��tϖ�v��
 �̼��z��q��^w;��,����vLM�����������$��c�*���6�\���Ef'	�Y�� �TtUƶ�"]Ӣ��Xmc��<�⼚!�Qx�s_Fs#�>k�Y)�����; �ܮV#,A�c�� �c �1`���W�2��[AP��&[en����NP.�*.��^U�'�J���׽��^i��a���Y��
Q�t�8e>�XPoY���t{I١��(�Ok����蠴��mu���Ԭ�SN�ޜ�Q'#|�`(^qmc;<��x���T4nJ;���&�Uz0�Y�/ͤ����a�{�,��)Vi��P^�Q��r�P~�h�8}��y�(<#��UZ��V���Q#U_�2S�"���t_[�.T��k��S)�[9È~^���.CO��.��g���x���$s
t�;T	_���	#'����Qן��Q��|��?��Ť����X`B�V�Qᇓ�e�1�J��IM_n���<B$�SY�w����V�Di��2����N��%����`�:a���,���2��	y�J��e�5���m����`п?ی{p��~`�sC�t�J3�%�̴d�C�B٨�R��0�o���1��1c�N!��m^8R�5����X�W�.�x�Ew���;�!��1�T��*j�#�rhBM}mB�31�7umA�_���Q����|�6;�갳l(Bc�+z���{���+o�⏞�>Q3� p��h���l������5�����u`OْMi � ����0�l��-߸�|�	��T�%����\7?_\$����B]���j���w��C{Tm�);3�D�R���W7���:���e?�� �~�k2Q��X(*���s��#i�1����2��5 �s{�/����X�
������Fxb+D륐=���*Jk��w�Wz�&G3Z�[OΦ^A��c:kLD>�ub���K��ן	bً)�M,�a`�~��4�$����E���Jh��D%��ԭ&^gv�t[�4��R0��E���Y���&5��������a*��c��u?Zt������J6f�R$܍ªE��6a�N����r[��:�F��\@� W�9���N��`�-C��۟�i�)�y���"BW_�_���J��Uī*NDS�)+�-3`��2�g�|�j�߯�6 �*����Ƹ;{j?��dR��	�4�p7��	��8	=�,���<�����=r��Jj�/ʏ3|@=��p�ӊ�	�K%P�U(�,�ϻ��W��T#E=��)�� ��fbn���ݏP��F�PB5]�������)_�,&��d�\\FY����7b��W�"��~��猖�d8�ͦ:Hʗ� N�Z1���)�)��zU��Kf�n뭒lofIa]Ǔ+e�Ȉc��6��nG�Zj[_U���r5��/�Z�9�|�US<�j�7˳@�`��!4C�%ԛu�A��9/9�a��{[��F3���dI���dQ�4���a%#�*ײ�h����^�f�:?�6����D��v�Ñ��� CE�����s�e����jk���I>��b��3F�'�{6�-4&~k�y�r��V����C���@�;�з˱p7�U|����C	L��F�Z�X���e���m�ÅT'
��t>��mh�G_��c95�)L~����|��Uz��C���������
*��kR�3��L
�q�4R[?�|a۠���E05!��xC�.P<���S�K�K</$ƍ|^=�4z͸��IdL?M���TF�N���<4rB��t���>�N��Y����=��9������2@�>>6���Z�P�i^}��.m��f��=�6�l���7����0��Z#`4ß곓�6�Jː�C�i[��T�-��������GYσ���{a _Nߔ�fJ�ITp�t��=K��
�ƙ�@��~��G�b�4��tz@��F�l\?$#6Ѡ=�3�:l�E���(]�v��n��xGú@L3���R�1
���,�<[�&���v�/VVSo}{�$ȳ�<�^�r���Q,._>Y�%U���p�jS��Ґڑ:Kf��E��G3�h���1t�L�2�S̡iRₕ�w&K��rG�B���V�������љ���|>B}�p�B�Q�)����s{�o�W��;z�bq�$�7	?���\�H����ۂ���g�ލ�̀���1xh�
�>������P�~舶��QOG("���s3@On��2�u?����I�8g�JV���R;|�	+�V��,�����O��!�t�w��T����]y�7��Rh�D�D�lt\A������G?�5#I�����wl{O ��*����K(p1�m/ӛ����.9�<�lM-�si����k_�A��p��;G����q�X�=A,�j���Ԕ�_����ȇ^�	�j�o��ܝ]�OK��F'��g��ո:_}a��g�� ��.p��������EG_�֙�x�K�yI�xy���d!_]<��|��՛�d����/RTBbs����C.�&ُA�_�P٫���/N���Zg�M��X��*�h�T�����@Z¦���.�����~s,��uO�
 D�"f���Jӣ_�u�I'
�n�-��\�_Z�o���H���q��"���k�����k/N!w8>�C��B�QoI���R�4�Aa�R��6r:�f�"(��W���>>W�q��_x[�48��O.��We�'R9Q�'o�k� {��דZ�>��O�t�
xBK��g۽j���3�P�+ka�'�<IŹ�0�EɊ��!�������Ql����`�υz���n�����>�5L�A]~º�=Ѭ�T��7����A��8!�L�<���ٱ�2��c���A��<Txh]��Z�n:-�E)�믳�Z�FZ��O�b(��=jW;���se��N�]}0t�����nUK�^:|
J�N���7�D���@[�2?��9�|��x���D��C�׀J	d!G�,�i+9k�J#�B2
�g�:����3�U�,x�[����=��F#�ӏ[�M�೷����L��<4f��w�c4h�Mڊ�퓺���+6+^և	5�h�?�L��(������?�1����x?X:�ݎ��"���-'�ҵ�e�˗1�W�5�(�d\.���硪�I��6ۺ��#QO��:PgP�[ϭ��}���E�
c���<�ힾH=o4��~b���Ԑ^6^@���Ό_t���L��֘��M�� s����ގ��p���̥�q��=���j8��@y*ݗ5
�^b���l�2<ɬ?�Xr#��rm��ș ���_*�{9R"�������˒�Cp�0	��9L*$G�B˾�Sޅ����v_溼t7�K�T���uLek�6v�'�#�Oi�Xu�4�Ւ����3���uk^�38�,D9�;���@߆.�V���"�w,a��>�L<���$f²�̮�p"��^��{�\JLձ�/��kD�1�=�`��ք�������\x����@_���l�<8�%#�̿j_���_�42T=P3�$T��׭��
�!��D�ئ��ܡ���m	s���jS�+PQ;��Ȇ;�ʷ�/i0��4A)�čO�N:x)�K�$��!�M>�3r����x��BP9�@�}��F��E!� &���逄&8���� q7���<��.�kgfD$�Ybh�44f��=�s�PL�_Cyu�w8̂_1EÒ�j�箙�Ǔ)���ć&ef`qet�(Kd?�!�u�g�s���μ7�H N*�����������z�q�O ƒ8:��",z��dn^�W=��'�G��R��x�u��33�b�b\z�\=��gg芶�����?�x��ȑ�� �e1�1�zR&?-q�W!��L��T�:z��b��b�����r(b�#h8Ҫd=��Ҷ��I�Y-��=K6pf��Z�(M9�u��uݡYhmuP��193��
�e]!`�\���1P?����뤆r�k���P�u�y�1�U��k�I	±��>/0s"ѷ/�@�	|H�2�J/�
"�w��\��ZbY�I�cY7OeS�oӝE`�����@��,P��o�="���s ޙ��%ϫ$�3��3����<�I��}ʄa-З)������.|�2겥Q�%w�\��j��dv�t��>�lDh@�d@�b�E�[c���ǹ�He�%j��PGٛp����N{�}'p5xZ/b���#%WF��o䖓��V���u�'��S�~T#�b�I�z[W�r��L�l�:�	��X�&���J�yY��C(�g����5z�晠Ϛ_bYp���o�q9����r| 6m,G�S�_���&�d��-��
��7b��(��˾��G����5�ѐ7�Kd j��+�<�S[�(�y���+m[�F��ϵ�4����^_�FTx�<�9^:� ��0~�ά+��E�`���ҜD�� �*-0Gm�6���S�����2�:}w ��bn�}�����?m�w�ȴ٣;׌"�d��ݫ�ve|�F*��iPr���J��f4�O���U�,�F��3��I�캠���ʉ���2��I�¿��X2�����)/��"��:�r}-z�q��(�>�a'�A<�Ƥ�J)�T�'f�J��\��u�\��:*�m09�_-�����p\;{Y=��/���	� ��]>K�-yU�Ƃ�줗܂�jqI��:JP�/h)�	)I8�1���xD@�X'� ��'=�)���z��:g[@J�^��)�8obnL�WN���2{������-g�����[���:�/���^kY���A���񉃄(���h�O�UY�S�tx�V��p���;:y|<��W<�b�'�.O�jhl�7\B��%M�������Bhy�c�,��R�6!���S�EC��	�X�/b�K4U7�Wf�Y��_�-�J�݄������
���I�ц+�e��=Ա=s�:�J<�/nP���C�J���d�(��o�\���ҧ	*�{C�U��7v̏O6�ʶadeSt]�|��*AZ.��Ǐ�������<'��x>l}׼�/��������Cu�����\� ��0���M��zYF�<5}���������l��;�b�X�/��
�5с������oȮ�����"�sW����;wX���Y8Io:�H!���#D�I��M�$[�J��Z�p]�,��mފ��ބ��p��]a�0S���� �׶�>�i�"������G��*��4y�.ҍ#�IM����N8㹷�b�����Ly�����!�N��C ˹�#�Tگ