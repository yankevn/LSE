��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~�>:N��c#D8�]GY��cN���+Qǹp�#�C�Wi��RΛEa�-$�p�����[�N����U�;�#�g��m�ն�u����,=Y5�`�9���a�qI�b�PL���� ϸ�1[\%#U�%{ ��{(^���wJ	Aj�P��С�w��s���i���s���d��8x��%����P�X_SoP��ؼW���TE�Q`�"�-��":��LF�I*�E�M~�U/�dy�×Jn���B��h^"lX-�,�L��#�����?{��%�CT[�C�W���J�LR�F�7������]ؔN�2Ib
)x��C����;&(��4�y �	��ٝJ!��Anh���<M16�jn:�`��4͖k���qHH>C:��ᖉ�@V����F�i�9��noQ2�jo'��	�	�w��cq ���?�w��ԓj+��!�&��_�\��!Q� X��Ӑ(y/����FX�E�OKW�L8�>��Yw@`x��0�𱌄R@�1M,�)_��qp�`�*�}�E�:�9��&J|��{T���-��2��N�s<���l63��!�8I��p1�fK�Ŏ�¿Xm_'Y��[z�8����9t��G�t�\S�+�d2.(A��/�\��?IO����,@�����"T��tX�:��X,��sW��":�9�wT��z���+N%P��q̱�l���W���z7�y�ᢺ��[�R����U��:� �M����œ�C�pj�6aqO��I,C�ɐ�&�i^�n��'&y{�u�8n��y��n�/�G��Km.明*�I�
��-����+�z�hp�G�J�Hx
A�ј�q(�Q�.���^�3]��.��D�ι��5�Y��2 1 �F�����*��~��;悅TLa�*0�] +=)t�X���Bd��e��W�P"s�������.B�a3���i�#6�a�lc'���ƤV3��;�WKX���e�˙=ɱD��l$:AӅ���ؠ�gF���(�Ԓ��
a؏lFǬ��x	��j��9*?�0�{�=U�!�k]�~\o�7>�Ē;ǋLh�������������*�}I�Ӏ$�j�����C��Dǲ=��Y�8�o�+�5	emq=>�/�ځB5X��}:�o#��5MHuۤ d����r�@_�,������e�N8�BJm��j����ltܸ4#i�D��..;lK�"�E��ߏ�g��1�>����;����B�x��%��y��� �O8t>�U\w��V�%��K����V�6'Sf��� -��Ĉ�.��1A�A�[>�]*b^����C���46��d%��/ԄM8�{ܦ�]� c���Ƴ�sȞ�[I����V{��)���Ĳ���!�N̧����e�/�H�d�6y�U����]K��)L�G~�q�5�s8yS�@n��:�bZ���5<���:{����қ*�<�e��xRoqѴ9���o��W�s	�����jGEC�
L��Y��ʴ�H�0�KÇ|�� _�9YM,��\��Y��KZM:ם~�ҵ ��|�'\�U'3��$��o�B����R�H��`�T%�	 ^�w�C�Tq;��8�G_���Ѧ/�Kڕ{�H���+����S�9]���&���Q�}��p��q�A�%���l�Kn���P�A�Rw.�������4��u�>u|m�����?Av �!���ߛZ���s��SJR��/|��	[� ��<�剻�wJ֩�=)3Ҷ�]Ux��c=E�$��Ø��������'B�Ln@�v��N���o8Mt5�M�j����!9C�I�h;�\Ȣ�L�l�Y]�2��
���ݴ�����nT�	�Yub<P�1��Z�M��>Qܗ�JѶ��@3��ʃ�-x-ss���u�h��!����>}r�S����^6$]�?i���|��,.���qc�Tȉ9IC����< �?�oI	�S�L`�������Χ�u���{�%��zH)InM@��? �(���kS�Ӽ̚E�F��E'�	�g������>dc�w�M�x����N
��*�l�p�i'�c�<�;/��˜��碝�׶�ɇU��&ͦ�*�v���>�2`���,jr���*��Ke��������ۭ�y6jYX�Bu��T9���yP1y��w!��vЬ��V�c����r1}�&��Խ<�ޮ��R������p�r��������D62g���`9�פ��sƷ����9h��.2eVF�9��48�%(n(d����u���D�Eu�O�\D}�gfE�H���߭�s:G7	(s�6�RN�>T�f%Ht��§q�y�@P�?�H��*\^<�c��ޖ�/�cW��.hc����z6�\69F�m3Fc9�.oD $S~g��.����-)���wG��FqwU�Ep|�%Д�땤=W�A���I֬1=��?Y��iH`pЦI'8���f9�1J�WE��Q�o��=5�H�"@��%��K^��;\k��~������Q�%��G�V�&�׹�;?z��$���6b%ɍ�B5X��P�l.^@F����8��uSl����dj��@��+�Dk�=4Rita�`��|��Chqݲ�U�'j�X�����!��x~�ӕ�-��ކ3�PXÐX�t5��k緙�V���������=	5����j|Jkd:�!�,���3�~nY��M.@�ȧ�C��xwO5|[�~ef�^zR����㣇Z��{Q�[c>8���+6c04 V�f�n�yL���Vl��b���C!���L�%�- �7W:������܉���m2L���u �㲌�|����q9Kf�[�N���4����jq1��q��k�1Zd�cM�mn����\�Yg:��w�`�j�<R�7V��SZT� ����!�����{`$�l	�N�)�*øm266��+.�����=�q�б�7�q����h�\9�s���p����W� &� gq��i���g;�����	ϩ��h(��|���G�r�$�UV���'LGyE��_[	��ۧ�n��P��^��&�F��o�,��MzVb:�鸳�{b�t����]H�C��]8z��6�� zɾ�v�sI�h�Yׯm<�<�TB�`9n���t���; 7��9��-ݍ�
G;�ݓ�xh��t�g�Spo���G(�6��顱�d��ʽ�����D�&'�v�x8�ltC��R� ����������K������	O�&��q��c���Ջ�;�l�G�0l�i�{�=��t�=��i,'6�滙��`_��ج�W����m��\�^�&�E$@���K F�' ���Y������]�E`��DDM�cu�ԧ��+I���T�����CW�gR�I�M�w �ۢ	2!�e�U4G2i���Kd�����u* V��[ݘ�3=��)�',�A�[
����y\p ����%!��-�4�Rإ�Q���͋�`���r��3�}kZp��	���^%�Lt�H7�b��yaa x���L8|����|��E�/W��ͼq|g���YQ��#�)H��j-<��O�1�)��t�lo�ssCJ%)���D"�*Ac�H���* ����?�fk��*�v��a�'��8`v5�dF�f�7o��8"�����gO3M;b�J��n^씧U���\X�ڊO���m�/郉U.;0x��l�	9�ɤ,!���z���_�A��y߽��3$�Ђ�����8����<3�i�t�S��zv\��?�>v;Uw*Y��Lȫ�c�4? �A��R��m"d��i�ޡ��}�9����	3e�ٝ���(�Ir=����-OB�ش-�|C�!-�J<�{wi�)NH��.FE�>k�&昐���%.��3yYO�a4fxh��t���0M�βZ3����ڟ[���h!����P�:L@S�����n���a�T�8~����K���[��-��)]���v�vFDћ4�I��yאj)��D�*k��0��p�JN���K�I�"�|Io�p���N�N.�4`S�_L�P�Ni����;�>u�E�՛pM�r�� �FL�g�{�@���"�������:���kdK(~�GZ/�@kТ����z��a�	[��w֔8E�G�HI[��?鱐F�aSS��Ai!�>�#����gN���/y�Vq9͑�v�L�cm�� {��8�ޑ+=�]d"�oZ1��4v��V��%=�'ý����x�>+�|����d�W�9p���ڇ���T.��`ۇdW�>`Q��v��0Wɫ*���O�l�� O��Ͷ��U�3�Y3��&��W�ŵ���N`I��"�H9�ۅ���M��_���4�SY%�`ϐ�$@&hך����Q��iΖ���,,�!Av��b`C?ӆ���;WDȼZ�����N����W�LF�J1��>�EVc�o8�6i� $X3�akp������DŶ����������m�.�g��$m���fH�^e�Y�I|��p��5e�}Mz�̵����W.ʓ��4�0E�^����ѴL *�3����x��_ٻ!Ġ.�-r?!\�	v��"4�\�w}��ݿ@�5!�Dxt���/U�T��ɪ���.��p���jC �㭋x���h�^UC��d=a�Y2"S�a��1���!����D�9�0�Y�'�b�B��*��p��ulK����d_��\_!����mnי����Z�O�35��<D�GG�pHZ�N�ۭ�����P�^�W���PMpLĩ�P������&p��8J�HQ��v-��?c��c���.�N�����ZH�NglMQ��ނ�D�����)ȹZ3d���Ώ��jcH��,���̢˵p9Z
��9m�1�[k�R�0)�f�zϬe�3�EK�������m�AH�Y}u�X��Ce�ī�S�K�]9�sw�<�_}�4*��>	�p�YS_u�W�qn�u�j�J��Y^�n��߳-�:���j6D<�[|�$�aƹVu��,�H�H���9f�Vݳ|U�؆��e��[�b�0$Y2��`�\0Ms�F����=�2oD�TB?I&]�U�"G?kj	�v����,%����A-8���f��vl�ms��U� H�*��d�S�� �֧���ۏX���V�Մɥ
ޚ�&��e?v{��\ަQ���̐��+S���)|�6�#x�Y���܊?O�4 ��"F����{�qP�"q'R������ӊ@��fϪL�z�x��U��X���YfHT�C9;�Oo����$qf�CIn#��t�������Y��І�8L�!z��wo���-���c`!���Ix[x�����D�����F;x�u4ɵ����H�췱w�L�h���.�h8,���թq&���f��r�5�r*�p(ے���u�ɡ��m��Zl1��|�Հ����p���\�w{���"wM�0Θ��h�`̛aO���:�"�m�n3�&�eٟ�$Ԋ��"^c�q�[�"�D�$o���`�͞���[pd�ˆ����\th�A�蛈�T�@���IԿ��zߕ��М���c�zA^L���l�v��2�R�ּ����3q�6n������~�������`���ib�7�ei?ܛ��l�G�Ӂd�6���i�*u]J��(�5�p-�6�9����s�	_��S�k^�{B��s�E���%��u��0I�d�<o�"����n�ڢͼ��%)f�)*� �� �.�:w�IuN(�u.�`��ʧF�Α��dB_�5�i�����$L�g!Dg�}Fa�H��!^u�H��aĤj��z�U�{� ��Y���n��7�<���KZ�?�~=�����Jy2J]�;�3�Ր��E�Нn\Y��t����9�V�l��{y�`���T���To]U�USt�A5�}%w�9P���jT�� w�B��:٘c�d�ryc�$ʯA�R�����:;���[�'���.���rJ�"<����C�ȩb��q{��u��&�v��'�^ 6�ph�Ȃsg�f�ej
�e��z���cBkTȾ����'m��_�Հ3��қV�<uI���؇
�-�X�ysu�J��^@޽Wfc�oI`]���d���d!��	�4q!1�v�a�c�㿬�,��כ����ӆ�m�E���M>Z/�]DW�D��0�r��V��� =k����2��
U X0��~pm��h���t�5X�c�+��]b�Ͳ���c���ꫳ��a�|3�t��c.������]�i�^�u�c��e�I�>>`/c3���oP�}1����u�<Wf��~���uaw��аm���]�]�W3>��!���-�F�Z�`��$<�vq�a�Z3���Yy��P8�D�������^I��dc��m��(��TN<6��t���m�&Rʂ_�;������VvH=�(�-�l�J){ܞ͑z'�CI���(-F4�M�6};$; �(k���;U�A�d	�9����q�Z�V�k���� ���+�U:�Wˤ}�8��Q©�f�W�]�V5#!�2J'h���O��icr�/��*�~ExhXC�
�N�X2w�R���,�&u��ؽ����(0
��o?E��.;�;���IU�:v��B�I���ݣ�i��S�Q�<p��1�HH8&b��ew-H�
�� ��"��$��ܡ՗3%i*,�uB�l�dZ<ɼ2�r�������-Pn�S#�j�J"�se�Gz��,��&� �-�n�! ��w$_�=1��t\|�e~'f���c�Tg���� � ��Y�p�G�0w��t`b�M}q�Ÿ�s@E�8�-�k-����0�"�����۸	��^�"�kG�l@�����ܑx�$�>���ʦ�D�=�z��k�=tΟ�[���I�p�z�8�l�u�a�#U��2��/��C��G�O:���p��~��UM��,I�Ww�d���[�_�R�z�M:�:U�F(�p�E���h��Z�T���zmr3��[ V%�x��8)s����nH ���_�XV� �tFIS&�Я�K-��Ɲ ���&����ױ���-��FP�,���=��S���uw��`A|��5���dr���K����{Kv�3Ww"R�}�§�Ď��=o�2�Oz���G�[T���o��^)��l%��=�0y'����h)x�~���Wߥ��G�)��X̥�J�QJY0'2��_L��{/�~Y�j�t�#����*�H|}a�#�`�D	��Ӧ� �q�S��bFF��A�x�?s-������EJ��[Gݡ�����4��|j3�7�t�+7U ���[S�$����wˌ�;L+�F3=4��K��J��kd(�w�������/$څUT;�۸"��Rʔ@񑰄�7�Я����y��j����x�:x�Z�iN�q4�<��02�/�L�8�&̈�d��L�;uO����cQ�c;�M�b�4�
k�`r1԰�u���Z�VW� e�6�*w�#��
w�>qs%Ct�	�٦���N���<�Y64mu�++P��p���b<��}cBZ��N4e�7�� ��&���ų9���EA���c��iE/�C�����d��_H�p��t��¸;U��Ȣ2�`ORǾ�==������9���2�f54��Ń��N|.�n�Mu���1�r���yzE�+�GD��k��	����9��A>����8^� -8?�k�f��� ��^�(�FU����_� �R���5���}H��ݵ���G��CĲ��ǣ
�3#t`������� ׂ�%g�]��%�#)���GV�*&`�Y�xT���|����������کO�>X����Nm=ݎ L��b�F�Eo�ks��ҒI�M?(:T��g�?6s��6����7��J����铒1�R[,�}�3:L8�t�F#K��m�b�tzN5v�I�T2�Ų�	\��Nȼj�O��_���0�e-�я���K $iScM01���H
�!X�����A����s*x�Uwz}��"���5h=����3��th�'�2UO�6���k���Q��Ε�Vh1l�7�qS��7>��QSI&,#�^�"�
�����&�rճ�����)_]#f�ɶd�
�д62��n�ߡo�>�&3N�
��I�,���:�=��r��DҨ���$y�Ez�\qE���&\�Z���--?O����]�FgQ(��tdf��M�2��,�0�^v���g�x%��m
�~X,�Z��M�����ex���#u��1&��&(X{�֡���`�F�
v;�9�YVmQ�/H�C�o��x�kQG�{|3s�\����c����F0׭��\���F$'H*#*3b�<����=�12p��,������J���x�cp�ݜӱ�oł���VX���ph�����TS�����&�*8����7�	�_�D>xD� ��-�
g��,���R$����2��dRL�o��Y�EN���K/�ֻ}��K�u�~U}�2*o��ԑ�K��v�� !$h��+?,�(�Y����0�?;�U} z{�GN��������y��+dխF@��RՋ��}-<��=��b7d/g�Q\(:����$�#	�-�c���s}F�|1��'ↂ
��g�� ��)�؊��>���ة�.C�
x*�+)rO P~�H6L�"ҝ��*Q�lW��u iUr���b<
��k��q'!�JF�J�vyU�(�YK��6�	Db���n��,=�5��=��5H���4:��je�P
̵̜Q�zA����b��.=5�O�����'�m����]�o{�*X\8�c��k��H�[	�*x�т��QU��$)����ic,��H��X��H���PV����/eW����pcY�V�@����u(�M�].��פ�W<z&��1��Vo$ǋy�wӌ��X"6ǿ +=�1h.9�uk�U�+���ˤ��
[�g�(��A#B�z����c�|�lZ~`+�^�Q{�J�u����3�c;^�H�;�xZ�W���(@C����c2ū����]}R��+�c�q�WW)�R�jc7>��Gg�����Tϧ��n�4��х��&%i����W��;�~�AAg���R�l�a�[�D��H��H� w	��C�`�2��������Z.�F�A�{�4��C��糣���*���(J!�v�<rէ���h�B��٪V���Y~e�4�,��|@�����_X��7C9J�&��q�ƚ��)&O���n���+�˴;S(-H�/�ʓky��;X`|6ɍb�[��lX[bt�;vC��9��.Wj���g��=>������h���a��)n�N�>l�(e����a�\oL�N��F�֓E�1J�~��桄���_~s����eζ���s�� [}��^봊���l`qFnZ4�؅�m_(�)��c�R9�w����Y�����$!��#!�wI7Mf�N��jY��Ǥþ�l>0ߥ ��U �R%��n0��2@&>7|b��ķ�>B�9ӡfikl	�yoe}�&��"�3T1"��t����<��F�0�򺤐K8T@mH�s�����u������W-�¥�a-���@��'1��(��C����|N"�g��f��x�����$�u�*��Vp�8X�#�̢jO����6��z3p#=�a�c��H3�

�f$��*���n���N:zK���eȌ�*`�xO�Oi�A.l��@{q�)]&�^�����!~��.=�5��|)�B4E4,���s3����� N,���-�7�)O0g(��t4�?��<���+P"��}�&���`��'^��{�j�%�t�.p������c�5�,�]�)�D�`��f�YucA?�8nto1�6l�T����h%�a_�JV�X�*F7�B�5*��ͿEZ��!�J3��x�&�R�����ܖɔ��N��J<kz3��[,c�0�/�[��O�։�l\n�K�Y�Kl��!�]�Œt6����e`��dM���e��@��ʻ~h�I�s��}�H�y�5e���ڊk�Y��07�j���$�Ȍ�g)�d��|��/B쾯*��z3$ɭ���/�I���������?�'Pk������7���+��H�h����vj�a#��;����Ư	�}���T�U�t��n9:˅&"�P�����r_�p1+�e}^�0��������ɗ:�%s�!���v�J�S�2% �CG$��Ռ��U;X��)� �C��5V/�7������/AY���F/��̄��n��y���g��{:�:09�#���2 �`\
 ��F�[q���6<_�#�͵>\���"�8����،,�=G�=�{J�#!�Q�ݤE���k��L	#�{�[��.oO�`F�ݵ����QT�>l
�롥�����g��
�"^���Q��d��ƺjpn�M���t�q��ƽ0T���r oc�e��"��xRlS	8�k�ǈ��L�pv�0K�(�1��ؼ���s{��9 �t�LԀM���Q#Jce�����1���s�'e�u����.�yQI��]H>�M~����jݞ(�!�(hi:���q2���I��-'�ol��s��{j�����S����l	�e a�^}���4��-ܟ��u���0� Ĵ�k��s]=�C	�'�s�����yVq6;�*~�3MHl����C�8�����/T�&�wj���co��o�i���/����2)�u��,��	��^���9�<bdʜu- R��:��vO�f���KH�H��w�5>;)�#��B��=�r�w�7d�X�����Nv�Pϩ��i�J��0{���ŕ�T<�lt�(�sf�8Ʌe헱5ǐɀR�>&�{�e�����G���.]�K����l\�"��w3N��ź�VN��H�H��\/O���wp��{��(=������ĳ[4
�'�uQ!!G�A�(tC��U�ˏSK�j��G@݋���6s�S��n�O��IHR^Kj�ߖ%aƨ"yն�M�J���U�W��ɭ3�y��룯p;�.�]랹h�+�e"a�D� ½S�v���A�ᗘ�{�]/�̜�@zt�Oi�E�s8U1`|�N�[���K�PD�����c\Kn�Z�r`��܆(�gb:_6�M�b��}�RV���XS���r'�
ۭf�=�o=��/�O�(fr&�x������ugqɊKLғ?�B<#�kP�
?�6"Ҭ�`� �!g�=J#:Ϝ61]�X����S=�kg��C��m��dQ��I,q-��p=	���㛌�t���(uHAǉ޲L곖�����y�f�/���t9u��ߜ�Q�?F������2�?]|�c+�n��(v�L�h�1a�㺝�^61��9�P]O����_���j]ԛ���!8 �w�V�T�����cX>?�a�!b����_�=�ì�Kٰ���qy����Z�gnx��3tEj?À?�3I()NGD��ʝ<�C�����O�?Dp�E%ze�X�ݚ�\61�G�.#)�{j�`3 �:�_�� �U<^�)^?֜?]�چR���?����.��׏�7L1�';�"�U�p��3��H�C�4�Yn��]0����i����=���W��k����3߱��"��������Ҝ�q�Gj�*+��=Q��F�p2�l.���Q�=^!A�r�[�W�D1��*�u���|��TZĀ����b��Pe��`u�NH��H<��	+���]s�̂��j��*��Tۼ6*����oU,�����9K=�M'wa���0��gǃ_��>m��b�9F�nl�F�*��'��S&��73Qq����݉���˥��`p3T���:<���6�hp�~���M_��n&b�N��̰�|>��k:1V|�O� �Wc^;�񡫺����df��R7Aa2����L��i�����J!�m�N�К���V��N�n�9t�Mխ."���d�T.�
@�����N���	ki�����΃�Ԣ ��T>��ˑL�4{��oN���Vo�h����ݯ�,o�����e� :-�"�b�#�ƺդ��_ok�lR��9��G��������5����Bښ�E���͚gr��}/t�؞�Ij�n�P�͵Xlx�E�0���L��%�c��)��̤�tX�	�\�'9`!��mL�N�:U�j�6�YoR匱�4��-Oj�."4��r�!���+]����J���_��f�6�!i��`�5��j�G�f�N�3�#�b�a�%�t�帖�7�>���m�R��h�`?V� O| �s�JoD�U鮄�A�UN��POA������04D��Z~3:���t���:MX�����DJ١����;A�}Y�Ӻ���Û.��lK��2����!�����E9�502�����I3|�
8Na�5�65Š2����X�q��q|�\��J
F�2I�/l�?an��#�9ƣ8$a�Qw�e7&kS��<O9�p�e���ؖO�΁@4�Z�X3%Ӓ�c{��,�Z���8aM��[LRY�&���Qq���"K O�Ѡ�$�Vm��JÐ�	��fp`|�%��%��g�y�+����O.�ҁ����y�i����������w�����ڢ�xUa�A�N���b�����V6�q�`���?רl����wm�αnQ���>7���B���ڷ������Af^jJ^8T/x��=���3�Ѽ *���M�6=� dxs�G�K�E^��@�ȝ��C�!��2�oP���|,_S����6����r�)�hY�#�ta)� 9u���b�H��'�`q������b� ��l����`?'��-G��E�����N(;��rj{#���w*
�]���F�[�d��N��2������yP�H";u���V��^{����gqM��,d�{����}c�F8,���C��)��h,�,%m'�K�j��1�m�V�����o�E��PJi��ܞ� �#���JE�i≟�xr�'I�tf�4�5�4pM��V�Z�i[Ѭ�]1-�?<ٛO����Ć2w|�0�ĒEu3�V�C��:�1T�����	w��йq�N����ΐ0-�_����R�)+���ױ2�0��@�:A�H����Xk����Io� ��qT���O�����F
���Ѐ�c��=��q�>kS��m,�
6r�`��Ā��1EOwad�2Cv�'��k��wq��E��KbJ%I�'M17��v:��9	��X	�!>.lH��.���v�it@(ژ�Bّ�'����D�3���ؓ�H���?%����Ɋ~���,�5Į��L�H*��?=(���/�T&8��o<y���Ӱ�/�&X��ο�M�pn'Lfp�ú/���ug�T.�r�j� ��+F��f��?,�ˁ E��Y�Z?F	m������-p��Q� ���jS����Xz��z�xLܨx+�J�-J"`��3���"��H�����4Ѝ=V�6���=�E�eH��6׊9��a��)���e~�!���ň�l��~P���m���0��w�����5�zѠhԆ+H�v�%���^��X���G?����))���+n72u��V�E�g%j^O����R��ЃD.U�Dh�3 "�Rn�s���ٳd����3��w\�p�.��0e$�ںS$�&�4-f>	ڵ�eM�EY0ɣ\�&͢�t.�_��;G����K���^i�;��^o������Ϥ�H�6b{{��4�&LL�O��$����c{N{�J���=�G��+�h�f�<���7���C��ó�5�Xaɉz��ǥkeP�j#�3ӿê�޾l�5{�P���<�w75a)�W/�Ҷ��`��fӀ������NX�ۢZ�K[Us����]�4�g� L����֭VT���o�|���\��u5��H(�7�ł�m3>�?pBM2mť�R#P�a5�:�?5��_�B�o��5*5�*�P�@s��75Spv|6kt��q��@A,;vX	��5�}�h�v��$Lw,£���kj\���ӕ# ��j7�+���eL�%��o�p�����QC�^q�)�~�e�<�Z��ip��V�	~|k�tG�l���S{��Af�w{�~�o����s]�ҽ�ʐ�-&��Fv?|'�<��,�o�D��e���q�_y���왡��֬�yy����D؂�#?	R֫l'xlL�&��c���@�o�^a���ѧ_im�6�D�}#�:����Ed��SV0od���ժ+�t�F�%,`|F��J��_Hje�&&Ŕ�� �PŇTd�� ��[�2������'�yY#K\@�E�Xj���X���L4��yܶ�1�H��`�f�D�����Ȥ^??/Y%p����5<�}�(�4-"dv���vt���;mp�+U�ۅ~�����~CH��0���*a�2ӡ���Wc w����|Qg��# ���c��]�����F���@b�y=�璉�jy&[m�#H��d�;���Ќk�D�e��M�$d����Q�8��%�-��>�Uw�y�M�㟃RY�VT�pMfw]�R.$���p�WF�W�
�hՈ{^ڠ�"�N�%���~S���<6Z�:aR?rnm�B�YAM��������
�W;t�Dc���'�f��mg~��{����~�w�8٣4��6��R��ʭ-3��"�U� N�`Q�ƙ�ٙk�`x*y׿�.�^A�m5��^��O�ەg,��{m���!�q1�UJ�Y�����q:����d���vՖ�.���'쉣�|52�'��++����{G�,��Ae�ә�E��jC�~�pyk��T�3�%����Q�y����1z!�bc'�ts��R�!K����I� �+cF�4O�RT�����,p��;����!�n	��k
	�V?K�f��#E�#\0��>�σ:7��U=uzd�!�"���|�V ��F��+�Z�/: N8�=E��d!TVHP�����_�f�5��4�U$X����dU	?!նX/�W���2���V��q),�dA�m
�}m�C2S:�d��> � 3�aU�fFnv����][��4��̎���>�s��~������M�<����Od3\%�묵40ޫ��4p��Oٰ�����<Z��.EZi�%�b�,�."�\�[�vn)��� s���N_h�����h0b�J?P�<��4�����z8p�]K�v۰$G����Н��ҷdZ�C��ϭ������T'S�'���m+��i̫WQ��f7��^`"�F�*����RȮJq"޾f���Z@�.}�#��%�h�a�y��L�U�T9�������n��t������/�1�!��iC��`d��l�,tR�W�o��-J�E�pW��T����p	|_���,�͒/��mz<a�Q���!�Z�ΫK��/��� Ms�V��R��iXl³���N���7Ouօ��������K�ٿ7m�t~���6B�$��oM���y��;��a�(�_�k �K7�-�7K[ߍ��p
21����Q,�(x�]<�p�S'��w�R�%�W�(|Lj	�*�$B�w���q�AcS���4��}���3z�O}Eyw4ת�v.i�a����K���5;!��^���8EPZ���׏����R>c��@�^~�-![�v�^�uu�qi��k&�|�I�)X���]��5q�=
"�L,2�p,q8�O��"!��� �n���Kr�p�����&U���
�Ŀ��0t���>�g�_����|թy��:��� %R�6��|���#�Q��*BesƕԐ���<�#��ʧ�n=m��L�8��9-���%kP�����3@�Cf��pC�ֲ[�����w]p�M)�\&���(�Ø)�d�v@%B��@��Fұ=}�����7�j2�7P��%����.�-��ALĨ%}����L��)���S��"r�O�ϜV�:�Y���/�f?糱�C��۹�a|��`�E ӶI;սD<o&���X�0yߢ��hѤ�E��Uˮ�Ǿ��y�W:,"n���� Ģ�Q����&����h(TZ�X��'�s�6aK�B����p^��U^���_n��u�{h��:�eF�"���uC���3���Whr���e�)��\��E.�+��kè�V�D�U�o!� ����9"y���T���Ю��ٞ�Z�L��T{�a<��J�G����� ��kI��#�edC[��A�"?�0�Ql\Ί}
iC�s�Vʔ�Trl�V7��$Km8�4��\x먊fޞ~�6.(1�� �?Α/J�z��L��)�fVj[���d~Qt��&�d(@~�7ý���W@���΄PQ�K�g1l���ZU�+�F���h���LSѐiN�J��-�|���K��_b|N��'_w�?�}Xe��	���e��8�ܣ|.ӄ����z��dh��
g��\j���:�DU�_�:;G9"���$8�CN���2�B�9T�<��JČ�l�q��d�J��&����$��y�n�8��J>O�Б�f�ͬ��z�6J/A� �STs[�w�F�ܻ}�.4_�>ib�q�=�������U�5gZ�ƴ�P��?Q��Ss�B��ڻ�g#�!��rG��V�'����װ��eH��P�x���7��6�Ѕ_�u!NKU�s��n�g�vf;1/o��K٠��#X�Y��P<����*C�T�{�Ls�#ؾe#J�$>:`���1�\5���`~(�\B)cZ#A���8F�>�i�Y:�R[��d��p�5qi����U�H��&�emZ��f�"-i�������z�	�@4����vn����̦J��X�UO�
����f�˸D�Z�k�O��L�r�V#�<Q���2�¯`�^�?�)����Bb�m�e2*�I`b��j�а���S�D*J�X����W/Z�?y��j<�䛻�RuI�IƹSZ[�X���R7"[�z�#,vE�-���z,�o�� �lR���Mg;������C�Z��2�7��:���&�ݐ�Rm��W�^-��Խ�H���9��璶��X�*g<�s]�~/I>�qZ"�ƽx�<��/�˕S��s���:F��^�=��|$q��;� y�e�� �^�6��l���9At���ɨ�� �#�HX;�G~��B�v{e�~�5��a}������!1���0~�:�y�8"���Z�O�ǁ=:vD�F��*?�F���"��$�G�)3?�-h�S�'���-�������V<~ȇ1/��o߸�N�������dq2����G��9�,��B&Z�K�����Y�>SpqF���͘oy��wb�h=U��3Q�-4:�Ey3�s
���"�Nt��\6�g�w~xH�^a�/�����8%����.�::>{t>Z[�ņ�0�!�Ƕ��~r����Hƀ)g��k�!t<�x0[;�g
�K��4;�T�+m��ڙ�w4�0Z����Id�=KvR�r0#r����э7]G�0� ��0�kW��i��L9�;�Vu���s�̂f���<Q�����F$�ր&lp�q���q͕�����lZnk1i��XQ��߱����t������\�nA�gr:`^�w`l>��7հ>� ��l��o_��%�ٲ]���e�%H:�_�
�[�L�C�q��u�?���{.@Aɜ��&\
�v��;�]�6�s�P}=Mm�l��5k�+M�v԰9-���3�����t1��(R�+�$	:sd^�]l�����I3�O�I^S�')L?	$�࿳�h5A�k.%��u��ӽm��w/��XA��8��K�^VimziE�݊+�h���^Z"̞v
f�ӕ���?�k�	3,���Ĕ<�C���J�f8ov��L*�/��Y�������4W��"����������K���ԫݾ)��t^GA�ᙩ]Go�A�ߎ�M"r����_M��ul!W{Z0�z���B�!�D��[C �B����&.~y�Ӱ�j����{L���\H�PĐ���剅 �H?�yJ�^��|�$�����2wfۙ+q�I���oggϮc֓N��|_=�|�זu��(2-���h�b�O�љ��C���n��3��_�����e|k0ڠ�f��=h�uL��Ԍ"6�:ԕq����d�8��F��3=��aT$�=�Cu����?�ɍ��V�sQ��k1��t��z��t�A����[zt.h��iޭ;�МLܔ����ֱ[ijI3��yߥw��D��GC�&1���-ҭ&3�nC,�B2����$q��31ɢm�K�ǣ5�h0kW��R�H8~X�'���{A㞻Mk��kH�T �xt��G�6���vT �h?����0�$�b�I.���٘�R}�KC��g<�E�%���#�i)�H�lO�Wz��k��8Ⱥ&�3�5��j�����e��Q=oz-����}��	Nu��!AZ�����i�����v� �<kd��Gj�%I�O�!��U�����oD��|�\xы�wة`�'���':3WG�!E��KYh��7���`��}'�����Q�?�${��aw-�+�����\d���n�(?�qf�����B��Ě��X����L0�{t|Y�����`�X���fDHe���`���i�f����ַ\��k��Ə�k�x�)�N���q2w���Q���ba�A�d���q+�P�j�J� �c�b�A& � }�u�#DG�b&���/���������:����Xȵچ���'��)[��9�آ�%�1�O���۸HZ�Մ��������O��1Z����T!M��⻗�n8�D$�T�8��`���Fe8�I�|9(6-�
"�G�C"V 2��	![�=��~0{ϲ�ݢ�]�Ns��೥��s�A�7*x��
�ZAkk�AǤ�x�����/b>3�`�Y��P�!�g�%�8Vr�I�4\�	�X����(�!<h�z��o�'�"��*vDݳN�D�5���vv�h���[��Go�=��'�����0bH��H�G�szzwL��5u�dBR`�5}��ךI�A�f���d.�i:��*iz��>7��� eAC���?��~;p��`��Ԫ.�8�ڢѫ5�Y��4�^
{��r�Z֐�