��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQ�k��s�#��ݎ�4Jh�}������!2����s���kW�YCu��ߥ� q��j3��:��ʥ�C0�S�m�lf@q����.{�.��Wgۋ���ʓ2v��K�U�@����vF63q�^�6��\��-l��P|<��K��S���]VL������h7����_���Z-�:K�ó/�-M�fX���I�S@�F�R��b��F�\��Ǜ��`��dS�L½Wǳ�/y�nV��A�Z>y��k(�<�W��^8���W��;�u)u]'��̱&�6��*XV�����2VB�98%'|��(H�%�	��9N�T�1Z��QHJ�T�a/���,,IǼw��l����=��B�&S����I�<4�@#U	8n�j�n}l��޼��櫐h�G��R?�x��i�ҕ�$Gc* F��%<	#c�b��M������_��{nГ۲�� �C�۠~��$���Tp'2�՝��Z�Ō��9������U�_����H�
�ȂQ����}���A��~%�*r�/T�"����4��}N(�t	���r�X��y�#�<�`�I�k��Y@�
rA����Z`s_� lc�O7��WcY��ö`ă���|�1�b؎�Z�	����km����3×Wh{��l��o���C(hEII ��-:�2v1�}�$�4��VY=*8����G3�&���������K|��ngG�S�)�|�t�zn�ɓ?n�L���99��w��?���䇏~��=�r�&'s����}<}k�	�e��*��<s�l,�J��3�8��0�o�v�m���:w��Wt�~�	]�*16���V�0!�<�=@v�����s�3yx��T�X�a�S�{��Z�HL)�JeT�D�sr��n��k��@�Ꞗ�I��]�IpC}[df����������OkY�O{ɛ���H���4���%�:0�c��^9�}���^)��&�qo��D
�hVlkl�X+Q���� �T�>�q΁�Z%%�&�a9;"�V�0�����c	60 ��Iɯ���-[��7С6�Q�R��j�r� ���'�)3T�y�̘���5`���x(f l�P	"S�Z %�`� ��z�>�:d��~�����*��c��y�u!U����!���0�HC{�ķԬ�`Fڲ�(F%mh�>�(�o9�8�tì���U�����ql?��gXP���� 1�[ګO����i���c��Z����تIU��e��Vo��"a�%F۰9ȗK�a1�*t�p���{㚫@)�Կ�Cx�mY5Ts�̻��P�����oQ��C���)���S��PBC� O(�R�T�di�B{��9�Q� ��G��7���cw����yɧ+�8A��lc(B�Y?5[6�l`�ÿ�V�WW;�84�k��#X�Fؒ��7�u�.A9R��{��6�S�K)��cU
#b�āL�aOt��.eL�b�PBA�]L���I�.��Y�|m-~AњSmdĕ[���=|���dYM����������n��o8o�Oڡ������k���'$i ���\��>9�+7D0�7�W�%;�~��d=�ߙ���=��������b�k�G~r"���f{���/����V����ez���i\ߝZ�C�$��VLg�?��e�����9�P�P�@u;�d�aU� �s8�l&=�����==ա��6���覽�־y'j�e��^qe��,��O�Rdd�j�� q��-(G�Y���P#-�_���X�T��d��:X\;�D��6w���	4N�#��q���L���}��]� �P�T�9L�ʿG=Y�v�r�:���p�#$���%�� 
�|���7��C����DV:�|-�z�߆2'*>��:l&J��(�&-���s���$G/_�� �ڸ%�C!����ޛm������2����(���ĨXiҡ�}��Ǆ�Ӈ3���#gTN���`AU�ɗ��%
�����b8ϯ�'2J~nxc��FܮAֹ@�0�<���$�P��e�=���*�I]�RL�BWT�?���jMt3YH���7\W�5ep��$���A�W�؁]F]���"p����1���Uzl�u����#�X��l��,��M��痽�9����,7�,�WQ%��� �j~��`���j���N�K���H�n�i�\��s,q;�-�W��o�	I���銕K�I��/'c��܌�y~}>��!��I��X=�����!�eQ?�0�Qu�Mm.������m��tF?*�&i�}/�(�-dr0=�e�_�ٸ����'�����$p��ʟ̺�-%���()d�rR�FE8��lr��͠��[���S�M�iˬ}�J��J[��e��:r��O:h�ǌ4o��M�bM�i��T�biq�a�O�3�
H���!��Ѧ�m�55�0�Q�0���~;&mV[(M5���k���0���Fɳ=%<�@dh[݅+�dp|'����U��}��J��z.b�ѳ�40"�r_;�e�Y����×�n%�-�q*a��� �M�n�/��6���㭬�۞I�
�l�]ҫ����-��|V�HCF�.�d�'Q'�d���i�h�ڕKB�q=2��Âr��*g�=9�*���r,�u�5uAB��{o��y������B��`һi�1 ������O	.\����Ds�j�\�98�<�����_�#��x����@zU�꧁IL��xL�E�?A��Ff�k�8t!�Wj����1(�.�:�p?h��9_ܓv��Q,
m������<�x�,;Б=0��
Vy��.ʝ����s��D�U>�XVu�0���n=�&&,�\��o��r�e=����H���UE౞IKƭ'JwO���N�G[���w+s�=���_��P�8�V���F���
g�ym{���;6�US������eV��d��ҢfL]�#u"!̶"ԗB�Ẍ��PAW�<ߓԩ���L��e�:��ʯF�Z%��5�0M�3?QRν:?q0��������MkBٸ:e6Ր-��f"I�mB����J��6zx`���r�(A3f,-m� હ���O����q���!n,�}+GQ�m^�)I>��_�ۊ�io���"ri��N�R���)�w�x��c��d��J{�B���B?��B�j��ǁH=�a�v�bi��bX_Amu��؀>���5�O���v.���^'���]Գen�A����Qֈ���t��3P�M�ݰ)�-�>�j�s�m���i������[���0��~��"�!��h�4��d'������U���~������$:&�vC�X?&4c�sj���FF� B�C��:N[�����mˬ=�i>�எ2W�d<����x��ߓAvV��q#����5e��C�ʎ{RY�z�m�~�?2�j%ʕ�/�?�o:zU�$0��%c �$�Gز�tK�4�|���f��Ge�ݪ�x�1�(D_�ߔ��yHX�خ/A=�z�6����y�I_��ǣb{}
n�6��ȳ�r�>-�D�%&Y���+O8���b��}�(e^y>%M��ۤ���B�G�}�+��!-�?s���)��K�Wo?�Ve�H�:��Ca�aEצ�����ES ��u���v��u� �#��T�E�!�^�Xi��5)�3��ϛ�0\M������n����tIO�0;\{������|��j]P�s�rm,�(2��y0��h�j�"�v��}�+&,�ʨ�kԎ^]����q���\��Z�e��ut���7?��&1������u7�	�wB���RJf�r����e��;�I� fN��Cv����Jo>J��w����@g��`�E;��rWh�;:����bEiGW�\*+��*����;R�S}��Ó��Ϗ��l�w|��d���R�)_�0HeM2d��uӏ�X�A�G����y}Ù��hh�ҙ�����*�,/.XN����T��-2�0B:0�v�y��Y���j�a��!�����M�Z�;�O,c���h|n*,��	];ԏ�buV�5���e ֒*�L�KK��_s
��y��e�|� ʷ�~�sUc��8Ix�\s'G�nQ�S�QA���0{W�s��nQۤa��\�Zm�n |_cMđ�a�M�m�jҝ1~�3��]Ph�[O8�p��%�g��-�(!{N�����?�ƻ`!V)K��>�_��Pw�9��E�c6k{��6�`ja���[�l�e��8�f	��coS
ӌ@��uQKR�3w�
r�]I[i O����0Z�b!�.��3�p���>X]���
y�y����az�U8�M7�A9/�B
E��1�Z� ڕy0��?��ݍ�����Nc�������g��˃~�=+��y�u����T�
о��G��@;���3����l\�O�XβT���i�՚�𹮴��.��	�"O��mV.W����c0h� ��!SxD�
!"�7���݊��;j-����Ϲ�2:Zx,(%����%�6�!�>nf���+���w �|�D�������*r� {B�����&+��3x�j�Q����k��PI��
 �������,h���UK?E�96X�kϋ�6� d��V���7݅��:?�3�̇�X���(&vO;�������m.r�c���@���Y�@W���T�L����~����,�zo���� j&���1c5+���w����E�z��������9.���.�T;?ÿo�I�ˈ������
 p(�,�gѪ)�^����!n}���37�T2������YܖQ�(VG��.��P`d�TL�:�^t�����x:���b6�"�Lk���|x�(�Aq��yÖ[�=���%����� LΖPh��T;:Û6<�qů�t�UO 
� �C���"p-����.s~�od�ʯn:�ad)7��+�ݕ	��J�@FP�q�˩4����;N��5w�x��i�.N?�l0t?�U5R'��G��4���$AS�	����ۦ��t�����tնڳ4B8���V�naI�[z �����ƏJ�3M�.���^s��YE���~���W���k+j��� ��i�1�bL���]|8��F(Y�o�@��8�����[�)6��<��b<^S Vϻ U��+��7i\��r^��گP���W��l`$�����z���Ҹ�Y�*Q�i4��5����;A�Wp܇h��ہ��R��I���`��sR���m�aD�$5�q�{ �g(<��9����{�����no�'���1'śyb=	ڱ��������������R�R�ݢ@��Z��X6�H)���0��_�� *=���N��6T�n�Qm#<o�� �+zl�/���Je-7ai��G�5[0ۑF	<^ZT9�ch�����&���>�1�Ӷ�bǛ�VDc�fw	�ݶ	H��X9G���ʔ۔�+�{A'cNp�gf"�'%�(������2Ʉ�	��~��]F�d��2�x7[Γ ������(tWfBV���A��'$-��'���ѱ�|Ɂ6-ȃ���o�n�N�&Ϝ����ȿ�*��P3-�X�<� �
dE'�z��q���DSwJ�tu)l�A��7EٿN�|�'�
I�.xPA�rZ�e�D��W_����LLUp���/\f���zѿ&��֪>�[e.CkmYq�
���4��#����@gb�D��9>�%�K�M?�SUZ�{ OS����,e�R��r�2l]J�!�l���.N��{y�3l����aY*�����U��#sd��s!?�7��:�vķ�2S�G�u�52����:C4����ЧX�R�ކ逻�p*Q;�ŚQ�G��P}�m{ir~n�#�BI�U2�ס}��f9�~��̇g`h�vɑ U��p����9tJI��U�\�ߧ����)b���MT�<;��yu�Y�@�ز8�ȿ��PLؿ���>z:|R���sRC����}��m�}��3���޻�{%������2,�-���G��6უ�Q�eH�5��?�AV�������%�d��-��kϞWJ����7\i�׭���/����:�>���ӿM��&�s���L�ruԺT:�Li�<.<t�
�לv5tD�X��OxK5�E��Btc1��s[�������R,7r3�|�,�-��wS���0���y����~�1���~�=%�_׵8uA�]M8��-�d��FU���%�Dw14-~i�3�H��]�cnL|$r�D��OKP���V��`���Y���lZtDd��kК>9A��W\�`��)9��5���\o�`��-�{3�ֳ,i8\�haJۜ�cqJ{Z��{��i%�i�\�4�����V�ep��G@]=�&[E�#6j�+�S?Y�~ח�����%$�d��a%V�W��_�|�-�I'�����Dn��AE���ъ���*��u8�gW�$?�̦L�*�ς�|�1���gA񚋢�j(�mc�!Îh�,�P!S�&g�^�M����(zD�PY�#�������ߔԏ�9�t��d'��ӿ�W�Z������v�8�h��nٚ�n|��$Q�G2�оz�����-��ō�f9Wi�-.W�v�Ę��	��J� K��덓���'�$�F��u��s�d*�pW�r�ܝ��#'7;��K��D�`;S;��H)���5;�g&�,E�f��46p�����ƭ�P5�K�C�a�c�f�5�$HW�Gy�>�V��dz'o7c�C���5�"�<���el���7�|�~���-(���$@}̔G�)��^��(-��uT0��9��uz̿���s����5��8ж=X�Yj�*]�����yh��#����W��q��5����X��t���?k#sT��������_M��$ȁנ�t���.*-�����U�Og^��~d�$;���ں�o��8�0��%�>���B����Ú�l�G��6��"��&����������ѲoB	�QG	�1@(}�w �$/�e߆+�u�4���k�?���V�e����0���f�ti��,�Ȥ�c�x~�U�q������*Z��?�P%�OT���E�9���9뿽���y�s ��h��0�祿�u��c/�vdY@�'�:5x�G�o�Rx�X��1v����w��:�{�l|��sK�DC��!��#�uK�f����p�!�y�/K݉�	��y:�c���D-��} /'+�M�"�`9�N���M�ue^lvu!Y4¿�L�6�}��PT�W;׸U|8�� ��	b��/Ll�
�2���K���@э�vB]0\�M7.|تP9:����0�R�%-����Wȋ_^�MV
�f��5�Vկn�.���:<�ڑƠ�#�|��L��"�r��M����ۣ"���KN�MIt]��[���?ߙ��Z���gg/�ǚ@���k�	�v���3 -����D���G�"�Gܤ�-�َ�E��Z�!��|�V�9C�+��g����jMAK�0?�ϣ�8L)��`u� �~��Ψ��Lq��tB�A�PS�X��-Q87�ԝ~))�O=EMN�� ��o�\償�{6a�W)�W~Q��Ѿ8b���O����~�fts��vi���a�Pb�XO��4��'�762qAϫ��.=n}���|�wqXu^�V�J���2��1Ǆ&8v{�<��.�mC�0���� �3;��c�B�,=��o�	�/�����&p\T~�e���p��s��n�|�fKT��Mgmq����ⅳx��E�/0�a�o�d�x�)�����ژ�
�V�:�����Z�~���69̂����=A��-S���r���>nrm��f�����c��<�j.lc�(R��~��+�����fе�6
��53V���T2���9X̝-���~�o��F��!A���:ԕ���o���<fs�g��4��Md����_e�hs\�nN�-�L2X��B�*�RR��Lު���3�A>{�9H�S[���50����p+Ǳ���.��)���|j&�7A����ہ?���J!Y�lk�;�D&���=[�RHz��Q�:�5V��}܅Ҿ��I�,�k|������!TO�o������6_jv���g�"�)���j��o�"���{t"��@��� ,}�*ְ��ʉJ�F�S1���n�yH��vH.]4j�P�������y�X�q��˰�YV�v�u����|��'%�>D�k����yk-�d*)$���.4�N����E!;�%f\�₈���!�zl #��}��̄�y�j�)س��/�^mHwR�?$e�H��)	)��L�׋7D�j*k�k@�*F�6{��y(
��p\m�s�0͔.m/� n��"�����FKH$��ۆ���������ߗp��
�U����Hg�ãK� Ys���ڇ*������������"�A���a���e���ɘ6
<���\藺rRH�n�L�j��-�!�c���G��q� �nw�Q��b��#	>ʕ�V���Rݱi��}Р�E��2̕J	����(��hdq����LH#%����p�5���R���M�+s۶�g�r[�>ܗ�]B�J �6�}��dn�r~������/3�_�T�G]��r���3��*Ζ���x�Rc�%<Y&� �Q��W�h1E��_����]�\�_M}F.fMn�8 �>�׫�G1R�w��̪a������g$�pa���h�/��~v/����	{_�-�]�3�bZ�ڵ�n%� �0�Yh5��7��9ms<$9��K����#vR}Hr�7"�<c�{�ē�Dd���߽ �U �bP�|��������hs�"Ƹt?;��R_&�����ÿ('�Ε��P�W* �J5��Ytc{��X�I�f�t��ROv��������K58�>��D�^(0�q �O�L�{�?�>�r%aX���]֠���w�m��h�f�����e�a(��� Qj�
)kmW; a9��o��/�g�8�t�
���(�};���I@���p��w�'��������r�����fޚ7+5��T������<FE�	�_jf���$�W���-1��G�Ѫ�N��8�H��+�u�u�K�K�6!2�� A(CYG�� �=�k$�+a���_����e�>��v�)��6���i�X�(���7a������6̽�H9�ƚ��|&�rA��;[���o�)M:�!ܪ��]�҄Y���3�$j��q��%�<r�jvց�W�3�2��i��C�P2b��)q|�oG��͛��/��C;�-��	��)� �8�J~%�V+-��Pq�������ʲ5�[DFD�!�SFA��G���� �<�����7	a���t_���(j�g�nR����9%�[��&g�z��@�&T��d��l�T�dj3Jqpp��*��
��?�{RV���C2��R V��f��j~�L1d�rVϮ-9�P�ϫ[P��'��0��%,`�?�7K����b^��f"(�9(6�J�M��1gi���6����\u�gK��Gw�G�J>�9�n��'4�a��>x���7����{��� ��u 4Y$^�IBj�&oǚ�5�K^��W����'��R�0M��͠�����ۀ鞭�b.�i��{-�`�r�$,zXB��G70��2�`|�p��DrA�1v��k#��6�:�{.5&�*�5��ҤK�Bm�������T�� ��kW�=�WH�~3�߃U�jl���+�_u�qZ��^���U��;m�vWK���̢bH�#�&�b�o���QŭR|˥�\#�G�IiW�	-Y��e:�\|0�vo�Y���;�����k㛡rmO^,T�e���~5^��lXn����^�h��-�������
+����R��g�@6��#��#|�#����w�B�x������/kt϶�u����Y�O�h)��ɕ!��z��6]e�[���#�O���;�KO8�{�%�B�Wn�^<M�з��E/�{:?-F�&w��]%R"��L�S//T���xvA�xo|\���%r��ջB^�#m@�oNmL�/E���51�͈����;~�,�5���J��a��&*�}wĠ!((��H�z�&�`a�Y�vM�ؾ�ƨ������1AՈ8W@��0C���07`��e�B{�5I&�%?K�{��#\�Ł��t�#�o�"1�<vh�0����R�*���]';�6 ]��s��1�M�>βrXG*��?=zݡ�ǒ��ã���8�w���qn�	�`�������s�R���<�����	"��Tm��_��_��X��h^ 6/��d�Y<�n�>^mf�����1�aީ�8���0(����WI6���q[/~��v=�������%t��}��O� Y�[����a\n�����if,�4��+��Nx:Zh�1���t��{��^|ҹ(���io����ps�U�����!�K���,k���v-���V�D��(�άah�*~ǲeʭ�����Y$Gd���D�5#0��R�T�g&R��I���h3�:H��/���J����Sz�&y�m�����i�j|��6���J̿����e��d0 4��<�5�xh,�!��D?���� u )����γx�cIы�9��c�����9�&h��9��"׷� 4kM)���F�޼��2%<���_����?4����4%�W�N��Z{l"܌Z�z��. `���.���fcF)ԏ�;b����+��2^CI���J����d�f��j�?pdm�ؐ���rf�&М�;b�k ��Y���3>��ߜ��2�\(M���d��e
<E_	�vW��f4?�x+��+�c�����8��=�eY��'Di�ʣa�vD<�r�*)�zZ�7�v����';��7]�O\s �9��Dj�7�4�e6*6<xV��;�2�9��?�p�������6�	�d�� !���dGF1¹� eZi;���t��m#[�EL���)^kP��l�x��������#�<�'k��C�%�S�J���(W�$##/��d���N�����M��}���z��m�KM3��,�(���.�`�%G�g�'&������?z�KYͱ�h�l-J���2��Ob�ŌX���bY�a�V�(b�a��&��y4��w�\��_ ��ǈ0���!]֜E�bq��,�-�.���W�R>~&�a��2���N��3kKH�$B�tj��:�$HU:mp����/�-��?9b�`�c��S�S�[aY�T�ո�Q
 ׮�Mf;/wW�9KA2@��XF��X�l���i�'�KO��R~�j�;�.D@��l���e_~�8�b#�D����KkO���O����]ُ���Dp���lv�fQ+�O���)��;�/����GA95� L��ZN���-��d��2�Z@cW��PL�Oke���R)���I��|����������TF�$+���M�~p�'ڛ��S]����Z��;{t�cV�޻W�~������T%~��~=N-Z�Ɋ�u�cAw�P>�.�L?bƎz�<��I,ڄ�*�d�C�$QK�E!�>_��w�_�K3����()$�5���Q����[c|:1M��Z���X�C��⸓���t��:�kM/H@ ��TG�VU�B�rG�K�D0�`&��C������gǠ����3�-�s�8!tɜ��O篠�o�cY�^0sU��ɗϗ��t�1!���L�M�Cq��r���}.���۶����(���+��/;&��s"U��D�	咬CL��Ӣ�ʤߠ�w�Es�B��ٗ}Z�����v�5l��f�d��c�\��L������8UP-�I?�~�gã�����8V����`��jc~��p���e�Ad,�:xQ��ϭZ�>���T����d�9�����S����*�o3ւf�g�o�Rn�����R�T�� ^)PẌ�dJ}i��|��qd)	%�Ggt�Ë2l|��I�%��-��ak�:��8b`m�M����0��#I��J�e��������� 3����o��XC�H�����U@~��y���C��U��U9ͺ���H���A��2j�L�y��/�u��Ԧ��b���Θ�W�Dj�.j���a���B�7y�H0g���j�a�S����<��)t�>��}��&��E��NH'�k`�w ��#��?�\H��2��pv^�L;w�eB��PRIo��S�����f��$�ފX��@�p~��|k:|-	[&�s����b�� �%���l2�'gA�-�6y�!��[Ń�{'�z�#Vl[�D6�?+nF�}P�_/ �3wd9XL�J�s.�
2��u�L��4�N����I�G�S���e �|���>�����G���XE�gP��"�:�o�/G�P�}���3LZ�����E[�{����tn��m���C����6c���;����%��h���ur�݌Ѿ��k�m�gQ��*�l~ĳq@"�>��u^�l������ު_��������TD�ʲ�\��it�H���a��F�ۉ)pÁ���mE��v��ѹT`��R���b5S��ӬR��zE�Vgjr�s7j�)�QXފ�ؒPu����C��ǂf��&�."CM ӡ��os�[r��o�
��#o���5� ���E���R�q�̤Y�d��ы
ȍ��aW�V����Չ��?E)K�mN)�Y��f#fg쩌ԍg��;�*��Ik�@��%��B���ԇ䯉kl���^��Fˀ5Y� ��K~t�{[p�G��2=��0ƣ$�]��ӱ�����ӲLMj��q |��'|.=:Sy��QYT[\m��AI4�
M���V�M��d�l��;5�����ž�o���P}��3��[88wOX��l墐^�e4lWI��b6mmە��`&cs7�K�9cl<���NJtv@ױ�!��@�񢓒#�i��
p>�ξ�����awZ"�h���:����7�j�ƶn1�ÿŀ^�}��L�lt\G�J�'GIF�8]57�V	!�����X|�����.P�j>	�Fv�20��b#�����%��p�<1��|y�;�|9([m/�t |�����*0�6�(s�[�DFoݦ��?잮�Ez���L>�{|�>[�q=�������ݛC�gUI/\�+���:_f��nhI�C��ⱔ��E�+�&�	4����D�z��������� 	k+���r�J�8�ωl@.�3�]�ݜ�^u���蝢X�-|z�*��Cu.��Ss,L��a݇�S�Ha��VV����l�&Yw��SZړ��jmq�b]/-��W~z����,�nT���3�
f��؀+e�2�D5K@����d��S:�I�]ֆ{|��i,���R�#ǿ��dd;9��4�k5�hP�^WN�I��֠��?:�<���V�*:ўZ#�TއMO-���� L8�����B�����si��;h��n�NQm�!-O �j�/&�G��iΉ�˩�?��AOcD��䓈	tQ�h��e�	����'�����}��Q���
\���ǥ{��4��Y��R�P�e^E;�4@�r��&bvcq�t���nѼWʼ��xy2<Plt���&�c�w.wnL�WTTSO��*�cJ��>m�����
ٍ���O٨������L�4���l�J�-I,*�n��p��ԥP:��q�t�wY��+���t1�`llu���}/��X����~��/��!@��l3o����;E�S���7�m��t!��*yl[�.~��m.�.EU��[��.�VS,��j�b�G�H[˫��!���M��G�&�k�ک����z�ɴ���04���l��F�`�C]g3}�]2+G<�t�z�ى
=R�.;�1��xO����#�x9�N=U�^=$�l7*��q�`*�X۬��Kp�X�)ؿ4���z�#��o7:�-��aB+����eBm�^+�A�ù�����Q�f�A���OhZ!u��-��������ٝyA�����6�d�O�8ci��T��f���*��n@8�B����� $,ɦ��j��42����&��f�k;,?8ǚ�����%��]��@�\j��@k!�#��o{M[C�ARSd���E�fwb�ڹ?Bd�h�^Ԛ�;��L\���xwr��0��e�� ��r�|�D�pJ�8vQ��Ȕ��	4�WƷ��:����ԧ%�kneBD�b�@>���p��{`=�d���?'��s�H�:�0c�7V$�RZ�h���.k�ƶZPm��2a����� ���z���������ۋ�ׯS�X\�@��8$����S���^����[��Mq��6]�8VE�Y�
	��aD�Z�E�lS[�ӈ=3���6�_u\%��6�m.���̉�@��<ϭ �<U�M� V�݅s�#�N���}���a�z���s+�zUő]�g�s@j�
zn	!�<�zS]#n2��8\=~|ʳ�&�@�xo��㢈�+�K}��r�%Z������k�3$�e��y�2�K!Yf�& ��J�ͨl��Ya#�;��;Wl�9O�Y������3��JBDV��$��z�����F�sUf�s�<Я�_}y�|[��_G��kdnɊ�[�U��,;6C��=|��1��ٱo�t��o����K3X��q;D��՜�磽+J���&�mW�dʒ��hZ���^"������UaJ���T���i������w�u�\�A4>�����I�&͂�b��bog��l�3�m�/�f�>�X�^Z��y�I�Ԩ��? ƚ���64�+�%Q���x��^F���Y�$�N��+�x����ؕ�܈��AT�\�K	����{��FU��ā���9��oڳ�P֑ڕ�N�D-������R]���1�x��jֽ@ޙs�`k��F��"1�?�%yuSb5��A5�)�DS/�j}��zF�`�(��u���.�K���(�>()4� t��c���ap�=-��d<j��Y�J��Gk�kZ>�(���]3��ϺqP^J��$t���5�s ���>�6��(X�J�U4��n�����¯(C��9�|hPݱʂVK��#�I�H�86M�?dtE�����Ȫ���<x���pu�<��	�0�t$^u�QX�G\��e��W<V�G��pm�z��I����f�r-,i�7ކ��;��-[A���=縋��6Y9�3�[.x7�-r6e����Z8_�d#�A��)�4f[�4ij�63W�I�<8d|x#�*����"��TO��vٚ�̀'�#@��g��A��*�	I�esLN�9$�w�)�"2����7 �0����$�w�A�Y���5|\���1+�i!�	-�P9cG��Kp
�g���zT_Yr������F�*5F�B�Fz_Yu���������2��8�A���+��c�Q����}+&65�z����Y��aE�1���8� Ȅ�١.ŏVHE���V�_�Vk\�Y�P��b5���;d��F�b=�nʞouC�MR[�P������"��C����h)oRn�F��� 5]8�,��k�WȪl��_PTF"����� Y�8��Ɓtz�rϔGyi�ݬ�4��>��v%�O��L0��~�K\�ԯt-��)W�����-	��\�^��ȹC੓j::m�ѭ��0~���I!�����
�m0X���흘
v�9�,[���Bn?�L7$R'�j�[(Tl~�@u�K�0���Ð�x<�M���J�r����8�ߋ���^`8����Z�P�1-�蕷5Y�6u#|�|�z��~%w�+�|���6��Ʊ����P��ݽ�k!�J:���m�Q(Gj6��S��/s�ڢ�N��(�YmϧJLn�=���ģpy����a�6��ؙ	��8Y�]#U�]d�2S�ΐ9>`Y@��)AX%~˺���ͷ�5i}K�y�y�9qpT�Qa\�qU�k5@bH�`A6t��G��_P��	�сu
ؼP���Pۭ���|�Bp;���B�0݈�#� ���a�X�sU�
��{�_�c�M�2��z��
?[c��B(Xt���[X &2��8��{��\Cl1��fـ�}�n<��9�A|�[=�%j� ��ތ�e��Q��ҁez^;�߰�mc��h5��I�@�jS�ތ��]'�����9���D����Pi�s� s^x/���	V����۾��0|`Z������+j��}'��E
���/�5�=<U]s�â�����)5
��Ę���RԹ����5����)��#lh/��Q]�.������E��"�B�| 5J�S�~�[�����A"h#�? ;��N��B��8D�Q?�����3p���Z�ȁJ˫(���b��Bq�?4��uה��� J~����ǐ��$�IV���M��5]�^}r8}��6Mܯ��������1�Q��1�-9ɢX������D�j觍�0���S�[��e�Ϻ��U~@�,˳4� �S�!X3��<�}���c���f5�`�"��і���y�L41��XА-����zƟ	�]�R{�f�Z�A�U��M<���|�Bf  \������:�Y�Q��9�����,C���$1l`�7�Q����<KV���Y����� �ȧ�ӷ5�}4�f�_�afMϸ������Q���2c�Nt��
,�N�ڟmU��n���ї��1b���S"����Xt�3�'*�಻�V�m��B@r8���no4B҅Ii_���+I+ R��M��3_eK��+N�R�w�D/�*u����NSƺz���mj��6V�n ��ge(�G�K���3*^��0#Ib��$q�C�V�Ƭdg4�Ӿ�l�:�`�P��v�c6]��*�d��t~ez�E'%n�8�L��Z?�iJV�Y.�Q��&��}�x��gԀ��R��ß՟�ѹ�Ќ��׿���w� �K.,��'U�=fǗ�%�jU~1C����8q)�ǫOwJR�Ry�6o$-;�Q����^�Ω��1���v�FN�>:����%�-�����@R��@�����f�kZZxy�T��q�2,=���Bz!���G|hW���+V����O:R���0�J����)�}W!�m?�����_j[�� ��)sR�<P	��.�n��^�� �۪��&}e������k�_f�����9��T�Kʜ�K �k�����T4�3E��nٮ�C�kt!<���*��b*BsXs�I-ߵ�):F�;��p���m�lRmJ�r�g��,����4��HA�炽�,{�n��ߏ�?��,;nc �HA3%�jrFQ�M̐!lv5��d(	wӓ	j$�)9��I/��8ќOQ���q������7l��D�ݤeu�x�#�I�pLb��RN1�=v:��)�b�����c\��8R��:*P�28Z�M㟠W���bc<�_�;��-H.i+'Ù冕��ƑX��K�� �M�ɭ�-�Qb��J��ϪiL�|^�1�8��%�mζv��xg۬��`M�k�(�(�,s�Ȉ?G�7����]Q,�t����h���]��m�F�����O*�%��~�NA�æW)8�zE�8ι�#�<d�2�K	�U������,}��vV��Ɉ�����$�HQ{���2/1k��@�ڽAU����!8u��TU�����}� �x-\d�����v�-����;�Mdj�p�SZ�%�[[�;.71��)�J�,���Q���fcn�C~xI��`$�5�`��%���,�C��Mm~�0~�]�%�IT�ka�"Ϧ�0�A��y��T�P #2��)f[����0�xv�h���SŨvԭ�s���tL��̷�y�
��%��n��N�����.���{�Y1xQ�*P+�fO�B�nEb>��Xu�����r�&�Bہ��#�tݳI�\�B�g��f
]ai� "�*K-�|u�]c������"��)k ���ߪޱB�8��K"��s�0�7��7�afӫ7��.5����N�y�寗v�p*ͅ��Zgl�ԟ':��(��t�?h�$ԫ�N6��5ؓ����T`n�����,^����ʶ)PF2�/�����jt㉰�LF���*�H�*ؽ�>��z�l]|6����Q�"O!�7��ϷD#�ݸ�|���N��K�Ì+�V@��'OkDTy�����2�;���1�,ٙ��#�	v�6c3_�.����/{�j�3���I�!o�虍�,,V��_����u�A��TF�]S-�kwA���*d�|�x�cPH��S��t�?�����d�����>, ���!�ue�^�����<z��������ap����u0^y�5I�	�:�puO=&4�!(f�S��UGܕ]�*&��D��6���R���LԴ\ƀ���Q�X�Z��b��;��M�4Q�mc�<&�V��O\7c�;�_��zJ�ns�2#
�3s���M��ӹOa������PB˵z��pd{�ʧ4f?�4���Q���ˈʪ��By@Sq����H��yBG�}�s��P�t�Kj�uZ-�������qE�H�*B��B��|�|�l��qI�Ap�Z��rh��zc��Ϳ��q��OCG�a�5��C���'a�ԧ��b����wd�b�Q��"3���Ta@��[�� q.QQ(�
f�Kd�g9L=kO��a��!�o	��M6S��a�S���!�m��V�f���[��v���H	�/�C�;1*����T���z�.�ih������%D�(����|�ǯ}��J^:s;h�O��G�U�y��ЁeI�T@�Uq9� =0���b�J��Q
Ƙ�%�~�
����ם��%m�#���@N��a������,��0�b� �{Ɇ����'�\�>%D���o��V��GS� .<K%���(s�A�z�:��׾���T���z?��kƐt� y�G���=�P#�cƀhR2+2t �@���h�ܲ���s�3����4�
��)�x���b�{�d���'��'��!��t�lk�Jx�g�N��2�a�s�ҳ�'1導:1}���i��G��Ʌ�5B</�L���s���7w�Q7�wM��l���Y����w�@���4����5�Qo�m�)�����6r��ѕ|�Ьh��*��C�'�t\�����;)�`��R�5���s����S��S�0�� 7$�G�� ��E�Ø��=���x�K����H���F�/Y�,���m�
8���)&R�E+o�iEg�@��Z�Kf�� ��<�[�k�aS!�YA�k;@�%yC@A����p�4nR Ȳ�5��.;´�3}����;<M;����S��5���f�\��m�EZ�{��u\7P�x��s�.g0-������	������©4����ua�����tn���K^v��Q|�wM_�97[��f�j�7d%�V<���9�L���*�{\�'�
k����YqP��[~��Ԙ��s:�NN��*���Q#b�{3�%�� �����[<Y$�����e�N�v��v��{����[Ma���3[X�
�@r���?ň�_S�C��s[Fj�F7c@���=�� -��{s�il[��It��q˔6�Do����"W��#S��0���t�{K����@S�S�L��}!�.��/%�E���l�YtHw��c���]+�H�Wp��@������	p��r6KYS��=i%�-�N惼U���H�Uu2:�׍�G�N�mLS<?�X@���}�#�ٿ��2�Jh��m��BK{^�#���2%��of���{N��j�Y�x�ܿ��2,"�}��m\�9���,$���L(�k��|�j���mpy�E�SJ���)�{4E*Y ����o�K;��0�b�z�(���B;Xb��A5��s�~W/��'�PB`���K��K����.�i�X:�(��ls� ����NBL^�L��Я�]p�赅��3�-������m�=���՝�Oy�I��7߄��=�?탮���#������t��CD�l5�n�`�|I��Dq�.��En���x�s��^�
.�>��Fk�&iCU�o�c�1%���i�3k�P9 LímSkq��.l!-A$jE�p��:C�����,���>G��Á	a3���}�YeI��P۾��:�N	�L��>%������r��#��9_�Ow�"Y�
��;),��Q��2��ޱ�����D��Ӆ�لO�:�G��r�&�&U[���
Ԇ|����Dx�hh��吙��]Vd0p��J�-Fz=Z��k.=�N`N��$�XJȼ�p��l��`=�S�4�cʼ�A޿0]�1�E�5�ȸ�dB�ߡp����pRڈ�.ĉ�%q,p�%d00������"��?	|ǁ�����I+š�N��<��pJto�����z��5f�,���\Qr�K�镴�D۪�)M��RrU=�$=h2�>
3w�,i��)tT�Ǌz�Ӳ���6\�󒯴�8���O ���6-��+����3��a�t-F�Q˷YϷ�ɛZ����5������)���3993Kt�D���L���)�i�g͛��������e���Q`ۈC�FsGaa"�V�#Ǽх���T��v@�u�GȧQ���������E��1i�S�Ls(��%}l����m�!ˉ�v����jY�Ѷ����)=ý"��v�"������J���S��C�F]ٷ��-�p���gS	b����A4sAXH/��W~]����ӏ����p>�i(c2:l�z���X"G+���m6m[�*D���v8_-}�=�@,�2��ZZG�R����d7ǖ���P�Lb+���ۣ���D�c���Y����tt��:��&��#;A���Ȅ4�64)>-��c��t�,g��4���Xt��@ E�)���2��gL��p�H2:�W?��FD�����{��� ��R��vm+9�"ǳrwdZ	�Y��"�{�
��2UYD�b��9���2{kA9�	���Ju޿�э@N��`t�-,�R���9�T�f�O�D�k`�C�O+��XWdI�$չ��`����ci�����]��
�ɍM"�ՠ�4����rf��VuȤ��a�5�ت�S�G3���=hh�tw����7�'���m�41z��i�S(*ǫ�$��٬.ݺ1��넫��U�,���	lh��:^��#��������R�O���c)s?�¤�N��?L�+ �j�һI���JӶ���~mͼ�J��8��U��"���m*�Y3��0�8-�M�C&��&����Ӱ�q����<��'���� UVcQ��/���'}�o����)zۼ�M-S�/�"��������Xф3��j�(h�c?2�|��sk<��MR������-�����\C�^+[U31<(52�}����H�����/!�x,f6��1^�sD]�|9�"	l�;��R5�����=�q���<lX��9$���yk�p�@5׼h�h��d����B��)�r|�j�Zh��Ѐ`�PTwc�y��L_�-���� g�j{������'K���h�����
��k|2�c�N�I2�1�)M�|)�#���J"2)Tc�𞲷��~n���а��?>%b�V��!����%������71�:L5���� ���6T��\��Oɒ;�����'�y͍��n�78T�PC�ٶ�������O<q�
��&ڏ��^���m/��`�*�0���	���8?|��4im-rs-Du#4�u/s{�LN�B�rsމ�A�Jd��JO4��c=|��n��<�,�_-f�Y�+4J ��)w[��!�Z�)VV�I���jo-_1䯪;�-stQy6a�� �n��U�z
�ԅx�w�r�qͧMWbX�W��mG�'�^��A�\G�m�6�E�%���x|������[�-��������2�Ч�q˳ R���<��<l��#�?GyM�7,�p�˗r�M���g&���/�m�hl6k뿖��=�������x{���q�d�����_�ɇ�� ,)z��v�j��v������Ё�z�=[�Ү�)	y�0��g6���%+�����c~Ց�V��eޢ��m�u��ɞ:){v�B(n����%`���[�k~�.��rA`�?�ڝ��<�F�-����ޞ�Q'f{or�tv�(�N!��]FG������ij�5�<,�K��6��K�w�����2K@�-)?ϐ�@�W�l�/�ۓ�S�=̌�4�}�4+m@��dV��v�4>8�>8BФ���J�ں��Q7��i2�q��ީ�`��m�9�_*)�>�}�~3|Hi���]��w?�5.���ð"<�yy�D	d&��}���x?'���S����QAC-O�/b�9�ݑ�A��gz?B͘`,�F��as)-/��5q:f� �tf[M���L���'Ra�?� R�ː=���Ў��fY���z[S7��L�Mm��Ib�
�=�6}���u��pg*��Z�$G'V�帜�V95�d�V��œ �H�-�r��]������F1'v_�9%EUs��':�`�O��0�y�x��E�:&Z�]ՙ����Y�
n|o�Da�2��0��=vJ��/���^w[%߿A��"YK��1ogL$��.�2^��4�*��ہ�.���S�K�
1���;�r�ؘ��	���iz �ݦ���f7�&�*c�`eq'X��?o�v�	i�E{�cy>f�+H�6A:c-�%.���s�͸�^��Dh�=�L��cg�Z
V�([_j����:�H����2 �Z�45�[��0Ѕ#�뫴�G����hr��jR�w��wY�{R�v�Ȏ3��.��H�6[�ٚ����{��8�]wsH+	MWM��D�Jč�.$�u�r֣P$�c����z�TLS/X�K��/����O����8�Cnܗ��p=�����r-�j�A�͡1���k�[(D<BS$�-�n�vb�U���UD� ������;>:Y|��	3bhŉ�&���t���w~�&��N=���� ��'*�#�ނ_E��d�{��_�E���i�����7Ӿ��9��-ǅU0L�LG���Xy�5�j:\��<bS�ux���]��T#������{�p���U��g%q��L[`.����̼85*�SGi.��Lw�u$)Q��(ob�Y����ѹ��P��Q}3��D�5�%�f F�z���;_w\���ߔ�1H�&ՙO&���t����u����U�\o�,������0vG�lvR.�梹�� �_�I�c匰�/T�߅A�,y��X��*'=�K�Տ�wO{���Zm�dB�e�ħ�b0�v��`�I�$���
[���n X1ǰq|h�#O����' 6}@F����O��ո��q�ީ��T �S���+�i����|���ABg������w�܆N��U�.h	���J�q��T�	�;t�;��Y�������-�~������kz��o[V Lwz{;f�����|�#7`��?�b{ j^�(�)���4펏� �u0L�;�WY�� C1�zk�r�[,�+u��%Մ����]ZًW��Tg٫��&����N^>}��h��������t�h���R�z�x�
�_$T�M�{��уE�8��Ț'��6(��9e���n�W������17�Q�㤹��xR�f)�l 9�Ԡ�l�������O�3�kB��d�esH��<�����(�`M8��U`�yr�&��bYx��qM�I;!!ܖ9�ۙ\�3�dx���S�+���H��5Ƀ�����m>�ueӨ�[�b�O�h6��[�2�`���f�������d9��g%��@�#�
|��F�vos��G�M�e3 �%Q����������c��j�'g��ṏ��J�mW������T*S��櫅��*�����yQA&`�����aj�\n�����$�2�������譨��_)�˳%�d�6��$�_���Q�B̙�=X�(U���y(���bv�bZ5�P0���f�T}���Eu�9$4@+c���\�^����:�%#�'�^ǗV����� }=�Ҫ-N���$�(Z�5b��Z�j2=�Że+��s�'�X��)U`�;�*_5 ��x[�� �&���EY�&�@��R2�a�7�HA1C�c���˃�S���hC��]>����B �#n_P^اz�����hu˿G������f>.:+}��a��!�~������5na�^x�T�]F��a��0ybN����d+�*�����Wl!�y\x����(�xN�5{�c� ��O��]9�'Y�֚UE���+\>�M�X\[g����FO�s��H���)����GX(TXЫ6�O��3͓)X���#���j�� 8$]$豚�Ź���6z*/K{��M�5�����No9J,b��$��c �+��9����E����خ9W�P�k�>���\�fP��˯C�R����+�[��E�Ô||)�6�q1�Գ^�ʕ�~IzE�E���D��s=��A�3��;K��>���5�W�	��Q�ϝ��9\6� �;�2���^�����R����|������= Ɂ}�s=P�q\åU�m��HgR1�/akc��� ���#Ajl~�d��e����!�
b���Ї
����+��C��Ѱ��e����D[�Xp��Rz�-,���M���e���Df�-AY� �)a�!]��[��Jc�K}𦵱`w�*�uS����0:���W��~;�G������,�xo/�;+�p�5�����FJa���"��D/��@Mg"O���8f�/`j�{�v�Nv�@�?�g���n�.������Au��>}�c���J��`+T��,!%�Gwy%@I�?�
�^(G�A?ؖ�v�y�(���ʇGy�����0wG7<�_����2@���͔������|��MR�_~�D��ɕ�:�\�}K[^���ce��8��=� ��8.�_�=�(v��a�L�I��J.��6���Y&���p�ґ�q�T\Fm�nh�3�'T3���83��K��2u�ܧ^xV�Ç�ğ�彙ȱ���$؄S��*$әO+��~09>�W�jL��ϸ�b?��Wݻ̮ DoO8��G��@~9��t��R��@��r��_\u|�@;- �R���D^�$����W
<R[`V��r����i���B��;��U.˴V�^���%m���t�}�,5L�K�.5�1^�� qCْ����$Utx����J*�]_�����;F�/~e���,�9�Niٵ��I`�zg�V���XdG-,K�&�_�����WD�P�o�A����i`C	�<�G�ut�i��#��l�ݓˏ�Q�u�T�H���/^�T-�h�^�SWl�V��Ĩ{m�jo�ۘ��
m������F�_`�?JEIq�{�)\Mg*2Ջ1�S�i*���~��s��J���ːH����>�Lr�nۛ>�b�zΐ���k�,��le�I+��/q<Q�9���%���k�m��Qo�$sUJ�eΚH���"(�ݿ(QX�����,/��%V�+n�����$b�T�Bs��d|��k��{�j���"�E��\��S�:��ׯ]2>�o>�JJ�f��� �Q�\�D�r�5�)�ZS�|�D�zzϮ��Ѓx�pP#7;2ܻ�A�ѻ��Cb�� ��Á���"�
_���R�lNE��Ȧs='��� (Dd&I��؈�b`����N\�bQ� ���r=�P3���S����ʷ&,�l�E]�lP�IU��W�J�T�0��#�n����s?f���:7�i<�ET������x�*I�"7v0ã;_o5r-�s-h)X�]̓$X�~[�䡵����YFe��4�����,��1N;� ?¯�{���+�)� G�ėV*��`�r:��^V��&F�s��^��t_{C���ZYh?<̩fK*5�d���kK��oAs�뗽�w1��K@�h�t�^�I櫏g֏�n>|\�r�����G�eL�;�Ø�뼺D�����?�Ϫz���{ɠ':;+ٰ����z�>4J4��4I���RMW��wrPJ6`�6�ka�'�5�%�o����3�#���/���ֻ��3�A�����:�.,���YTpBJ���~7�y�<�?5c����E�W�y��,�1�16k���:�q�>hO3PT��/��h)u�b��4Y�/jh-h��D�Mt���̀H����O��X�kɰ6����/d�:8x+W��YC��4�"�>R&2o1��:f��(C�n��3�����{xɯ,�R°W+T*��GgNo�o)ɐfT��#�THY_ڃ"Q�)�z����_��L��BhV�9C�Q*hxV�)�MPd�`X �t�6���L��F�G`IBC�@��L����V�(��%g"������?����$o��=+r�c�"L�] #4�X����"��z�h���ue6B���[�#�!����o�:6`�m�H���L��n�D>�	�lbgn�X;�a@�c	��؟w F�߾s-h��xF	��͈nB���C�9�|S�^�K�F��P"ܛ��PV��Ҥ.ɽN�ys�O��$;Ntq��s���e`��0��6�� !֡�[��U�M��K��M(��u���5pY�vשK3!)O�w����hM�lT�^ ^�`@�PCi��B�Psʀb�$\�ZV<�]�T�q���t2���lu��W��.z������m��&'��C��Ĕ����iDDϳ-9=�HR�<��Q�iA�#���[1�: �&��l.�^���jߥ��/x;pҮ�&�,����t��A"(�'�^�� v��"�|J��W�����Q?���`����TtrO�槾�:L���~\�1���Sg��O	�O�0��*�x����Q�0�%n)S���#�xd�(�F��t���a*:�wna�ߌr]�>��m'ύ93���XU����e��pȐ?"o�\|�lhe�OwhdW���J�<p�B�y����
��~����K�.����U�^��m �}�v6�xW��]�gC��8���Go�~0�zl�=�`���c�%��Mi뀞�QѶeȍ��lN*��F�u��T���1�&ѫ��p���8>��+e���XTN�}��`h!\!�ij�g�{@a~���� ��-p�96����OU03�����gS�,���Ʃ�՜�F�o��Z%��""^M���|���FI��g���z:[��3�`w�l�C:j���0U���Z;��q�h`q��hl.G�̢
��a�KiGyH��L�Vl�3h�1���|�bk	��+V��o���y�}d����oao�w��pD�Uf��H�z�ayAJ�3s������x�cQ<p��ĺ���)�}��:�	L,�p�i�`�n�ph��R�����r�=i&8vT������*z�W�x�����Oc���h�x͕��`�?P�`�2um��H�݅a;�?�6���D�Mw�`��7"ZH�s΋k�+*n�$��=��.�jj�/��	��n8���tN"�&B"7�z�,��Vla4{�q��	:Ϣ,�~�A0�"Hh�W�u�l�n<��S���\��3|R�i9��l�ĞQ��og6�ʦ�]��(¯u�Ntx���
�C�f�n�l*h��*�� �Q��} � �����o�e*�Y�z��a��a��I��5<��s��q,�t���e��޾��̖P���>��XpnC�"p���H&-�V��WS�g��.���F��!	0�ĕ�;kCJ�Nk��pJyir�k�����;�֌�[�/:�9)��+�[�^<�wS���Y� oLe�, �l�Rocؒ��MKJ�����A��1���p��U
^֥�2�?jվ��x��a<QB��!�U�Sv[ ����"�"'ަDhc�����]������0޺람3B��8�����l�i��g�QI��(�f�b ըD�7N��"!�c����Kb�~G첵��!��d�J{ʡ� 11
�>}��f�<?�v=���)`6�;	��:I�f�ׅq7� f�ێ�}��-X��B�GU*���'�[�۟���IW�K�4ͫ����?V�t��DC�5�ȟc��Q�8_R_���_�Z�J�6lᴮ�����ҝ���p[h<��Ժ��C2�� ������t%Û&}��̡�O���ߟ9��0:�h���|�0�(��2�Q������~����*> S�2s[�]�T���l��&��O긇�#�F���֩$� ��5�.�#�[��#��!���R`�y�/�l]�(T��-�̖ot=��o��Z{��c σ(+�e%�� a�`���E��,V�4���l̓Q��Ss;Zb9�q�)0Y�I�[�xM>F�����ᬆL8l8��y�b9y��弅�h߀.27p;:��+1Y���|��e���,v 8qlsTAü4�ܪ��b=$CD�Pm���+��!4���WºU�~z���t$���GLW�E�r�I	ӷ�#���A���!@#Qt-�:k̊�a�����n+�T�ˌ�Kb����Pw� 3��r]=��1���v�>���)6v�Ǜ��cR(��!#���/�mHW�<�D1n�F%
��>c�QO�>���~�vr��y=�!F�U�F�w�O�o�m��4�2�s�G$W�Vm��U�Ӂ�F�+�Ge�}l�vW�9\���MJ&�i�Q-����oaV~�6�r�������LR0PY��ke�ݠԘ+�qu��� 	DC �:u�B!����f4:\w�}�d�ւr���z�O���A(2+a]y-7F��M�Ӭ�bF	���L��B�L�q�e:Ó-H�"m��'x��V�#�ۗ��ƛD0��8���p�g#G㟄	͝�£�|P��O^+��<T'{��\a$�WGm�`i��p^'�w��y�yS��Z�����MrJ]�J�L�f�N�_�����l���)�Gm��z8�e��@�jI 򤋯8Z�ڴ��]�b�Պ����sE���\]�Ժ
��#)���n�Ù#X���_M�ƌ���ц'm�o����ד�yE�ɕ��7M"Dك ��;�i_Ӓ��}ز�����c@vA��)V,9Ha�f�l�$��<����|��zV�=���Il�}��?57?�S<�c�Á�[m�'��c�u�r��K�ԅܴ�~�ip�*����O�R�a"��K����H�ˍ��o`6�m�#���]u��l��چܧ�C(�rP����嚈�Z�E"o��:D�1�t7�����D"I��e(GO��kk��,IK�;K\�c2��
ٮu���٦Th]\����6��s�a��?1@N��Փ5'u�ה)�X��~�̒b@u�|(?R�֒�K�Ɋ.&�Vߵyk�j�]�Ĝ��7ȿ�P������H+�:�f�'�1Z�|���ހ���2����;�9��8�N�����B���)�\TP���3qX��|#;���#�dyx�Q��2�V�W/��BϏ�Źo�Nܔ�*�5��=��ʮ�!ߕi�Dŗĺ��I/��UT.�{�mM54��њ��ȩm��hA�xm��7�A���=��b��I0p��5�XS{Xo��Gz[���τ�K%O��ˑ Y��v�����3�*�R["�OH�P�+�b�FP���lUD��^�����ն�i"hl�r��ׇ�>�c8_���z�8�P�IÀ�����ߠ��w��mٳ�lq�h�^�E�D�n&R�)!a$�S�'�Fg�OJ��&5��G�l�����0��y�JZu)��Ѷ��EEH5rc2E*�>}����NL�S����;�?��	���[�*Hl6�9����d||D`-z���>��7y���iB7Z����XF�v����i�T��F�u�.g]T���uj�Ο��Fe;�PiT�C���/�ɨ8%�6X�F8Pos�@#��"� �M�x%�>J�_����ńe	���v@{5V���ZW��N����h�p,���C��P�q�~�0�ۡ7)��RlNIKg��e����4~'���A���[0m�r�����n�Yt��Eo�q]� ��yG�3�� /���A3L�w����;_����-��v�8�q�>s��r�y-?���(�m�
!`�lR��S�	l'�����we�& '�դ�Y���bF�ݺZ7?�"���7~�����H��.9�)�$�n?�j��P8P*$�gʯs��2N�i���hHֶ>�b�!�f�`�[)@��9�&����FF<�l����
�qEL��e^�)���c�P{1/c�]���H�f&��M�q�BU?;"��Mރi�3� �|＄��x�������.Ь#EB�%?��D}�mp
���B�3��R���h_�v���:���w���S"��O��.���!��tV�m�%��M*�dU����O���1t�~�\�*���_�9N`ς�k�į*�Bz���Ag
t����;Õ]���ƌ�ϡ/�/ڌ������j�9?_�����:�|c��L�g:��ӥ��,a`��ت��wfJfc�t˒�m�V����W�V��U�pc"��l���(g��QsϞsK�J镬�6�U G�=j�E�,2 ?�]���ٜt����H�K3�ƷI)�-)�pC�؜����f���!�i�8�Ϊ7'HbMĢ~ۋC�q ���J�:��6��BZ���`�%2��;��[,�/Z�F�h�"+C��qݷ���eWr�����סS�������1�X��Y(_�v)51nn�O��B�Q_��8>v�����k$��;�����4,o@ x����_}C�ոT��Y*��Jf�e�fd?`��"��/�!���B�)�  �g��jM�ZX^P�u���5�v����}��J�����V��A+K=�-Y��yp��_Zã���9prg_)��Nx�$}��j�c/���pz����K"Ųz,v�K��Q�߼��]ԣV!�`���J�+�A��A"~�7�("�cc��P�k�� fA)DM�a��/j5�O�>ο��5��l�!A 2;0#��ς�̔7���Y�Z���_a�+�O	��W��2�v��+�Ы��cruh�4���R���u)WV �� �@h[�����!>�S�d��[?%�&)]Vd�d4͑*WR;x��*��kHM/��[1QjK�O�࠾����T��kb��ކ�2��zQ�ذ:�_��P����꼑U�j�_��B��@Urg��z���6-������QK=��"LBȷ�BB_HLF!���$g-R�O)gJ`Z�,�����>b�*^V�F��V"k���~�K��h��X񃿽`:aJ '��7ЂX��ȥ��A�
-�)��bJ&|��b��}G�V�Q�)�D~~�'HJ҆+��R�3�4��-�p�Ү�IF`��c�TҢwK�mz#[۲,�:n]{�`C�'G���:N�S��lWq�����L�U#U���������� Zv��P"���c�ʄ!���Z*�H��_���$���K�0��kAr��,Y��%��S#����'A2�:5h�'�<�QX����ׁ��ʛʶ�ˈ��B����A�.����ᡅ�N�M��s�s���kwޣ�z&Lb&���n�P�7jR5s��V0��tK,��b�XZ���&�d�iY��\=i�o���yv��^�+/����)��	�?�_r�d�c�=t�ah&�L�AQ�+'�Í�Z;�%5�4�0��1S�������%V�r�$��qu5a (_��� JZ_�x��`�!_D�!�c�*�]eSi �w��h=�v����T�r�f�3z���cAS���"e��4��������0sW���\����5	��8�Ih,����I�p�U9�B�~�*}��q�W@�_�蟷q�qx��޻:�D+�������	0���5 �4��šJ��u���Y_��8�V�9Fͨ�B��Ǣ�?-�mo��_��3�h�G7@2�FIM��-d���({��>��ڏ�6�y��8�)�x��Hr� тiS�]lK1��+���y�6�2U��G�!��`<�&\/$;��֚�'��.}��4$DCYۿ_��K�[�?���}�ݬ��+fJ��s��?�Oz.������Bg�S�՟D�� �C���(�_V��[�$����7PY�Jw����j8oᏡ��U�ر�C��5���*[z�B&��9:����}�bi�B�N�+�b����2
p�������P�: �J��`g�2?�1�"��L@�Cɨ%���O`��W�#��Ј��8�=[�FdL�E!:	&�Z(E�����ʹR����۝����y=3i1o�����z�I�/�L���$�^��F%���ʅC� $(�����O�οT��a�ێ	)��jU/Q}����`�0���
O8��� @=z�:]�~��%	�Hr�1/�̙��&p9G�8x(�T��nf��	�E����Ȕ^���Kφ���u�%��e�?X�E|R���9SY�~�̪��r���ECB	^�J~o�WÍ�2�W5Y[&g�&�ds�.)�V�[�w�+m�n�n�im�����P�U8w~�Q|ZM�����y��PZn���XS����`��ޠ�Z��zo��f��sv�P�(��jLO��EN�@"�֏�"^ē� $�>��P5�.l\7a���d%>�I��J�j�y�*Np�yB��,���5�ă��_,�߉ �s�CrM�FK���%I�δ���{��XY���H^�P��K0�l;a�6H��RZ�₽�$QZ�$�D<V�������]�1��r�"��BG�<L���%�͉�M���)]k��e�v� ��)���*�A�ƿ���R'8�]��؅"Q�v:Ѽ�aKUqf�5�O�=��+T'װ�2a��J@q�������-4_�j�M�+kJ� y~oĭW!m㜆��?Q�*�{�^DJ�|څf1-�$�w}��A���9�n�#J�-�=4s:m����:O����Du��#6�1�Ӧj�/`��#�z�BLǽ9��b�P��u�M4��a e��X��Up�?�e1��L:�г���G��{t�o�V<4'�o�/�vcj5�b� 㟉W�*,��
U�2�8�� ����|+"ٍ��X�� 4�-�WZs["���*\TX%���&\8���U�+�nY�oC���]��o	�q����!2�U��s�b��N
�)r)K�ON���4���Vʮ�$�G�����j�=���4O�$��7�/��놴=v�n�>	���|ι2��#kv1��:9����m�����-�sS9�B�Z�����c�	R�.߆f1&NA;T���
��k���1����a���;�]	Az�3D},���d�W�Ts�j�{L�c���mb�;���[�n�%����
�P!��*�	��)��*�"k��o>)��r�/ӟ;{�c9M���� �#"�L�.(�͡0��?��G*2#� iz��}k��0ҹT�|�ҍ�@j�g�\Y�P�e̘.�\q�]��|s/�ojQC�PؐaU��~K�V>�ɉX������ 8v�8;v�o�� ��La���\п�Q���%˚^�_jN*�s��;~
����)U��1��.�@��!�S�~{����!��W��ؕ��SXV��T��jP�fuZ`�h	5RR��xmC39M���66/�
�f�2�'�v��b�csV/�R��6�0-�J����?NFjk Y%T�+��r�#z�<�&�3[��@b��X�l���R�K<���X��!(���Q{ ��=�o�u�m�J���k)/	i�5��Q�u�TZ�v��؍�8�UJ4�[�[@�A�Q��P����1m��u׋B�4=`9l�r��d��Ge�H�R��A�Ň���B��H��E�,��\��Tz�w�4O��6�r��Y�]�Ƒ��*��{���23|�Ĳm�aQ��O\p��y�^� ��]�h��Ed�e�M� ݗ��e&a �py0"����OD��7%��� ��cN��(&�����H����l� p���)]��(���i�g4bCP[�Z��_B�vM�p�@k��;�F&>@9 ����2i���0��с�w��#����""������Lؙ0�|��_���B֏/(��U���q��+�3R�>�Z�\���M�I�PK9R��b�&)#��E/�.',ڭ#9�ǈ&"ֿ��M�d?�9��a�;Jgh`)��3�����C^o*ֆ�}�mŷ��BJ�h��( ��V���Җ�4u@�ؑ��ΞMz� *O0A���c/��.�#졃�e�t��ʟ��������.��l�:y&�Q.��p.3��4��g�,���\��^�W{w��o�pO)`�hں��X=X�e1,����.uf��h��@��qH5�m̡5�lt��p��O��1��6VBm5h�_��%Wο�^8��eM6&}o&p�Ŏ#	��\�zZ�8�|�^d�����틙���-s�Q��j�Bz�1�^q$�@%!�@O��` �\]
	qWp��g���r�yyo�AX�Q�y�u�����G54W��a���L�<�`tYS�~	��X��)���@��B�;aݍ��~kݩ:ߒI�ٻ�뵥�ow��w�9X�Q�2��O���Y���qHrӢ�Y��;�X�|�3+���Į|C�؛}P���V�+��ȗc�cK�N�0��_$34˵XTj��z^�ź�`���^;@�!��igG���������X΀�.�!��ѓo���`/ѹ9E�BQ�?����y�#av3o3�x�U�Λ��T� �M�<]L��_�X�������w�S
�����_ܗ���aZ(��x�Pڄo��̵���o����������]G���C�e ��S�E# ��%�����c��`m#4�&�%�)��Vڤ�s���u�]���{��ui0}����g$��+�ɔa���F��#L�wq0�ĩ�􏾐�������C�|�F��U�Ǖ�!-X�vD�v�ÆEǛ(M��p��$ \��˸���=��&໤΋w�|A�9��b�^��	06O��զ��
��D3�Mh���0�@C�X�".v�m�g�"��3����gI8���vn�[T�v�G�4�I��H�`�p���ze��Bn��A[ռ�h"<&�}�
BC���L�[�z!�3�����%M�6	��S7�II�D=I���Ҥ�ǯ�I����#����t��YdqJ����iF�?�j �< -̀�J�hN����x��R��҈����{^[C�ὀt��rg���@���e�J��́q.��&vS17�m^8B���������%&���pH�L�4æ�������Hb��Ur��!ܯ��9]��Mv�}k>�}\� �ɭ'0��s#�˭v��c{&#p���Q���>c�dِ�j�y�4�{�����B�2ޤ*4��X���2�}�kcX���%��\.�GrT��SHI�^caY&J_��R�����'1n����5,Ot~˓	ݯ��B�jNĝ7��ִ����0��Z���ya�(���?Z�G}��"/�dq��Fv?f {ˠ����&blN�e��7�������0���J.͘O`G����9��Y�A����u,K��p}���a?���Y{�D�(?q������[u��ߢ��E[)RF�h�J����w�gtx� _�.�I���]����_tO�N̹�w�[�q���9�������x��TX�q{D;�5�\��a��M@�%GkƲ��i�'X�#�3l4n ��>�
�"h.h�r�^�C'�`��/��@�/H����]��QF�1,��6%@6��� �Ɣ%܀w��'�h���irR���sM�T/0DnԲx|z��	6��a��}T���'#?SR2�:?&�����s��Uܛ-����c���ݴM��;U�[�O-��@�f�Z:T~����+BDnf����N��"h"�$��
��pI�or����0�����@}H���0<�J���<��1�+�WY�~��q{�����}}0� lE����l������]V^�s2 {�v&܆ږ�+e�qy���X��t�ҵ"W���+���q��ڵ!��(6Res�2�A�J�1r��_x�Ls�x~0 ��r�9����c�A��h@�~��a�2�m�.:���L�ѭ[�F��mF	�A6kW$�NW��*�PE�T:��&�����Z��_�����|t<����FÞ)��v_��p�5{G_�5��q�QI�w5������C�N�k�@��
$�9�ˏ�����?auw�Nm|��+�3E
!k�΢Zj�Jj�ɺ��Q����|A��J0��c��q̻�·j�?
���g-���@88~�c�ݙ��*M��H���꓅-'G�a)�X5�9�:��Ob� Y�_� p���Nu8�W����L�M���U�����C�+�(�%-���RT^�Q2����bқ�ER�~��<�ä��+N��@������§c���A���qb����@�R�yó� 2�2�%���ʿߢU ��S���2�I��6� |����%j�G�q
��������p��U�h���{�iS:Wy�&I�#*��DO��x!��M-��$�B	�����{:ε���^�t�I�q{DZ�İ�Vuh��9���\A����	��83�ZF�էtP,����1��Jd�+8Ifl�g�p���((�x�qS�4o2��HQ�L	��U��^R��Vߨ�E6�m���Y�Vç�ḑ@:�<5t"s������㌀�����b�^>������ɋ{�j�l��5-ԭcs�DX+���5D�z���߅�-Sg%�iv���] ����w�$����>�e�^���@�6���y�"�Z�m��4Q�p,�Pz?8��o_W�hҵ�ƺ�S���
+m��^w�8"2~CPz��J��������{#��X����	v����9�p��,��JUX�_��Н�VH����kX-J+�b�SɺV�ß�V�̢w���t��H��j\ߙ�Mc
�ISw��O�{g�4oT�%���`�dL��NҐ��4�h+R���4jd785��Bs�Т��G�����6�Ei����VRx�|Rt��u�U4͆H��'��.����ީx��P�զ��bǨC a���vO�jL1����
�/���I�HY�n�&����	���摅,-�kL��$�,C��qd�@��~�{n�G������?��Qjp+�����ײդ���C~�g8�<��ْ��PZ�\
�9D�o,��2���Fv��jm�֦�v�1��I�|�0����:��o�� <D����7��F��
Z���K:�M"0+P��K��iף)r���T�����t簌��>�*���������	�-��Pp譺����"�=K���8N�9�[2Ku4���mc9�?O����¹��(���p
��c�����k�R�1^�Y�}�ڬ{V6 U�-�����Q�c#�ɂ]c�����g�H�]�%��]t�r����6(�W�:��~�n!q�ۉ)�l��9L@ʓ&l��s���^�pW.��	jM`���͟b�-��m��`/����P<%�u麪��>&� ���@��+2-vr�Y�׿�k��ڽc�8���A��!rk<�G*�+�d_�>e���� ��t(���}6IIdJ
=I�$�ߌY�/�Fw/�t���} ۝�,̚q!������������.�,R��V�/�xYv��� O%{aI1�
џ�ƙT�������\)��$�(�=*�ϸ�t�Q�_�x���(6]�a��
�Y�ӦC�nX_E���V���`)�+�t
�����w����s��B�<��*�i/�^�@�1>8'���j�W+Q%��1����d�,�2����b���0Qb� ��Ț��r�y��2�Z�H�g��&3Ix�ζ�1:�
~������SJwOm���e�4���e��k�&�9�
7yW6�O�A}�"��b�ʕ�f&9�1>R�ow�&/��E�Mj߂U��p:��Tn�F�=A+�1�=��>�bt�l����������|�^��.L����ŝ
�zG�n�n�����@sZ�K�G��_�
�W�ѹO���ǜCK�v��1����r5�ӿWo� ���`�!g\���)��f�a�ż?R�.����S��qtl����?���'@	��c�#���X=Q��:j<��o��˖�9zl��fG�}�!Dz�n�q��(���Ϙ���.2�a���u#���t��7^ՍL�Dezu Uү��(�\�P�L>��v�������������M�ɍdM�E�wόPu��Q�鞣Ӛ�0����&��:t�nj��M�ݼcA߅��nX�B�(�f�eel�3;�gj�S��8&��ư�@�}c�/}x�&kVt�gLL�gmӾ�a,ӭi�v���=L2�k�gthuEʢ���#�Oؽ�1���!��r�=+�D�>D�;�vKքJ�C����������l���2UH5$}���m������"��)ɦ�3�S���:�6���$9�Ye��zh���s��ׄ[>��He���SXg̗�L兴�w�rAE�`9��txyK����z8V�WI�c˓8�^N��X׈�Mg�`t�a?�2�"�5��>/��_�LC0*�p�n�5�+����m�e��2�]G�i��\mЇ�邾��������� �����������p>s׶�k���XE׭S ���r�G���-0��N"٠4��(���ӥ
#v=H�����-O�V� ��!��`��K�$uWk�� F�48�I?i��F�U�[��?��wR(D���Me�s���C�-��_F�
��u���.G 1��a�켈d����aDG�p��d�7~ YW�*xH��$��)'{[�ϲ�kX%<�w�L�nɅ��bc��0�ְ�n���i����F:�7�6���B��j��T̹�#��z��U�RD&�8D��r��T>ڳ/G��;�a_�C�*b�t�6���=����"�@͘��U��|�T��Ɠ�[�gw��{3�n*�
r~)�!̒�@W>��K/�xQLXe~���ǵ�cyocF�vH�*6	�2�hiEҚ�~���,�l��n	~yI)���j��u�b�����*،a.9#=�u���M�k�;:�&2�1��BNAs�)w�i�{����:>蕟��sצּ�����R��ߴi|܊�[�����&�% �i�����r(��c
���� 8�i�)�|�ȥ,�h'~������o�FTc�A@�7Q�ˡ+ٮY]5M���f�w���w��Y��Pb�)���u���y��P���;�U�@�U��D{^L�%�Uac�õ�r��S�̟e�	�P4!*�E�����	y�D�w�$챬�c7m�$[�� 6�����?��3���#������V�L���H�;@���Dg{��Q�$j�^�w�?PjR�L�Ȩw�P�b(WegD�S�߾�1�܃�'�+�qw��ا���|�����kӯ��Ɉ��o�L:1�-�4���W�$tϣ ��D�jI%|LHӭn/�K�L$�x[f�Zk��L�[�N�rb�{������+U@�)�Dn���i�06���3�EZY��2�AT��0�� r�.�&bJ���b~cinZ#7��#���ccUv��DzL}�˃%���I�ۭ!0'c��)ˢ�V��B�Kh��=A�o��N{��*�wV�^o��P�8���;/=�U��\�dJ�Ѱ��.���j�0p�2ҭLj���0���se�윈>����+e�g��}p%��i�]�ڹ/E����6�:'z����R�3�E��B{�*���\مF��Du���S�=]me��w��:J��ݍX�BrS,G�����/�_��s�F&x��,�l�#g���(�l��06��; � ��ո���f6~�/FI�W�i#�q� ��YoX�tz:��Xᓽ�陘���J��g�
�O �� ��[�,d4OM�<���,_eP�v{6��Ow12so^C$,'�coI۶�"����gM���&���P;��1ٕ�s�m�v�)c8���5�C�p ����,Z�<ϱ�ו������.��Ҳ=3$a�!i{�r����=	/9��r`Tջ������ai�, �#Ԏg pO07�l̞�R�#�o/��j�pէ��Թ��4O���-%<���B�E|��\��`پ��#eqd�����;6���[�[(k5U�MSU�%�&9��l"��tc��J��y�N6���۳��~o�z{jD���@{ �My�}��&�&�Ȯ>}�5HK�A����� ��o�����^J#$�f�����6����H��M^V#W�
&�z����3F+o=�"_1{� &��w{�{��|2�?�3�O���[8�+�_&y�?E���ҰrL��ޠ�8^e�Ǭ�s�4�W홣�u���#j=~����ڹ;t����c�k�F�.�3���ZAUv��RV����$
mٞg�Q���/�E�����.��ꔣ��[z��y~���U,��rl����f�Ks��P��O^4C��UP'�T��a3'x�~��2��s�G	y�|	�<��	 e
	a2*�by��MYa���e� ([����g���ϸ��ڰ;)o�~��k���pp�'w.�uE��gO�f��z�CXw#���ޕ��>"I�e�=�̖yV�5��m�-�Q;�kJH:4ـ�|"��H��Qqr.a��&<B+�����	|����=e�'��+�W�40��V[-���g��8����Y��(��~+Q���i_�R��,�)/W��e#ܧ�b��_�J?���F).φ)[�s2Ħ�q�B�a�4������J�w5:es ��I�G�a���߰�?�Q5�\�����%7L�³#Ory��ef9�s��	��ٲ0bz�Չ����>5T��J3:˩HZ��5x���3��u�ꨐ>@O-��f��s*�� �T!~�^8����ڱ��&9��LQ4��i�5��.�.�)��fŤ�a��l�A�emj�k�Y�j�?z��CU�3�pJ��E,�%y;����3��T�V����/���Iڷ(�'���� im�9l�R�x�od���� ����t{�G��n ���+����h��h��܌N���Ѽ� 8���>�m5���o�=����:7}� �p1d&󉁅[{�iZR=����
�{y��'��뻴���R�Jm�CqD�K+A��2�����'56���Y�W���/i��T�x�`J��,�����ź�
ĥV�]��˺��U�E�`ĳ�0'���:�$n�JVrdB0O�	�47����`h��q]8GF3F�Md���,$4ⳏ;]�g��3?� l�RU��r�.;t�俑�{��+�*�2��ٶ(�C�qO�e���1v���͓�ކ�X��3� �ɹqdok��n�PNcn��ӏ�<��qq�-e�ov��A�^�{C5ѳD��ǯ�TF�|������I�d�qj����_���>{q��o4�+J�	u������Υ"��?�73�����1>h�����uנpR7��yꈬ#�n��-e,5�O�P1 _��a�+s־�1�+�7�S�����j$n��r�����\�7<�%c��t�c�"�Ԍ�6u^Ǿ[�F������z�$��b���t��g^v׹@��$�&Q�1/|jFR�,H�\���J�������*;	tw�*g����z�<���R�'�Mz���X��%AÙ���׻fdD@C[��@���Ne4������N�n����$r��ٷ���Ľ�N�,�OZ�1a�Nd!	���S��[2�GOH���þS�Y��3��}9��XCi�@��T"QQK�}Q�@�8�e�au�릕{
��R2,��I�pCQQ�L^S���td��z�]�[�Z���c�H��zQMa=XP�@�.v-�'�3�"`.�|��S��%ʻ:�6H~��Ig�I��le�K�F�_���9�}
gT,���.ʔxazv[�\H�9���*ԴZ�Z�i�R@_3���2`C�T^��
��*���6���\�籼�>Nܑ��5�:��a4:#x�I�^���e����\i��wWqB�
�._M���<�Y[HՂ�����K(��U_m� ~s��	s�f\w�Y�=�)�j�^S��&�l�tp���͓�M~)�S�\_�U��x�d�_�Z>_��b�Qv�U�_��v>���}�Q�4�} ����2L��"/��)цi�@�tL���:옰�g 9�>�!ࡑsL.}8�a�o�t��֊��m�WoA�"�Ԍ��-�H��k}�&HJI��-�~�ZJ{�%�%����<<��35^�EV�,'�B �m[ $] ߵ*���S��ҧ��V�Ɏ�<:>�m>��tO�c��n����_,l��;��.ڑ�4 ���57pH�D�zb_.�bve}���^�g�q�˜��W_��8�r�,� ���q%��|��VB�{�z"MJ���C��3<�%��Ffu��
�UOPۿ����� �;��2�UkE�� �����ˮ�ԛ�w��ܞ^���-{�5�o T�zq�V�d�F�ֆN-:p���T���ߐ�~��
��ѷc�چX���Z�s��a� �$"]�=�X�|�k�[@6>�f28ꥡ��F���|�uĒa��j:gZ�󇈃2#:!������C
	�������^	I�L���B�����_� �lС�������1��(��_��n�73*f�S��Ú&!�	�\�E�O��cP�����G8�ϼҎ.!͌1��@�(�t�dj:m���j̢��o`n�2N��&N��i�!����{�΅��$uѭ 71�!mO�j��t�JQ,E!3W�ު�L$Ȭ����&G�@VCJ ��K�'�[h�:��V��P�Q\�Y��ֳ����.��Pً[�3b�C3ƃ}w��Yh��0ѕ�F$HC�������_#!�N���
��=��*��$p�����丝�0D�-������6
�JH�IO�i�R�ɇ��� � ��hӈ�B�|��DE-�̌F[��I�~.��6� _�8!>��?�kO�x���L�R��/
o�%w�f�X���B��$
{е�[C�\� �#�����B�{��� �P�d���\��-Hd ��c�V������1Y�\�:�@����H��Fv�m$1������	�"]��}�Ӂ��Q#��s���µ3��[��_ ��5���=c=$��쀜կ슝]/��&�ĕ���p�wK���y֥��ù�K��N��ϭ�f��3-�\�'��U��������a��Y���L���v����D��� �kl/�(�V��@�ϯ��kU�um�^�s��i��w,pk�nX�>�Y̇�h�$���O�:s���q�,�\9�)n�yf��Ki�c����b+ŝ>�>��YH"�#e���<h���v�E�G�~��X	qd�
����r9�|���n���s�甏���eJ��D��!0H%�b�w�^G�ʴ��q�U5(4��&d���m��".�2*G���?-�t�|]��@9���D��5�+2�8)~��Tx[^�p�`+wT��a�����i����	���p0�9^����� ��Jz<&(�����L������1���j�~���df��.A(A�hY�� `�1�E���$d>��t3i�.o�9����.�5����MEB����[d�(���31�Ng)3�:�O4TbZe6���е�C%tal�8�y����}���z���(��E$�Q����?���n�^(�
bA�y9��w��J7�ƾ��x	�2�T���Z�.��^�x�kG«,�9�n|3N�� 00���d�k����vfY�j��ޭ�qT���N��F�ڀ5�V��ڻK����Zw.�N:|I������)�--�U'��̀Z����ڱ�.K�s�,w5d��M�E�Q��l�JC��
�nvz�IOܣ˭�~����~Gչ�P��������sh{�u��|E���,J�����XcJ�Yn�3ze�������L�ƚ}l&�H"���Z¥"������'�.���>��w����T8�tO�k� 5.�R�>�G�:��=�Up��8r[�9u<�pp@m��,�����T�D.ڋr�����p��r�9���[��x���s��q��`����F��sOɰK7��'̨R�M�Rb�gn"eK��Zm��U��i��u�t:�ikPMT�Jh�.y�J�Z�ʆO
���i>�ə��@:�T�I%�{��oZH�9�R��*�U:?��g�����eUu����"6���^a0����<�N�ºC�d$�)����~܄(B���,v�
��������������_0\`k�)�NUA�UiA	͋�0G����J�R��
A��h�>�����]��VJ�Հ���Հ�
j涞~�+luyYS��S_�G�;ĥ�7��ߓ��$�.�b�;�Z��X�O(8�w�O7<�5�Ѣ�D�����c1#ڲN�GQ�������+F�z@?��w&]�ﭡ��6I2#�ή� O���C�Z\BbHp�u���4Z���� �?��c����@R�>h�gz�~��@",͈.�^H�pL7�8����7F��F1�gGbǙ(���-�(��x�l|ɩ�{O�%�
����슌+�ݣRA��Jn!�c�wS>Տ"-S5?���ԕ�0�>�3D{e���p ���g��8o��K�'pL��g1rdOh������m����c�}�O>z�M"�I@�' �e"6`Z�@�@���X�biE��~fn���BIz�x��"��U:0iؘ-[�z,�W�i�u3�Q :�i�A���}��2P�n/;��9+�������O��b�]�D�I��KB�"�4(��l�8��Hc�s�O^�j��,FِNχ�sN�&~��l�\}<:����M7H(�R��+W��:JƢ��|�?f�ɹk���.9����Q��(l* ����Č��r<:l����kO|V�l�?p��[�������V^7};؈��H�[�����`t�XO�y����(Ө����ݏ�|s7v-GM[�g�4Uȝ�E�1�����]ov���j(�!Ք�[�h�偕����Q���dj�
��M�d	Ar��x	���*�>y�\Rf�F$�V��P���e<I��"�.h��k��6!� h0T�� g�z�=��"��p�D�U�`�'Z_C�@fw�hk����4M�6B�Ś���|)�c��(6�����~qk7HP�+�
��kq}���>F�q���ڸ@XC,��������۪��~Fu0�j���5�n=b����CjV"#�>���Q{X;=4��U�!�mT
fT���.�ƣE<�U³��������L�Żg�~�v�]uBx%�|��͸F^ ��Sϫb��m�Z���R�GǺ	d\v�������*�mS�EBX��|E#��Yo'��t���ם���w�3�8�MY��-j�K�?Mb-L�Z�Ќ4U��y5�$]n�<4@6�y�+�9)��c��:'i?D�\��X�Tٲ�(J�<�R�?��|�Fe�n�	v���d��E&�R!�t���"����a��v�]&��"��V*�����X�?��ҙ�7��r�ϸ�|������mu���W�~�s������HѺf�{$~�!C����7�lx�7�[/:�X��9�=t���	%�`Eپf�&�57|u�J�݋X�!Y�&���F=:�����9n�T��-�J��ܙ�FY@X0c��
�y6'}�@`�u�rȲ��QUA��M���U;2f[+V��X���E��BAH- �=]�q���ĪZ3Wd�]�&ϲk�v�Rf V(�3m����(���^D�G��_|����fk!ܖ9p�&�E�y�V	=I�!�Kt��w�%0UZ�L�X �$'�� ���-®�7c���^��LR�Qd���رUg<�(]����lO�+��`W!<�*�/��஁K���@�7�H�k8#�4�.߽999 ,]��P��`�,A�������m��XyS�~�&� �YF�������dD��j
U��[��&�_vC,�"'EI�d�	<J�|���+&vJ.oUT�n��[��[�}'<$��~����$l��$�'@�{�^m��f8?�'i�M����{�ž�$q�������$�wԜ!sG_1�O �C]z��p�[	ޤp`ڿ����g7�+B����N�3g��������z�<�rO�--o�{�������*���������{��@9�Tb����lS�����?�,�;R+m��,6���r�F��Wx�M�n��b3�3��/����339)��[]1�n�"��J7,1�[�5І��\Zs��w��W��P~���}+d����f�3�^�mgK@ۄ�ø^ Que��+�B��20S�>�$qu[f�����<�_�s��Js�oW��%�