��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i��������J����L�.���w��)�Q�%������r���������ɗ���
�����|��S^҈�|�9��Aޝ"	?�qHa�6&��҉qь'|�!�/xqˁ����&���׆=yh�S�Ϛ-�d�ri VV�D{� Y�mw���NoO��GQ�� H���z�ѷ�'�s�&���vc��๒v���Rifҝl��[򥍠��z�\�|r}�zi	Rr+�W]��[e�T�ϣ�Tn�Al��
�}��:��tY�u��$���^���s+�v�|�t�A$����2�����k��Mb��!����p�Hj-��x�#2F��G��T�B���^ G���Fn�oN��K5�������J#�(���;la�C���	���F�d�z�a�-"��`��ea�H�Ŗ�d�a��E���C�_Q.�љ��7`⠦߅���<����c%.8��N�k?��G��4w*ؙ\�9�a �Ÿ2����C�P@j�|H�5���dBQ	`#�V*�/���Z���6W� r�bѤ6�h��LJ��P���6fv��n��XO4�c�4�rl�6�(�>KkC�
 w�s�_�^�.���X�7,\#,XUύ�D�' ���f��lrz���8g�/&��� (�<�0k�W��ig� �|����)���^�/�Śja���n���Ŝ[b��jD��q1U�x.o2R�(�s�k<�y�?56�L��z��h���É(���F�]�0���ҟ����h'�k��3���Ã�N-�����X=�a������িb����2՜=����@�W_f
��L㲬?�W.´�ǡ�LXt��f%��3^_���r��M�J8����z�.��Ⱥ<L����cY+�1u@Z���]%*9�o�'��;��Tc��n�L���b��t��h�a:�(��նGb0�F� �e6�:�NL�c웑6;�q�c4PB�ļ~8"��&&Ɏs�+��|p�ʋd2��+��<\���B3��R�U؃� ��Ӄ�:g}v��z�K��U`�ll�W�y=����kx�^~�Vr�_r��T��s�H��D���}��:����������|쨌$`���UԌ<*���P�A��uӨ6�_��E0��z��|�,��u��(	%��$U2��$�)��=�Eۡ?�.i�����Ɛۦ��Z�M<
�h�H֢>rv���\���~`~�n��3�)"�,�|:2g����+��p�������4���fh$Q�\lh2ry��)�@�Q�+
X�zߊ�-/]�:0�>�N��C�把�XK�c�c�Om�oo��w��t�%����ݝc�Q�����_���[����z�Ok���$x����uC��g��@������9��O��-�c�`8=�3��bzU��V�����y8c����0!�. ��D��'�^��>,����P�P��)Bx^�0�'�"2����m��$���8c�Q�|�bC�}�4(��JiGy�Z��5��/���.�u �'p�m���.+��¤�`ca�P\$ܻ���M�h�S�BK��m?P�ĥ��U.�x4q�P�⚁u�}~��|V&�#����󮦲Q-K���j�@)T�����m�)g���t�{x�ɢ�|4#�`��O���JCK{����Z����<��
���|b�`dNy�M��^a��b��߸7~���iY�cɶtI�Ƀ;tÒG/.�[^3LVcF��B����v'�vGw�[��Ct��@��y0��u�j(�v��,ԇG��0�8:��!U��>�CP�n/�d2؂����E"�1%���8q��������+�t�F@����>���\G4�QCg~�����dw��$�}E8��s�β�������;K�@ȿb��g���t�֣^M�r���,o;S�Q���Ë�|hJ��O��2%�M\=w��鼐9�KN�ͫ0(}%���1�y�Li��Ym���5�&k�~��ɯZhP����3�Z�`U�$>!_8��5؆E��y�WU�� ��;mJ�ڴ�,�-1%$4Gxa[�x#�Po���ͱƙ�cV��ɨ&�g�%��+���w��f�1V�3i�ßY��^N�o8(��A�srP��g~ē����2�Kc�ٸ�|��C�ŊwNg�з�}1�AY����ދ5A���g� 4M-�#��`'H�U���ƫ9X
Ͻ�Ï/��rĠ:�xL�b0Igg�%����O�_���u_��dA5I�&y�o�C����E�M�2�v5Nj%L�r��6�����y�uÉ�%�G^�sk�^���nj4�l�v��?C��	��v�*`6��A)����sn$6"�b(nП�d�.$̷�`|H2*F��J_�5�����bQ-�7c׭1��W�)��W�=�,(�.1��)�뎏:��c%��Oq럕�/ea]�" ?���lFAjT�GCp�r]C��]���Y|�(L��)��ǣ�ڷy��08y4`�c��v�@��C�����J	[���Э[��'���G*���ۣ��
�	�L�1�V�&�g $�\� չNA\u��9�����\i�Zf9��ҧr�Wx��V�y�+�.�,��b(���^�>��_�kS*����6��=8�u�!k���n@���L�;��q�c��U��=��qEXj�5d����I��#[��5�ڴ��
���|��?T��6 i���������勎���k������i�֠A�Ƶ~)XLc�(7���� Տg�Z�\nR�~m8���˷o `�{��w�uj������O�V;���p܌*#��zi�o�>-�b�v�2M����ʦQ�?�/2�ژh<8P�n��B�n���ET����L9<T�08� 6��v� �.�I"��G�@1���1���[D��\�9M�aI��(�h-Nܲ}\�����ቤ�e�Z,��#�n�4�eC'm7���uT�O::�ABI��h�E�ʴ&Ӄ�_"a�[�_8��هPG��s�Pce�%µmw�� �e%����zvu6����! JuJh�[gQMv�ݯ$��C�`����6�`�7�x9�Oo{_����d}����'������s�2P�Y�-�;e�j"r�r�W�wK�<uD������313M��5઱�sJ�!r@�E�g�����5�L�Ωv�#&� Q��>�)BSt�v�Z�tZ��]����!�p2��9�l��0�0ҿ�ޫ�缪Tvx7EC�o����y�^.�!�x���k�#�}
������E�o(�@���Ȇ�#�+8��I��J���^�n����~��<J�y<�c����P �/��O�ߪ"�,�)��Ɯ\�{ku&s���h���{X�Vb�u++��m���_�l�+��
��½�a��������Ka�~)�����9�H�lGY�h'�z+����Y ���w�m��y"�R�rS��%���Z�Dΰ���,��t�!����()*2����5Z__��j�9����=�ĳd�<��`QXY�q��b�t�-ˊ���RF�V#���ʻ��e]�y��l�v�@',,O�Zm*�G���Ar���>')�������>�~{uO�уi�*��B �fC}_C���,ER�U�d���& :ۧL�Ӥ-2�lۙ%��/�����3��#>�F=(|��4�G����x�D'M�=toRl��\���^�9��˞s��EP��|�_�k4��p���Y*yf��~9_��A�g��"�UT����hS�ep���Ka��A,�͈�M���Ǻ��gv�k����1a��k�B�9]qV��O�x��d1HA��F���ʘ�]���"�tJ!g�~�BĀ���ye���]�����+vne�-�"hb��� ����u^L7$�F��k�^��F�/�mx/��~BI�a�X-SU*:��+=0N�;&x�.	V��Oo����M(}E��MV܌h+�6ŵ6�T/v����� �=�9��c�M������
�ZD{*�}�v�H�cI��'@�"���:Ŕ)=��^D��s�������9����p9N�a
�/��蘝�V�T�@�믓�A����-��f�4;Z�7�)�D���u�b�R��}��YW�ݡlSo8p����@���\.���:}���8��f�Ɛ��De,fQԡ�JP��h��Qz6�G�;�*)��r#�dΊ
��jw�=�J����ܪW���*܌(ڛd8򖇁η�%�GN���R� xƠ�6��9J��a��Gd-a�W����=$���"���O�ƨ�o'sP!�E|ƾ���͑]lK���YT��L�B*�Dr1�c��c���F�\x�goH��-���h����0M7C���\p�Vc�|���aJ<-5���'Lh'���D@���M���^��\8�3ܩ�r��[(��C������E�#+Eh�(+D9r��=��������yV��&������������w&m��8kJ!M�T׿R-�M;yl��lA� &[�����U�k�|mV,٩AK�(���r��U7.�7,�D���)s�?ߵV�m�,����y(q���0t`���,���?/��K����H>l�Sp��+�7r��f���b��T��t@O>���ܾ|E�o	Ov������k�J�~EWK� �a�%f�N���oh�xm� t}#�)ۿr�߀��IL]�,��ݔ�8.Q�o_;�Sw��X�a�8|d�#� ތ�~�$�sx'���V��~�jp���
�ޜ7y�b���!N�%L{?n�7�\%�5O��GG����K�-c��#��& �;5������y����t�Z) ��1�).;+ �pN/Q�Ieh������� ����P`^�x�5>s�-E�-mh��(`��x�~<bՀ��'�meF�m���8�.;_n�0N�6-��\K����J�r�i��;��^gY(��]����,���x�~����iυ۳��l���8+�xZ]�O|H7� MX?M6�.��b��q���G����~�����n9_�I7Ci,��޶ ��*/��{@���)&�6P#�!��1�,-���ef:hHx\:+����`��5P�9~#{Y�����F�y�{S�S4Xօ	}�9��Z[}�-oU�n��h�v��j�U����CMu=˓����V�\����`�J�����������o���G��O�@�����Ω��e��w��`��Ujc	�Rúm\�QE��~�&�� ����i�	��7g� ��<��4��Q�y|'e`� ���Q(l+�Pe���Uk!�t��u���8���A,����gU�Q���73[��K��|�P�&0�l�Ͻ�׉�>.��@�����ޤ�c�G��j��Cyc�f�<��i��-���l��~q%
wR;�H��:A�)>á����̯�k�vÞ�}5m٨6m����L�{�=6��|�D��^q.2t%RT���[E������4�^����1ϻ�����ﹹI>�ׅ;\���j[یUQ�Y���l�v������K#�*��W���%�~`�Jk���4	x�f3����9���w$��`�N��ތh��o4��e�� �%Zd4Q�����n���l�hf��9<���j�#�M�RS�Y�Hj�?�N(YۏM��S[F�����31{G/b�
�#��u�'G�M�v���F��G�3/�BH�k�U�gRߖS$l���o���� x��-�Æ���o��}�f�|��l��-��Bz�؀�K\��E{���7���ԃK:�]�C�dH���0~����Ց���m���#$秵�"EO��iߌ�9Vo���س�׌bk��0j8Хra�߻$���
�z��MJ�jy�0�=E]��+�L�(�r�{�|��?wTA�_���A�5ir��e ��.��mn*s`#D1�9�j�#'�i��>�)����?��9,f�7e�R[�9��d�|T22)��U�&���L�P(��/gr��Q�i�ꢥc� ���؟��4b&~)'�{�W2���49؏1�i�#^��B˨ �U���-�Z.�1��������h'~��"G��6�+q7����9����R �%�ZY��J�p�P�W_�l���c�3u8�pHP��z��d�m�d�u���J�����M�y�L�'�E�m`֒L�U�wbr/j��X		�A\�ҏ�a����w�rhAq���K�;��X�/��_��n�)kb�!l�j�FH�Lh��5�C)�"�����+rf�����Ta��t��+zn��`f�京��,܋c�@p��ƀ佚�N0�A�n��N'5�����X�l�7�lSM��*Y%��I��W��Pjk)�:���1DA����5"��1y��8���L����)72�(���!`����\S�W�s����F1Y��	֌�I�ReBt�2�a�4����J{�	kR�EE��֘���Rp{�u���ٝ@oI2�{b�wn1��m%V�t�Ծ�Z���BD���"�1�1�ҿx@�2b�X���(#��_��gΗ��9eeۯ'rc���z��\�F0Dy��%&9ppY��)�Dw-ä���-�*�X$��7�@�q��/�.���v-#(���q�f��J���9s:�%�=O#���6�� �9�(�D��ߢ#{4~���E�<��d��i�e�@�z�>(����P�/��\�g-nY̦n�wK�S�E���XY�V�ǻ��G��#b;���nP����F,��#���,`{�51�C���q�Եs��b�m T���w�0>���
��oڈv�K(fU0�818�E7�u�+�~~�-^z��ęl�1Z9/L�x�n\F�3pa�J�tgF.�6�`.�ڃ�'���ϫ �u�@�n`��,��Rm�{cln�뱵���:W�����
&��}�5ȋ�9�������
Qk+�t�u�Z��S�Q"��ڵ	_�(.��n���/�ͳ)�ccQW"sP�w�!��h���a�22��tn��{G90$T�k�1��q
j��şܶ�4��H��n��g����O��_K3&�gD���bD*�ř�r8b ����-P��z�z�X9b�?�QaY"i��JS4y�_{%�f4��ehD����[A��d���j�ŕ�~w15��[�n(�!�`�J�\脘4�V�z�9=c��kTIXOIq�Omq�q�g��~N�
6�.�R�$��! u��zA�ɟ���V�*�ň_�����&hG�HJ�QUsu�������u 7;����7!X'���y����"\��;@�%k�[�M��U�p�SW���2�aĉ�kH!���A�m�/-��#���\�x�Ez(��u����u�I�!�Pt�=��7\ԬOⲾˮC�S�DE�� J
�Kw7�ݨ�y$3~�񴴸p1Z%����M�����8 j �d=z�`��Z�^�%���4����Jc��>��b8V������5��>�B�T�y���wI|����/��v��>b!�9�o5ui�2��x�r�"d����#�)(�ƓW�Q�{��s�w���Ͻ�9r�?/z �m�`Ug�	,���(V<m����Q3']~��ᘿ��p���Bȓu7���^����{�.�&�l2��n� �]7V��Ƀ]�OZ��E�X\p3��=����W�E��ų�/��sv�"�Pq�WZ���?�gۜ�_�?4i�.�%�c��q����a���S >V7ko�
p�-�	6U��	�� ��&�z���,�u�6�G�_�C��Ǌ�o�h
�@����������|uR�1�jg�x�es�?�����ah������뻻VTi�d�L4��0�����zA<��7��u� .D�b��5�5P�R/Bi?�e�G��^X�c���w��-XO���B��+jc�����5].���������Z��6\��	����1�HJ�	+L� (1�o�6E���N�����+M��K����XI�1���!"���U���wC �}�s��yA��Q��`���C�j�\:���tT-�r1�pLG~I���p$�L���cH%ـE��w���.��b�sI@��6���s �Zd��|=7���Z��d�������K�S][�T�Gǀ,x��]�ZM��z�ʟ)��-�	��%��:{�)���Q�M�/�h��g���Rٖ��2�\��^4��Ќ��%�Y9�����yA��ӦU��C��V7�zVH�V��~5���VB�#��ϝ[a�)���^�6�;$fn:0�I�S�0�ƴ�E%�̊��w��Zh 1�X�64Ջ)���+ut��h�lM� �_��F��.�J+yL�k\S��p� A9E�5�HΤ�rKnh"+�`Aڪp�$a�X��&
�8��A��y�/JL���<V���jt6���:�a�ԉxge�x��Lp���f�`�!�PU�.&�xa:|�
�!	_��|V�_k�(ѐ?f9`�B����4��J�T����R����wbi�.Sc�r#0�e���J/p!�h�Jԗ�D����΢ ��[O���2TJZ�3M�c��
0�q�Z1��2փ䷛��� �Y�Z8�ko��5��k{>�גSm@�:�"�,A���Xy0[T�K=���À~�#��^����9ʘ�>�:�������a�Zզ�HL���҇m�͋��[�ُ����l����ؑ�%��Fs��fxV��Y�>��)yA
��c公;N�|��R"ҋ��2|�n�[#�yt��:ƺ~�A�*`�~����6�c�G���qη�ߦ�8&"�K}
�\�$�u�1�-���$̛�-��dZU�@Q��t ��w#v/Eͦ�� �Djjs�3q��0�
�{���o���40ݯ�As��G�a�����H���BO����ޥ��f\~����s�o�K�K���9���<Q���C�5L�E~_�o�<����O.��C=�~Es���<.���f�V`]������ݽ2A��f��?	�V�}���I����
�O�z�F�rO���ioH�V�{����<V�8J��<Ǯ:�C\B�q���h�hn]9�)�4CG�펲�p&8>U !t����o�a�+�U�=�0(wt�*��`)qu�ЏÂ�s�<_屰�\>9�5�(L\�K�j��c1GA�&���U�3z�q�9�OII �<k�U�p�[.r<#�	��-���:{��g���B�/�ѹ�,~��f�n8���o}*�D��:WK�NBv<(`�n��]��c}x�ܖ�+���q@'��� &�i$a��~�2���]�ac�cdW���
���.�j6t8�u�9���-o���n}o�;]/{%q�e/�p67n�Y7�`)	�^ֿ!�^D�<*R����D�帗r-U ����At��ǃ]̀����gV��QV�54�4:e�c�yI�`pk�W�?�j�d	���Jn'��ʂ�R���1?>.�Ji\஋���i�W�'�K��,��q���d�N	�Հ�P�����-$iM�Bj���=�f��Z}�$�VG���dI�!��f�O�B��0�|?s�[?-i�Z�\��*K�C-¼_Fvj΅?��z;!��cĪ�qX�0�";��V���MDr�҇�hM�ݫ>�q7�=����9���R�DG��"0��`]/r���.A�:�A���+����۴B��`vM��G����#���b��6a���4�D%`��Y�\�h�.��{w/"%l�Ю��´�F�)m�Z]T�s�ȁ_�Ma��J<�L�"��	�*��<�w�L_����R��L���-8��k�A��P:�:A&R�6`�p��Tu��h图Sl&�\^����|���BZh~�ܪ�H������(&�o�A'�[����[M����У����.p���{�)x���
F��<hJ���c�jy�Y�i����u�3�sP�@�<-#)����O�S���O��GͬVO��0��*T��j~�'��kh�Y�C� ��������E�Կ�D����f�3��\���@#��(MxW����|������㑟���8����
-���9�>���e��4R�tf�͢��7�*j0/OO,�Y�����Kw�?{�MM�)��O
��hpd�姱�mұi���Fo�(�C����U a1���$�I�T������
����ջ��)�vS̱h�����,R.�5�}�m�\_Q�bp7�!3��Rq~�Ҿ�܂�@�6�<[w�b|<�`VN�Nvc��I��������:Kl��J))�B�WM��&�x�����4ga��ϫ=��|���-W[&�e�
+�]I|_�/0��ϒ��sa1�7��ٌ��Jjv��Bc6/*��D��f�,�����_�h���$?��!*��E�*�0���t?�>a_x���^"{hP��V?�5���M��;�4U�Mf��>Dꖦ�[��#�����7��o	1I��D��t��4'_F�}��q���8?�J�FyGhJ�! |>�sύ�*:�|6�����dR�Z�$���o�j �|��k�|LF�{=������~��9^���M\Mv/�	�e����:�^W� �TeR:���.D l�k���h4�<��T�s�2y���u��C2��Qn�f�?H�F~Ps.q|���c�9�X�+�zxp�#x� �����)���n���;H�!q�䚿,�8H�ܹ���g��(dr� 9V�A�� A�mԪ�d�>�{;�I=ۢ���Zk냜Ǥ5��Z�6.�Ճ`dbp�C�Ľ�5��):��lU�h�W���H�#אz`��\����)t����(%~oE��O94��WW�,7o�O'r�)� ˋ%2-�;F�5� �qSڐ�w0l�{^����t!;:�X�����O�?BTG�`�%}1�C����Ҙ�����^4�IC
����dǕn����o�#N�y,��d�~�Z�R�!\9�+m>�~�,z[�4�Naon��$�5 �x�<lo�D����h�~� By�=�	]��˒�A��-V^�̇�ſN�;٤�،�1)CEE�bu"vVEZ�B��@(� {��ٙ��1���O��LqSB)������5��p,���U��w��'-0/��[��r���`�~��q#�~���ѝ�=��Q�_��,_���݃�N�t����-Q�3WP8{٩������vU�Zի\�Qo�0�fd��>ƒ�Jڋb��m~1���<Ed�v�ձN�ss�����XzIP]4��4���ESrR����uw�lt�+X?s<`�p6��v��yXH*��-���>�[Ҽ�A�	�*�.VS1��0g���2���?���p��L��	hm�6�R�Bˠ{���������[-�V�B��t�H��M��� �q��B-��� �s<y~�{O�����To�QU�¤�2�M�7�O|��K`�',��t�>?R��7���&���xt����9H���c�S���������e���WHW��x����]6�³��Nb����,�}�v@v�s�Ưy��a����6M"B50�#��n-6H��*�?�>�h/!+��6F|�r7vS�(�����v��ţZ�O��ڴY�j`���>��t#�kC���'P4 ������=*]w�`��J����������P�a�Pϗ/�y��@d8��h}���3�����?$��$��g���@�'�w<g�v)8���y( �e�_XX��V�>3�.��u��B�B��i�1�¶E�b�kɿ�S�s�M7�lK�^�R��FMˑ�FQ�T�NɟB�:h��ǆR�6�b*O�5�>�y�XJ>n�NlJ���6�/���|/�ƙ�X�4L�W�?�������:�ZDĄb��f�T�g;�cU��'li������
1�n�3�:9�Н�L㏌�=�If<�"�x�W��� ���%�XTA����k�gi�Rq���02u�7"��Ӯ����!z��X)�8b��G���\�ǭu]&6@��u��G���`C��H��W�J ��%o���C3(ĉ7��E�M]r���Y��BJ���黮�� ���9�E���R���$|��Y��)U1�� �]�2�(C���ć_Rqd����N#be�W�D�t<��a�g	v;��C}�h�"�,�Ϫ�
���	=JOo�%?�m|p�߽�������}��C��>s\l��rO!Q��8��dj�Ǜ��;ל�B�%��٠7��j�a�R���b��x��)a��WCYx3z�[�ɷ���#ڶ�3��6�^�.C�B�!p+������؍	i�#R�~�Z�L1c�D?3��#����4�eY���K���㬚�pXN� ��6P�n���]tmz�jg�6���$��8ȇ7%<�)�
�8f���sb4t;��a��*O���Mg|֏b��j����KJ|��j�P|����`?�f��e4���dy<3$���2�_*�d6U#k�xk��7���~�9�M�Vm�_{�4|<R�՞�*o~�Gv/u)Yg�������X?���ɉ�J�:8��pY�W�[0���F-�Y��ǀ3�(�^5VmH���? 
�_��F��̎�9��0������j�g?��[�??��tt�
@%�'/o�+�DÁ#m�h��}����?���W�j�
�)�F���Ok����ǂK��w\dv�C��;�{�R��Z� %ʚ~��|����q5��]iX���\O���l���{�Z��uZU�p�LQã"��˜��YN��`�*F�Д��j�"�Ā/֠[�#?d�w��ء|kNzG��3�ץ���Y�f�`�C�8� 0տ�7��Z�+��o�y^z�kW_	S� �J�}��*�Ak��B�#�j]�K�2��o������1X=��$.�k�Tp�5���+�3�>�=��UX[��.��~�f���ꈭ\�~����s�&����L0a5o���'9>O�0��gmy�1S�Fb#�#�oˊX��8�DBH	��fut�#ڏ�j�q�q�1���侑9��TKP��*u!Z��9�|���`҈+`�;�S�����Q�=�Bǡ��Q��-��wF��d���wg*X7�j���R��^�0&�'�`��]N��&�g��\]���f�>�ȓ
�����:xA��ztJ��}8S����T:�v:T�����t|���n�<�� ���l���~����e���x���̀��M�X���j��|��>5[i�d��3��
�:;Ckf��/���!.�O#ha����=J��F9sᢆ����T4ǵ3��-kB?�bS�u`��C\����ނ��AuO����7K��'#��|����[��ٷ��q^l����d��J}��A�@�n�����2&�����R��BJ��X�ٗTa�I|���"0�|+�k'�<�����ß��߰i�.ke����׍���{N�DHc�G���_���m��Px�b����zI�J�i7S�4��/@�7�b޸r�<�yBN*ƿ�[��e��3���hc�/����w�|�[�� I:�߇�%�K��#=T��rmu!�{�!d���9��P<:�Ŗ�cc�!�p�z�}���N
�.�0�6WN��B��yTv�&ׁ]结����ʒ���@SX�G�'+:�������W�Aw���'aI���4�XId ?�Nn�A?�kK�6-�AR�-��'~PX��"��A�]��nd�:C��s�w���J�);�Eo�:Fk���~��QC�J��w,��%=�	J�.s\R��/�(%�L��0XV��-���!���)l�M9���$����b�B Ȅ�f�n]�^�U���ʹe!L�_�x;��U���4,Q�\rJ��y�Uj��Z��*2#G9�Uѝ��U�񨏖0�w'bGss�C����2h��X��z��M",��ϛ �� 4f�͡I�꼳��pi�7�Jf��*�� ,��%�r��Ez�-�q��[ 毨g��JU�rpĐx~�4�@⸢;�"r���R{��w�tW$�3��ͺF�U�@�מ٥��g���U�$��٢f?]��K�����Tq�ɳ���Օ�����U���cs⚀s��1���A����}]�>���2N�vmF�ޜS`c��8�]{��dU=���"�!������?���9K/�Z2E��f����� ���wy��D6�QFa�aF5���pYٺ�`ܸU\2W���BS�0駠J��mH�n�B����f(\6�<�����vg��B��Ҋ%w�{�3��:]m�k��Y� ��ÃQ�� ξ�" �8�JG��u�l�k���я�j7����򉋬I��T� ��$����E���>� �"���NO�a7�5`b�g;����.��:n��:�M*!�h� ������Լ<�����+���Z��j��(�K	Py|��V�,]S��o}�X�m)�7W�]���:�����a������g�ַ��@k�Q#[S��b�Qp��qڒH @��ɐ8����Gi�V�2:7ȗxK
�Nt���M���%�MZ�ѴZ�';���7�����[�<+�%	4�U�r��PXC�����֔i>��"Qۓ[��n��;J�f�^����I�w���26�ip�`li�\�X��s���2]�W�lj�J�"��;�ڶ�(�]�I���c���V�k���?ѯ�Ĕ~2�G�C#g�h&�M?�(�a��ep��ď(7��[H̕�g4d����Ԣ<�=y9%z�"]�O�1,G�S�>K��)K@dy�~Ps}����x\�8 t�[�	��lq�'��o0�U�o�Z��	7�Rk�&��`�T��cC�x���B�R��Wk���G�:�
�sA��9�d��Y�}�Z�� x��U8k���|��.yKu2�ˠ�Y%����S�	�n����,�6bF�AFZ�����#a���9i��cȂ��24��
����u,.4��o�	@��8p/V��%O�Z�2V^���6���Nչ#_�U�),��^7F>�b<|Y}�n=ڢVDAT� �V����������M�=��F�ߩrCd���y���f�o�|
���5Ϡ��؆�3��-8̎�'���\�:��%��`pX7�W�Q���Ȟ���.>��V�1�{疜�CuvM�1������O	��A׌q䤅��CܢzH+lB[���d���Y���xtQ��5/pe���[���e�
�����#���)��8�Ǥ�ED��tu�3$u��)fuG�Z���^��"5(0_���q�T6��V�ԥ�d�@R�p�=���\:H��yrXҡ)��"N-*�|%����f�`]6Y���e��؀R�� �W����\(!�?�k���Y$�>)�Z���Ŏ6�yCa����D�v�.'��v��L+��[/ki@7���3�Z/eH���n :`���6	�M�� ���<�S�go����6�y�Z���+^9��`���Q�a������w.�������q�(��v�Ux��R�5v��6%��3��BɻX�������͚=P>sS�KNC���B���G���܋���)�%�XX�����B ��ʊ!���<��J8PN-{���G}Qv��0�2Z�����4W��<�v6���?����3�?UuKSRA���Y�?g�XfJ2?1J��t���#c��6<�[�|�?�p�oZ�#ΕLPaX���*�s=�O�`�5��^F��nR�(�}$�v]"�o���r�,W�!H��c=�5�NY��F=�ۏL0�@&��c�t��!v��;���:�ƾ%3��L��58��9J,X�"�ʦ���*k���0��m
��m���fy
!��BF�mE��#⤷X�KcxHg���b�
�� ��y��8����Kw�C���Ǫ)�����hb'���M��c����9
 ��S�2��W��q��\M-7\��6:Xȫ*��l����.e��}_ۻ�ߋ�����o��u/H{��r�z/��T��!���r4���<H}��ӊ�:67h�*����c7��e�<�+}�^o2��Ƕ2a�W���"��'cah�\գ:F%_��-�۬^U����2�RvkJ�${�c歷�p�.ߟ��(�&���[(�x!�w̥���X��W��X�6���Zd(d�_�a�B��T. �em�̆�C�vß���(a+G�h�@�Ǻ}�{�	d��������qc:�&�5��r�U�@�ntX�t�s8�
�>�Sk�<#�U�2��)W�9\G^�~)Uq��n_P:���w
�\�`�l��P��('|n�]�� j2�R��X�R,ނr�Gu��Zr=�e	���W�p0��Wr��z�y���,YZ��H=�����;�y20
�=`�Z���&��1,��(P��:�Yi��.��FѸ'^� �:{��6��fAB�V��0�}������E���"՚Τ�n���$Yz��ӓ�X�/N��jW���G/��dr4ڋ�k��&տ�H�u�Pr㮗�'�P�Zh�a���ɜ�r[���B�L9� ��խ�Ch{',W�䈕�����ׯ���G r	�;W�{Qt)B�
�V=_��i,��$X-r��L�#�/ɮyr[�!��?ƺ_"nJ$�����R��a�Q�\�77<(x7ڭT�xuUv(ۖ!5y=�	�`pg�Y��?_����`bD�I����V����A1���3ėo���N�1r�L��nU��6xI�ָ�k�(��߰��9Q���vݱ�ݕ�\���wWB�� At�S�UW�T��ք�;�-���/X��*�`������e�f�9��Kq�b��6�g��,igMAI�U/�?.�u����;�ZϹ2,�}��}����Ά�ך��L	���`:�`�&�=�	cS��o[B���3ڢV<D�4��ål$8�n�}������o�6���'Y7��U�G��(��|��j8�X<�\�s˧
 �9��X��G�C\_�|oLĈ`��'YH��c.p-�q��D�G'��b�e�� h<��;՗��`�֟��.b)$�������kk)�_�F�Z�J�̐YB��Zy.���r#�9Y���?�'�|8�=I����lJ!ǽH����/���7�2���y�Ȫ��C���x�p/u��g:����0Y����c'�bg��
��[3����[��<Z�����P:>����\�g�� 4 �8u�F�ҩQ4\�?����M�,�KyN�hm/+r�I\H�&$Td�\��8�<O!9p�f1{�!��|�Hee�������E|�BN+�p
�n�)4�/ �5�+U&����+��h!����j@�w5�d��/���٧R��H��Q^y·>�`Z���:`�����iV�xi~3��Z��;�p4��rX���"U�q�8�pV��Ϟ��� 0��F�V�#�p)��Q�I��xw�;�j�t�5��B�Ғ��ի�$��pt���/#̌�VF���ڸB�L�,+�����t����(�������M�ZU�5O�2�sw���GUS�(}r�����X�0xhI�~�Z��>�"l��b��. ���"�\��h���?d9Oq��0�]�i���j4����1�u��H�r �s|!v_�O,��#B4c��������d�K��P�������u6��%q��b��9u�cA��V��<rz��bgb3ǆ\CTXL���Z��6V�n2p�e�qZ�.�c�@�l�}r�jˣU�:J_�q�Fz�/�І6؜�:F��.Nl0�|*]�8���w�ph��(%ԕ���f�#����� ;[�r+M�%h�*-�["˞�ß=E
�E0�>�X�"(�$0^z�=}��$�v�
U<r�����)JQ!('���|VdN�ݍ:���,��y�z��Nb5W�k"�Iϝ�[R��tn"e����u�X����G��	k`CV&�Όi�Z��ޣ_;�ȱ�v9mڥ@� ����/�b�M���p?�	���|w�wL��-�ங�C�A� R�ι�F.�"�-��μ�����ea%��)C"F�"^w�ءc��S��Q�Ŕ�.F�2N�9�̇Wmh�vd0m�*%� �O�K�	��1"ӷ���I���� ����T���r	4_����|�%|=X=�+��(V��1b�^��m�h���S�����]Y�3��2��TD�P�~���g�6:�m��	.m�= Ġ[^Vq~�e���w�
SILa�|�ᔌ�-7kԡV���:�����S���#s]X���+������Y�Č�[��4ּ���:m]:+>h�L���)fVo>�����+�w���. +c�5�?"�Cl��k։��5V��]�l��Sů��<TPى��Uz���|3A��(a����Ӑ[�jb��+D�]���q�GZ=eTm#0��I+�S�%�����bM���Ci�׷=�� ��K�{�A��Ï���o�U��]�����`��uV��&����k.eO������ܴ��+Wq�3�Π๥s[z��3F�=�y�S���aΪD[b���`�tkXz�Zo6�Pg8��mF(���Ks�ذG]�E��i�3у������5&'���t�y�)�^^��?��/����1�y��9)�9��1����D�����I�Q{�H�3��_��t�W;Ps�D�-�������	����u��g7���?)���n�Օ�kÇv۵�x�̭�����{���k��=�{�?��RG�
I��,����qK2�3�Y2 �'�@L��S�6V�E
�ȼ�s]����i���B̨��)l��Eڌ~�Ǧ�U�/�`1{�u��T7���D�g��8z�3�Px=���*���nX�H���! l�ƥ�Ņ�6u\�{�� x����U�(mw=����q�����fk컒�<j%N2�S)�K��`7=��^��٬��I�@IX!����;	M��.V���:�����\`(:�S3�ܲ�\�+^����9�L������֐�/�w�L����ct��� �����������Tν�=+a�;��8�b:���:��5�l��"ā@Q} d-��� -Hk���V�hza�b�g�S�=??���%]d*���/�ܭ<�����u'5��2-U�c�w�NP���V�鱱K2��/�'��LϜi����2�B(�p�������P� ]�vI��p�����ynn�E��Z�����g'Z����j����ͦ�h���\�o*����@���\:���d2Θ���h�@��O���T�R��Q��]L�eɈgϿT�% \�mdV9!��	{�__gk��q�J��	�E"I��9z<е����ؐ~For`Ve���ս9�B�2�mC�Fb�d��
��b%�h��H=$�����#P����3�]���󯰓
�����a8��4 ����~�uEآk�Eϡ̍���L��&��\닔S����q��H{N)EI���&�f��s$4�'Ҁ���k� ����_���&�����飠P�m,9��C�k����Ľf5O׌CŦk��Z~on&]X��I0)�PIk����$�eԅ�m�����7�W��1Z���{3��}����aWQ��\���C4�M������c;�c��ޮN$.?�&�AI������c�f�	(�_�RciQ�XN��\u���S�h�f�v�,%h�V��lBk���u�0b���.�J�1	�}���^Z
-��\]��I	�R�]�FN�_��D1
�s����]�y_p��*�+,�܄Edmi��^�/�d����1�1�h9 �S��~	�[]����H�������D;u�I���l�!r2vb`7&�&}�N�������<`_C�Pr��)>��0�ט�;06
��\^� ���7�="bJ�f�֑���<�������f��I1s�$�>}0�V���kw?"�s�SFYUO2�?����i��U�+G������8H��/�g���v<�Lh}� ��BV����|M����?�<Z���{n��P���=h�\� Q9!?�@8�çwv�KN�2��%��^���	��3!u,���ڵ?��[��E�.����� �nmS�� �%�CY��>�ۮ��v-����Jg�(sm_��;({d��:[`�3�a���xA��y�t����J"�	t�>:�8��k"!7���2��×$�T$O[�N�w��!�߉l�m��J'a.�N��p6U��6���
��,������}+q�Ŝ5���?] ��4ǋ��UF��+�e�Z�Z�޿A'sG����� Sf�	Yq��v����B: �Z�T9���1�	`�7:jG(�'�:�#Ap��F@��,,���K�1���xq��P�8ʋ/���3��78�E��'����`B�7m���n\�ց�	�m���"Ԃ��|a�繞����?n(�a��@>Nw��L��S����m��E�i�����ə']��:�G���X��i�dL+��^S$7�q��"��o_��&_]�w~�Fr�*��Y"��^��sϛ\ʡ'߯U6���÷�z5�Cg��}� O�ю�e^��b���\;@[�-���0�`��k_V�&Q�l�Cܛ,�C�8�5�������M���ʲ�����x��֢@��ӥ��e�	Kj�oݨ�����/r��8���j}r�CPq*c,�5��V�����˖xv��]\����['�gb�]�ŗ!���㸢LoU��D DW^j��q� ���/����Mv�9�[����6�4z�¡����2X��K�Ōz^��LF�|X����A|�}���f��>�}�X�{9���g&���%$��JG�h�����J�^6�*�B=����> ��9B�wȤ�b��	x9L�Ε㘫Yo��]Q���Zk�+`-�g��ّ����{�ۼn�Qi�3,���CZF���by,{e�(���X���hB��#��P��k�U����)W����$Ǿ�t���X��ꝗ��.o�7T�ǚ;���+����fX�QK��S��D~l�BVo��c5?yJ�{�?��s^o��k=�'N;�;��U������x��yQ~Y�}*��4R#7�Z�Ȥ9&���;CF(
�xX�
V�E�)!���y�dg�OBԯ+��epsP_�[�݉�����e]^{��D���ĭ�䪋5`�țOl��E�Z힛�K�v����q�7��>����Z���¯ ʇ|F�O��ZW�`�L��=�`J<ql97:��MG�>4��=�fG9w|�3~+B��%�VhI�`�]��L�E���\5���(�$�� ���_`��B����9`�:��98�P��1w�Z�#䠍LY�bL��$��Mسr�f|M����������C�|2�D5�c��k�@;���FT�;����iJV�?��2ڰT�03�O������qi����.����Ǿ3C	�8����Q�aL�l�glp$W1��S�+I>�L(�j}N>U{,0�˔��E&��Dm��"�[�����p��+3H������?[�X�CDd�ˍ#[֑��z�����&����^y�wي >�Q��
X������t�j~���>>ko��R��`:���o7�����.3ߜ���XȪB&�Dm~4�i�V�@xSR�q�/Gx��}���Y�UD�:N�c���C!-f ��YZ��T�������A}�B�Ȗ?dX�ì�#~��^.��n���I��sL	��g���H�D�U��;Wt�--��ҏq�S*����_zS�]��[�S\����¯)i~%LR+iS.�����dwX:P���{���4��UM�v����_7wgb�QU�0�'�s?���I�Fy�����Vߴ���_�B��:��<�ǜ���=n3�0կxy�d3n� g\K���ZQ͕$*�1�%�J�+���[I7�!�!�S��O�ŽU2땾v_�Ȣ��ޢ�ƿ1[:!�����|�D��u�F�5Q*q��=x���\i,#�C:p*�A�1��8S�^��o&C�a��i�>������ŗYVU{d](V�k2k��$���\2K2���h�������1���b���qBVw�8��G�9��V��_�>�Cņ���:�+j�Fܰ�g��!5���CM�����{�5g��j\/�޾@N�#�l~S�|@e����!��=��ƫ]����܌T�.4	:�h.�����0�l
v���|��=lp�@C��nkjg�N�]��d��O�)���<(�_����Q��h�x��H`K���Z�J��1�����!��~��x��:���g7�Nx�Y�{��"_��&��� g��%'{��,����ݞF�[D5���G�����2��X*)�^�U�K ���l��?�D����Pƒ~��	/���#��㸉�_���G�`#���nT6�c�;`���������+�=0�^�:�FV���&m��8��U�v��H����]��rsٶ���5t�q��F�B�����9��"��,�.�R6��B�(���)s.�/���='Lw8M�:�c��|E��y�%RAƺ��,�۟��b�Z�%�Wy��$��Q�I_g_W�M���>�_�ĸv`}�Gs}q¡۳�۪0BV�q���YN����U�2�	��[����2Lg4'��pkZg����p�U�4��ʭu�DUK�x�-c��Ԕ�.5�4���S6��|�����](��7B���_��w�t8����h�h���\e�4��=)��u��i6)O�@�_�d���gBT��=��]��E.��D�ˣѤxa�f���r��Wn����.Cك���j����VD�ϯ� ��@�YݵV�G��F�~t��ڊ\dn�a�v��y/i�l�JY��/����=A��jJ�d:X��θs��-ؕ�	�\h��P�곀����8�cN����� 5�� |j��U9O�>���%"��Чo�mQ��oP5�tsr�ru�B���0�D.J��`�-�nn�v։��n�v������Y�����n�D/³�nGj���8Dc"�!���<��ye��Y/�����{��������M㕂p)+Ώ�c��t�
�d"<8)�����G����b[S%X~�{1M���yl�C+%�'���' YS�'��Y(XYZ�s��[�E�f�.Q-�
/^�V(c��g�9��>?v�I%�u�[�Ū�6>� �-��׽�{9��|��V�����ի����<5�$4z���1/��'-*����E�70>l4HN̋��UE����4�U'?s��-1_*,K��>��L�"_r�����i�礜�d0T&w�4y�B�>Ŧ���La`K�1h�p��uh#3�"�Fzo�">�z�يO���uX${�q*�T��&2*��������8@��G�1�����Ȭ���THv��K;���TsNR��o�`����kKJ� {E)����b�^|���*�@�Rv�sgZ<>�Mz�K6��{��U�����0��zf����ze�A�o���^Qv��I2Q�C`����1�fP�"�K����>���t�7���ч�����8r�ҁ]�~`K���E^�HFmr<���A	xhOJ�	����d�C㝸w�:0�c�ޫ4���V]*װ�OB��F�^T�l����`:%���m}�Ĳ�<�xQ��ǎv/���5��rFX�3����������s���/�n��55��Z��[�Q����'����)���r������p����p����?7��5\X6J�JR��L���<���$"~��f�I}��)\ kD� ��d`r��K]�=c��F���Upl��#�"o��'W67�M��H���|������ÎF��{��Ix�sKl� c�~֔��'�.<�/�8����-T� ne���׸��X
 ѡe��d�����7P�ư�rp
��������yX�[)���r���y�
4W%�����Ql(��ـ_��Ұ�٩w�֧��z��� �_��8*۫S�C��ٟ)�F�'n�PxA�
���$��ߦ�]0pփR�\�څ�og ʪ���4�۸z�8ވ0��Js��f��	r���ΤW���y�;o�T��J���8b�T���� i����Ild^ ��+�dF���~E��JB�IH��\�8����w����~�q�������̈Xi$�O������C>�U ��s!l�d�uXW3�Z�|<��7d�&ӷ��O6��>%F��+U����O��q s�FQ@��(������ҚF4Gk
"�\ch(E���7�'���g����{6|��
��|?ٰ�>�������i߷AYd#��0���
�ͫ����B�AbMl>,��㋆tz������j�γB�o+a(�w<��꯬��)�а3v�&�!�w�1��$@}J�Mp�U�M�2�?��Ƚ|0�e�1�I���7���0����d�������J����7�h{���3J��n6��2!~�i�K�2����4\@�p�nIQ�+�����}Y6�.����R����'��gv����9��%MB�8]e1�ؔU����X�-@��G�s5��Xظ���=��.�Y��!���Z���̣�����������D�B�S�����oK�3�F�|iFE�E�m���.muc�!�g��ۂ�p���:����q{9Z�Q���aF16ZŖ&�f麙Ob���FA����7��4Ԩ�?6E�՛��8�N^U�YyTL���"+����0GY�m�\C	��P���3?� V��Քj���-[�AR<�Z.0���']�r�\�vIӣ���+������:���I�������~��VV
�Niw���J5y�wf�|Yzf72�D��bdS������>�?~�3	�:�qP���d�A����} (E���Q��n�X�qP�6�� ���9〛Dp_����JK{�K[�����2�͍ޝjˍJ��*4{~��6��]�K��s�	C-��ZeJ���l0��~�E�~%��;�����*��prg2���'5s��XHzEe��`����f$�z�~�_�m4l��~25bOF��V8�la�?�]k�j����Q�ٟ�QV4v�]cV �T��*��zW� 2(47-�ح87�����y���֎����ە�p��WuV4�N�M�CAd�J�q�L1f#G�m�k�4v�����O�9�@,���d��o�M�h��$[q��An�(gڛ@��q����<��߉�/⸅���}V��r1sz
��n�R�)����i�B�y-B�+?.@n�>��Q��r���]�������L����Y��c�b�$�{�+{1UÇ���G����[Z<ht�f���O#�\�	T�Rd��߻>���5��ZM����+�ns��V�i|�.�C�$@��J,WW3@�:4�D�Oͪ����,W��98s���[Z�V��W�W	=�e��J?9`A��B����N}䃘��kp��&����[��|G��^o�����I����ʅ�������!}�V��fy8�F9YЭ�D�aGSM0���ܻP�V8���p-��'?E����?β��>���%5������}���B�7P�H����4��K�,l��Ɔ��S7$����[�L��k�a�%� ��N]?���b����\��>D��ȑ��n���2HV4՘��Ԍi3[��N���x�����mZcZ}��\Aӓ�H|f�*�Ͳ��b+�ٝ���¨��1��h�6#�-I�]�ٔv�C�7B�C��"Ge�p�ڝU����ȼ�O���v��5Ƽ��L����їB�ʖ~�>[���AbW��E��M<��L2%���S�(qqjE��&�(���u~�d_Gi��C �Z���gY��$�)%�:��2�����o��pZ_'S�_3s��a��5�v�  �Eަ��g6��,����@dV��A%�x�sR�*��=Z�m)���۪�-!۰j�F�-�РI��6�Hd�Lަ�{��4�U�o�gf5=�EҲn��2ɽPbF]��|��pv-<�!�%uDo!N�aǉ�2�T�> g#H���<��-�/� �X|��>Xc7�����7S�����P��.,Xb����b?�\�^J�_��8K��$p�mwa*�M
�Ў{��<8<e�0w�U�Q��M����n5zږ<���(|��v����,�08)�ㅎ<�*~��ų���҂S=�%�D����:�g�QT�-�^ү���i��z�),(���I{�x�G��P��7\K#
��z�<��a�ua0�K��k[M0U�C�L��u5fK�`�O�UE\8����$k��eT�}���� T��-٥^�:�TH
��F��v��� �V��ط='�����#iڂg�=M�be_�m���[V�]k{�l�[|_'J�߫�����Z� ��]���~�tr�wؿ���ldg�(L��XPP3�U]�(b����XZ��m����2��.օ�h��<�ã��(f��'vtq��ה�L����`�sqEa����0���|H��������sh�Ņ�g2�J�*
 ���34��>�Gc��pb�0)j;U�S���f�}%A
�"(b�U|,=�W�@�˜	����=�U���kn�5�C�n~�4?c��.�%l�!�;�ɾ�}�`�s�?C�S�!H)o�LȽk�8Z���n�b6�D���6����Ш��{H��^�3�_*���Q�΁�.�*� �8g$�[@�^�E������{�ן8�uT���_r%\���>�=����^��d�����O��*���%d�a��P��Uq���Z,�����;>���^��qqK,q����8	o	�����
�},������)��Lm�"$M�����I[�L��~^�F�?�K��oFH]����r�O���.���O��I�*����.7p0�"c����3*�W�c�樢�^�.er������bj�r~�K_�s&}��G�Q�)�@����[nu4?Ӫ�h(F�]�W!�h��F
$�T$�kvwm�1�Ee��������#/Gt.��4T4i��EE	��n`����7P��@�ݔ��f��(���ܜ��0�/f�
7�JYuB��w\Q��벾�Yh�VƧ�G�H ��[��<�������]�Z��`wv���Iy�t�l+s�5��5\E�Zy�h�*��=E����N��85�X,��qoOc�7�P��(�㘍Y
�7��rc�p1u,#�dg���Ԋ@5��M' x(fYz��D�(+'m��/������!�T;�����>�-��Ʊv�a��G.EW����#<�%i�}���7��k�����@�4q[���'Қ��M�F���b%��c��.�7x�0y���� ��84��B�$	`W_�]+.��N At��s��R��ǈ���tR��Z��hy�M�.�Fv�,�](4�K�������	�,Q�.��[W����B�]�3Q�� ���U��zr�����,F��ȸ�4 �a������Ӏ� �����H�tD�����m�����Z�U���A��*�`�!����Ӝ(�.).)ײe�h�=fa2*q�m}a���*���"�є�u� �K�ǥ�&�PwRH7w���r�)ɳ��5�사�z��:Ϗ�S�(.'�t� 4x⁫�#��P���?G�+2�g{�	�'��2Q�/�����*c���s/��o�&(p.�նE�|�TiF�ȸT��`�����y��*E}l�H�0}�T���w��rBSD�F�vS�%����![�鎌!���=p	z떹Yg!�ZG<�q�T���"�$ޅ�o�{V;���"eT����硼S�k���
��D+�����\�hǨ�p
ԏJ����De�6���J��EƦ.rk��ec�aB=+f�<�a����� V�J���Y�N����)�0A��l���7?q�\T��Cf�CS6�����kO^v��W�X���S�o����q�/��[���lȻ�B��`�*�޿������);{����-����۲磕��K%���ߡb�Yɺ�1\)�H����Lp&|�>~�����'�� Ѣ�#^g����BU5�P��ƫv�A}�,�[K�F�}�0��Z�a���ia��_ks�SiCJ�n��v@�������&���@�-��,�nݺ@#�@!ٽ:�] J���'�G�w�q�b����O��O-�s����������:��nf�=����RO����	*��Da���ӂ���.�I˜���4	�4x]?��N]�o0�T����$�����\~7�
�5�"��� Ż����-1?1����s����Y#nZ�d���\�G.�B{Ǡ�PU܀XȞ����Z�t�H�D
�	���a�#�2��1�s&~�v�n�!~�y}$�����O�0r�}�1������NA� 0��n;��3�y%t2�Q��;RӜ{�᪯�s�G��� WR��������k�	���YB�'�RrBA�&������v1�3F^�`�1e�&"! ik���m�K�������	g*� &4%��Ho$.�ѦtQ�w�����eCZn<#/R��;^��;s�(_0e�bY\��VC�E�Ǭ���n���(�ǉi�������k{�e��8Tm�x��ۋ�O8w̥9Љ�s�
X)��6!Ƕ�ߤ+@ y��`�ov�l�l��ע<��{t>��O�uVޖk�&>�'N[gA��$[���U��?	�9M�� �7V��3�/M��7;����+iR����6��`8?�TI�e�	�E����e�t-�
n�i��6*��m	�Xp)�|���_�J޲ ��h���5�����Vn��t��9J�#�3��o}s��T��!��+���z�W���z�\8Efٱzi֏G�����v�_����vYA�mb�ʙ��72����}�i��gXV,C�܂����>Ƌ�;Ț�:�v3ŸA$����]���)�f�B&�!�<K�����3Q��o^�ڝ���@���2Q���Q�X����wm��X_�5 ��P�7��p-*VH0�#ʉ�	����=��UF74��sr���Jk����~;gWT�4�J)��ZO_�l���z�l0U��|t���ɋ	[�<�ϣ��
½�[�m���<�������N�k/ν�Q���(��{2lPc,��>J�Ft1Y�B�NJp)�L���~ ��¦����]޵��H�L�E��E�b3o(��{��E(��a;��H<���وr���\s�<N����)>j��&T�����lQ��K��U�$�P��b	��f~�q��ǰ\���]��q��G���hf�v~�6eԂԠ48ms�t,�׃���W�v��&/�SS�����K
*�WG������*ҡ��/贖��k�R�<�`�wi#IÛ5�d���(chp��D�u�K�L��a;!����_�N�l�O�1�AxPu�!e�����qki�Zr��UԊ�7�c�+:U�-�%����"�zd,F���L^/JgĽ�KL[iލę@r��N�����)�5���I�������N<bb���##�סdǤ���B�V%Bť%Cs-�l�01����w �CE��F@����n�c�djX�}g����"a�I���HG�����_d[���s�d'��f~Ye;LVڢ�8���MҴ'o�����-�n�~1�У~={sk���&�y>*7�I�:1�-�G�rY��<��t%[���R�շaG^�4pS��P,4�^7��7"��=r1R�r��R�-7CU��pL�TB)�3A��U�����ڢ�0�y�z�5^�����՛�����b�ych/�W F�����Gi�%�ܵ�����,�7q�T�IdK��4��H�)Nr"l,?!6�Ta�U*����r{�ɞpj��T~@�*WV�-��?u�zW�|!��`�&���ω�Qy�t��8k�Ko����2W>3S8;	v{LA*��5�Lvoy�q��}�I�#��D;��t[�p��Ef^7O
q�q ��'�/aB�6���M�{����!Ϛ�f���D�҈\�72\*�+�L�%5w#�j��95)�f&v��]Y��<`�D������ 5qљ�|\O�%YaP�M�mA�^b>�.y��x�q��iH��M[}[�Z�|�V��.�����h���}��֓�Oz��EC�]�$C��`�v)���!�#P�;&�i��I�@���@�{י-B�}Cl�k�&!�1�P�7_S:W�������������!x�>�!�Z��02c�^�X�}, �< ւ����yX��G��Z��B�tOӂe�CC�J$����?�����o�9�E��Ns�Ck7"���]-�/-�S�H�y�4:�Rՠ�<⡅�3Y��P�Qݏ��^	��p2`c��N|�̵�u�H�����ڙ�A�M����~�" ���F�5�0�A���q6����윬}�k�$p��s���� ?�2�X�ʸ+��6����U� }`iF����m�0X6���#����mIO��O���n)f	q\e�."_�iaxϷ
�$pĵ����R��./���0\��O^���~!�e�%�0��0�x��Z��lo��/��Kb���'��"UͰ���k�AȪ��զ���
o��+*�3ӓɘ��͢O>@�4YE���lɎD�'#ADDG��bu �E�S�40遼�21�Ώ*���w�9����v�ߟ><QZZ���?Ɇ	)F������_ !"u��������+�lHݦ�*�o5NKAm���1P=@�z;[�ݴ�/ٹ)1Z�P���o��n���Q�j����K�@�d���½ī���e.���I=��4�J+Jl�����(�r�K0�3Ʀ�lB���fǮ��<G�6c�����*���?$o��������k^�zq�7��?6��Hc��0�.fH�bfމ
��m���\2��ѐ��A�f����'�6�K�#�y�8>G��� �� !�4&>�s@5��)�fC.(�e*�uYs[Ϣ �e��i�S�!���ۄ�g�NOӑ�z.�������;��A%�#�*p��^�f���	�Ǣ��u�jEYν\?_��nE\���r�<�Z�<3K��S�<T1ݍ�=,ᒿ،@�|x5��)v|B��b�Gn�M7b��?��芬��"��jE�����T?Q�	�2l$�QEÖcLiS@��?��t� d(��!��a��k���L�@�v�����?�3��tn��|Zc3�xq#>d�=����+g�mw�\�����ΎR��.��n�q���rbCan%i����� @ @�󯸪��7��<g��ࠀ��WI�E���k���l��"@JI��K���l�5k�⏽�^Z/���}�8i%��2*1��
�@֩�~;j���(�;�9����Sn������f����n���7pU�����}�D����j!�*�����j�u蒰0���ǝ)��}��!��ȷ��c�E�
=�P�� ����c;�/aM�a�FS-T�6��?X.�BF�iQ
���c�<'�j���<�ۓ�*fQ�sd��8c�����>��3�6'O�
��*&u=����8��7��5)�����'I,n$�%Hc�o���Хнz��]���;���0�����C����R��c8P����N�V2cY��K	�F���Q^c��5�Pq[p�ü4���gNj�T�2G�$9~�n� �����o�h�9����f��^vYd�/�쵌��/l�gm�U������U��*�݅�g�2m���O���Jf�������pupͪ>೧�7��R-꽏��-�?q�{��iR�8?�UԮB��D�i�=�dnSY�y�o�s	��ᅵ�%ka�ߵGe��ؽ��l��U���&vY^��dP]˶7\�'l�k"���u=�Z����4	T~�cU D�����h�=�W,�!���Ao�W�0!��|����d�Ɠ��lC]�b�yap1?q2!�\z�]cҩ��~'���Q
pf��L�Q��U ���=<W�Tw�_����8u���o�����b������^����?�6�K,fEL��t6xx?�?�8�c�E�w�i�@�D�bKEK=R(��<x�����仚p-͒4�^2�^�Y1�\& �tT`�*�gl~y��I���{8{�dv>°�IR+W�	Ùy�e�h~M�Dd�kC��/�-�r<-�=8ꤳ�Z#.$���@� ٖ@E��LI-�J�,�Q3����C�K����<�Q����u�1���*2��S�+�:�}%��_����7�|�a��ޕ��ڤ𻭠�9%�х���(O�/��HaȠ��QG�������nM*��zn���o]1�$C+"��{l��F̥�*gŽX1.��=�--�P��0���q]��o�'�K;|\]Q|�ѐy�Y���
�&�ٽ��*�dtoa�<;�$c���j��"�,�<�n�0���g*�{��]v/(�#(��L�WeV�Ox5���j�9ea*���r0P�,ї�ְ��֙���<4�7wR��{����Ct�m�.�aN�u��	l�oZOn�7�I�.�q��f۫*B�����=b�������7�;G1�"$�T�I�<-��c�
��(g^J}����0�й"�i8��Vso��ow����-�5)�a�� �Т��J=u��z���p� �:�A��A׆IL����V����8�1Y0�����O`9%aK� =�_-QzA�ފq���5���h��sS(�9��3TY�4� a�ׯx��J����\��@����G���%@�֜Mf��,����%J��qS���3�G�p������MR1��@<j� ��:C�.��{�ic8���B�m�\��e$���>IIް�z�b��h%-�����6�(�+51N�Sk�/Yc�c0k�{�䅙��P�w��ԴC/��y�p�w��������6�d�O+�����-1y����}���.e?�B�ـ��>�ξ�6�.��|ñ�f��%�~�*�C��Xi������IMϚؔ����}�-�
[��T�Tzp	��7�t���������MP�=؉>7`C
#���~y��i�b�2��zN����(��XX]_�°�J�2���T��bk�MW@�X~�Ϥ���t��h�سk=CW&���k��yT��K�W	��4�.�)��Fz9"6ct�gkT~#�e��Ε�ed�ͤx�p4�f�$�4=�K@����#sNg�J���V�k=6���!?��5`o�����o��DSҖ���m����n��|�����ۥX71���/��m�f����;V1��3���E��|�')Rq_8z&�����I��~�NO��N)�	�	U�� w&�'3�p��xP҇@������&H�h׸����E��:*q��lU��]ƒ;�ΗM8��Fi���E^��ڎ�OٴS�W���CyȂ��%u�,u���u�`�Zp���
�n�͟4y��{S��hQN�	�r��vC��<ۯClR� ��� Ro����,��7#��V��o1L"5����YL���pK� x ����N`m��2�+��tǩ���o	��}����^�Ȗ^)(-D�EeY�Ooh��E@l}1��z��t�&V��&�
+��s34gQ^��%�u�S!L���<�}���p��Ͽ��E�#�җ�X��:�A.o"=h��]� 5��!k��������N$��zH��Z��^_���%��ΩŐ�H<䂄oZ{�1��4���}g������d�*J1f|�!v��T��!��C��
� �`P|��K�h�DE���f��ep���0Eє�b%�3Dcݓ@D�+♗�5h�����l����+%��kַ�X�I�('m��6�k2�b��^jT���3ҏ}{+x�'G*��n%��+��O.[^�B�����9�/�'�v}T�XI/�R���jW�SS�GA;e���2����o
��m5*�S�lt�I��,��@ �>S�Dk6z'����!lN9��QS�b�����8x=$���������ȏÊ%�Y�9&eh(�(��@j��Go70D[�LWK�uAT�i��~�2��ؽ�S
˜z�e�ba�ا�`ʟ�;�AT��S~��e���S����R!�|Q�K9��[P)@*q���R�)�^����� �n)�բ:s�^=Z�M��]]�Z����T
yid��(2���5BA_&�)�}�et�*Yjݳ�C馏�:���&�G3,���>E�����ޙ���ʙf�e��Fr��Q"�Р!��`9�������ۊ��o��X�!��Q~�q�ᯱgP��k�nZ��_��"�#^n��Լިdi��"�i���F2v�.�ð��S�����'z���q9�&J2�䒾���;<ҍ>X�+x��YU$E9tCg�O~57�j�|�\��+�ˣ���G�DۚCyn٩�s�|�{�J�����I�]� ��ΣĹNտ��A���}�s+{.9����mL�!T��E��RZ�TF�j��U��*!Ⱦ}8�Kar�z���Jj�CS�߯�1p�K72D��Ƥ�VH������~5�ɓ��dU�S��9 ����s�-ME����z:q����ؿ�p�XP�c�٬�;=�m�i�r?{�6ɣ�E[P=�"$��9���.v�p�����S�c8H�8nI�E�1�h=��1nJ��c��A��-�#yfw+L
��V#!Ȏ��R�ՙ+�r�Y�{�h����*��Gt����=�&w�dI�9eL*�Ь���^Ė߈�%��dW�m"� ν��-"{��@��"?�����Eزo�Ë<'�J���F:O��A�n	y����f����w��jO>�����"3�!��MFe���N�(�����j�%~�k�w����p�������u��AWH��%�2=%�	sf���A��fG[�(8�'��{o� e���e�u^�HF4apB���2������̈́�n��4O�j����S���y�׊��2,8���A������5��usK��;WQ-r�ZF�V"K3F�{I_�p�Mi&7�۔����c�n�0���Ћ_ ������H�5�F�R~^�)_�`�٬�0=R�0:=�lr�&��/�)�yȄ`�u���o�{/�V����cM���hM/�0k]�{�����l�5�
����.�8�5�eb�Zc�E,z�ܺ795�x`Ƅg�����O��yu`��a�I�H���(�b^-�O�Ԉ�7b�x���U�Q}�@�xۮ���]%n���W�y��1i�:h�aaOL7��A�s!1�+s$a���H�k���q0T��5���L,�DѤ�����׷��X�Hh�"��<��\�m�S��J���c�.������&�]G�d�����q�EY�A�0�hx=�">�`�2vƃ��&�Q}E |�/�ؙO��ҏ��%�6�U�1�"qU�f�g�>\���߁�޶a*{u�ͫi+(�s&��� 4�$��j����p�[�:iL�<@���z����d�T��,/��>�3{��Z�C�f�Ş���F3�7U�`�s��朖��*�)Z±�Py|I�G����O�1���'A��F����)��?��U��I�ӄ�OR�+$�-�Z
�Dq�B3u���3ջ�'~�i%���N[�u�Q����(D�]�tH�ځU[u�Y"}� 8���3���Ks]�������#�2�-\��v����.��v H�4��Bxㄑ�?7��ͱ�F�(L߫�셴�q�b�o��]��-�⣙�3^�=&F
�1���[vK��k�e��潘�2G��C��1���o�������
�8B�k��4<~�\�J��;C�n��i�}	�ʻ�fR):+�d}���-L���P1�O�E�xޱ)_t�cyS��@hd�C�_�ˁ�S�U0f��X��G$�����W�,�T�,�(��w�C�)/��b��Ҏ��-/��}\7*AC5�w�+HA���o��OuNy΀�S"�x�r�������r,�G��Ͻڜ�Ǯ	���L�H�7j�&
ƪ훆��)q�"~��a4H�y���s���M�S��h��٩��)����ǁ`=W��86���u��_d���k+��ú��z::�76���s�Q�(��SP�r�z�?��	2~@�ۣ�d�L�����;��{��6Ɂ�c��{寇��}>��rPjf�p�P�`�&kѸ��A�2�/�j�+|�g�s�b�9��������c�	�3{1�0Vq$�A�1���"����}�e�x�+y��-�D�h��ͅ��o�`�4߫BJ��=�_�*153U�V��}���-��2c�qW��0�p-Hu�&�I$����_E��d�����.�N���*�jhLK��>�@}۫"[�XC�2��ti�*Ip@���~��Q��1�������L���cy�2���pt5j��4��s�c+�r�K,���rtA�r����z�D�-��o��+&�|�3�;�hM|��K�'�s�}.K�5\Is�so�x���K���U�qpZf�tj��V���"U��KGX���L�w��6�e�����ӌ8����[��:�L�߻]L��$Y�4kx�2��E��M�Ԥ�ߑ�۝eVyw�������K`�To��y~��74�R�YFed������5�9'��4oHZB����Е�u�r����i ��x��j��Qn����J��A��6x;�a}�莄�S����=W,폝�°J��*�P�����| �|�*�	��B��ޔ����u�fd�	\����e������5&��< {���^17}X� �fx�Ր�,�U� ��5���Z75��%�.�:�	zf3*� ���e�DhfW��mI��D�'��ݦ5k���U詚�$�B��2Eb�dA�jf��`�9	0|'
�ȶ��a.�=cp Wv��a]r���� X�ƨ��z�<���@oO���f*	�� I��sbg���i9®R>�W#*�(3+{�뤱I�Or�,93E�jP�MW�𷇲�uqumvR1�*�H*bUKy�I!���Q��/��.;�
R��ąeWu:���_Z�>�g�2g��l���ԓM�Fȅ2W���X�-9F�3h��`yo(�ռN��c
�)����uTo���z�efU�ߥ�c�\\���:�r~�*�^��Ͷ����6MoZ�{�Ijar�?��cX���4br�����K!k���I|?����$,���wB�0�d|��sgQŕ���E�kd$w�*��Hl���;�c�)�n�p�t�~������&H�_M~��M�;*��V���Eb~�}�"6؀�Q��n$��X�ޠm��B^M���?����9��M�u��|��Bm�]��c۫�4^*���)i�U�z����K!j����[���B[em��#��3C�4�)S�?0.K�,�>��A1�#1l�n.�����s��F�ҩ���a����f��aj���|�(��J&<(�jR��w�ڠ���Лe~���-�8()]\U��o�}mH��Ε�[�>�WE����m}#��w��j�1K�N�oj~����������_�Ɨϰ^ ����Z��g^u3Z�bMB%U��/Ѭ_\��L�*k @����c�Z!'
Rb2�|M� νhk�
AM��kbv)�OZŃ�q-gq���
f���'��K�#�'�s�·��'��p;ﹼt��S�PuUY���]'�Q�=��7<�����
V���Vt�?!zV�IZo�N;P���ŕL�"JE��:��l���s 1�Yͼ�u�a	�l�Wdr����!?���_}�K��F���7��	k�c�8N�{������R��<��x��QYE�B��xh��N�,&��A�#P	6;��R���UmZz��?�=��3ڣ~.OU(��c2MQ���3��@)�B�យ��c#-��w&�=P���[c?���3��;^y�����ъJ�"�!������B�P�	�p:<��i�O��P+2��D������R;�@���>��8��k
�}s�����Ȣ,������L������6$�^�+\��V�i�O�}��ո�$��"᎖�'�+�@������}����l��o�FT��fGT�d�~�7[��̜�H(��=5H��	����J��f[`����T���}�/�.�K��-{�M�an�m�G~q��}y�F<����Ը����Ѯ�)Ĕ~j�Uu��/�
��j,�d�ú}!܀��)۳�t#���3���T�M����1���H��(l~C��`�lA�a�s谗V#��tݜ�'��,���h|�N�Yj�sZ�$��Ս��T5e,g��4g����ܯ��J|A��?V�&��fk|��������l�B;8 h�SO��G!��)&\�)L\IBn�b�xZCˍ85�K�3�Û�U1P����=f�N2��o�<BU ������JO|%gŉ��I�k�d����TL<��=��d��J�t��fi�J��o�mQ&�}���Zc����������7��?����(E��ao��Ӯ�w���+^ *T ߔ��T�X��f���,'@K"8�΍�U�5�ٖ0����k_�y&�	E|g��$$�"Xh���,/%l`	ժМ0:�A�J���eq4� |��9OU����ܤ�L�N�e8�g8�%xҩƏ9LS)��ԕ�2�/��"���]�Zd�P��wfCH(�s��y\k�w�
Ռ3�M�4�iP��L�^�b$������QU�� �އ������橲��A�,��*`{EJ��j����!u#,��\��Ƈ�ҸZ��t�Q̵bmb�c�حg�&�a?9��v��T|�$��Xh���-8'����w1�ⶡ���Q#�	��!��S��Y����{3�oC���� /����n�Y��/u�[�P+������ �;j	��0$~o^�Ȗ�&�&<����X��yߤ�e��!ιg�a��ĉ��9�ݗ�ޤ;��\��1����O[Ɇ@��s�{�T|(ՅǓS���ك>�Aq���E-��ۧϛ���W�2�#Ѳ���L2pDIhd*��%�y���n��A���������������� 5�Ir��>��	�����E8�$�Χe+���"�FU��˹����yC��OI�A�K�Y�Qu8���n�~�L��`�� ��2GT#E�F}�'���\���eTէ�8t��=�V���sg��,d��.��ћB0�ę�ڇO8l��R%�1��kp����I���5�f����L�t�+��bv�W<7�4`��>�d��i���|�5�ni��d�V�^�#z����s���Ϭ��[�}ʓ�ɻ��9�;�y�1L�b$���v>޷��cRŵU�~��Oh�+�~��KW֚�$|�CB����L��Z�B3�}Qt�-�Ȏ���\%R@ГyBײp��bZ��}�����E�\�>ĵ����^����	���D��%!��Gȅ-GAgQ�~H���Zx|�z�n.O��),
�xg�K�y7���i�ۻ�R�S�<qe +Z����Z�����l�I�5(��{�����I$���)��GX��K��*z&X�(�����i��.)�.w����L��eW�'Sy����m�D$S@NF�*�:�0�������Q+x�f)�s��k�3�&�|qi���D��f��H�q�C��s1�͵-�Y�'�[��	���
�2m���ǆ��=����3�E��w�2c�X*7��1a@_l˿���^�O/��^s���� N�?2�	2�r��P�V'��B���x���ٌ��׿��kw.Ћ�٣v
:����dc���°#�yfؕ�ˈ������M-���v��Z(=b�K�d�㩁?8+R���6�t$�h�U�_�َ�Z:R�o���h�*��[r�U"J��P��v)C2�v�jC[R�����B�N���!��~Wm�|d����
��-�Qn��"����nQ�~):K�a�W�/�l���lJ2F��C6QP�"�ؘ�3��Q�pY�X[�h���~=E�ʙ&��ə�㬈u��.7�L��ǫ�BJ*��쥃6�]1��/�@v7�"sh2ھ[�6�pC"!���H�[���8��s��[�H�Qx~�L���npJ��橖�o�צc5�]��~�N�ad9�g���b0NC4��xjY����O���xy�Kz��nzޡ�|��I�Ož��1�9��tv���
���C�K��q.	;|�����^�OSj�#�S�`�Hj�Yd4�yƧZ�8�	�6�{���H0;�Xq<O��\,)c�㹅=����s4h1Of��6?J�,v�Y��p��м 0��N��t�;(ۮ�ܲ�/ks�������P�)�c܉D�p�hs9. ϊ
����J��/S�����
\�&�[t-��N��>.�
�ee_�"��pOاA�'q)E�^,mӬyډ2��N��ǹ�h����5�|���2�e;�����'|t}b�"��J�yn��l�l�0�WMZU���Z�i�����z�aMԖD2XcC-=.�}���\�Z�o�:r��/x�1`��>�T�1�������?���Qs��D!R͉&y�u&ض�DA|#r6K��{��9�WX9��fL�̏���TE����zٔL�"!줏g�z�x�>��g�h�{��ȴ�c�g�"F�+F��ĩ�3��p2��}�����}_�\Vs���x�B�d�����;��=��*��Ɓ��q�i��*2,��6�Mg�'Q�M�K�h����������&��o_��5������l#j�UpǇ������R޾�Axa���hg���qwG����p��C�s�o��˾�����o�0��h��|���cX4hj.��x���)
�n{8�	s���B�T�g9�Y�	��E)D�]�m)�.��:��M��:w������5Ăނ:��?֔����ĥ�b�����>�zgx0-3�����y�Ɗ��IqA���Rl��J���8�+xIR��w�P��8��u[��.�uL��\��I�K��3�&�i| !�����1�����C���]�gc���ݽ���:��l�)*r#|<l���j�8����z\5m�*ʨȪ"��o�$M/�|�u�Ĩ��$��Mк'�J}���+��r�)�\D���̛�1�rH7�����4��k?�k~\$AqM�9MO���$������4g��#B<�nR�I�|�J���#��1���r(���$�����H
`�+�W`���W�[|�q���Ǧ.��:�k�����Nɇ�>�BB��B(����|-L�\�9��x��]��vf���B�|`�}�搼Ve,dڨ*��D�A}�`L�9����J���d��4J�V/[�����?hG�}����K��~5�t`"=| ��v,̗�Ç%�����7�(	�n�]�������h�J���L�}�=/�p;#�9���7w	��|���6w�V�Q��w�b���G�<hz�̈́�&v�fhIzu�*=KIQ0����}
_Q��^8ʴ�I��~��(0?m�F:��0��L�Mw����08JK�w����Bf$�`����S����� �c�HliD��$��~��C# j���?�>#���m�����F���-]�CyUr��UAa�
r��=�l�ɳ��L^����p�\ϸ��X�hNM\�xI�~��l��c�.l��Y\n����c1Gޏ��:���_eԹ�9��Ey�3�Z9Q�f�v!i�ٰ�l����m��Ͳ ��n�6A��T� E��p:[.A+A@Y��Ve@�89$7R���i�ں��$�m���G/qR��ޛ����ܷ5L��Mm���J�}�Zk��C���:w)�zT��V�C}Z:����Q�+�# ��'���!�VdhN����G4�(82�]Y�^M��r��[��8�D%:�dt4E�������u����$���Z�5qTz>&���ry��O��MM�~ua 0ۨ�̸8�Pu ��s��P鵬�,9j��$z����L%�_}S��" ���	r�����n
	�ߡh�l+E{�.��2��C�cNf7�<�^F�n��畷���.��0��nQ~dX��Y�Ɨ��B�3��4�-H�M�w��i|sZڨ�D��58���h��hX6ʦꛧ��Av�y�� ��[j��(U��'xY*����c�2` T��R��.&�Y��X��%!?�%�K��	���"Ϥ_�U��oE|}�0�Tmx�s��7Y�:*)_��跭�o�֟���T��Q���jzvy}'^��	}yG����������D)���1U�
c��{�"B����>�~Nw	p�1)� �K܎f����B6P�~FU�|���q�/F�kr�Ј��r��9�՞+|N�AS��Q*2�`3��]qJ3q�P�E�m	d��%j�j��F��,E����R]��m˼��+�ck��z�����-��D���W�a+�pX��q\l��֊+:L5\\K���[<#�;�����PE�:����3wჅ�st������{c$�)���k-��[d_Ϙ�Wٵ��Ϊ:���)F������Ppԫ~Q2��t�0hay"��R��+g��I�}9�E2���Q#�S��]O�t���{S+�پf��s�k��U�:��^A	O�e,�CB���^�� 9b���Ì�?��,��:�Y���l�^;�4�5c8\�����S�0���6!
�i�aBޗ�<޸�f�(i��<_G6��gl�A��;}��6���ڳ����N��Z!Ker��9�DYu�X��M�����Δ�vA���x�Re��ѷ>�C�@��۹}T�1$]OG3v���W��R�ys��@���F&�Hg��N[����e)$P��k��.Yb��.[&���5-C3�A�B����P �^��$0�	�D��d���C�g�O����~kYc�PT�K��1դ�ig9י�l�1���׾�-[=ٙqmZH���)���?�L�qb�H���$� ����fW�@�����#�G1!|�R��/~��^h��IVG
�``%o��db�%oK6n��z���RCKf)9iܶ�Ӑ���k�A�c�TƇ�2ЎvOl���B�:��V)�a��G��<���\SjJ+6;��NT�x�O��+r�Z}�5I8UA�%�]�RH�al�r.5�C�t�͓Q��$��Wm��=r���O��y���N�]���f�&BNI�!�f:�y���Ŀj��G𘯯p��)Ҍ�r%�1��Ёx��"	[��VF���=
y�v���ȅ�:���ق���I� x��6Ѐ!de�7����������Y,~�pӻ�3�N�8�|`�#����mU���^�&�B1�A:�tR��3,_nO�5�G�m��Pg��_�t's߃6��c�ߛ����;�� ����p�<�b�[�֣U���+݋�%���ؓg�ì�C1��QxR�)Ha���rM,�r�MH�F.��F��G��([J���6��7������&O��d�N{WB��J�� b�g����ϩL��W�*���q�e.��l`R$b���pm��Ђ���˔6�䞆��V����fGyn��耍'96tO���)��+���Ғ�i��� �nm���u��.L��w��b��'{YSŋ��OƩ������W�O±.�${I��A��e vDVN�e���b���S�gO ��<<��d��F��<��N(L�mϜ���R߿v),�v�q��~y�agՕ�ȳ��\��*5� �$�,��|��ٸZ=�gc�.��t6����D���p[�D8��Q��c����Jj]t�ᴋ&6"�����O
+N��΍l��ok�vz��mȽ��o�!";����K�!��PeJ���&�xH����^�Eop��lZ������F����r;�Z��P���2���Zr\<A;<�T?�e����-�;����̿qZB1�<��P�I��^5xT��wi��dm�����M�+�����rg��K5�<�{���!^Ahk�e�,���, #�le�>�J$����֚<$��Xݶ笈�1*M��<e�.�zڤV�O�f���g��J��8|	 �K��lX��P�r�f"X�8�����ў3�e� ��"�#�IH�^'�����v��T�5j����#Ds����Z�$T�=��K��h���d��Y�Wk�(����_�K�׼�ͺ�	mbh>?A�J�#qɚ���b�0���᪬U��dVWa�_(�~����N��6������l�N�Ό-�Ҽ��}M �QB�p�wQ!�R��n�ʆ;���\��{�����mva�Q���m�Od��B70^���#���A#��gI�M\E�W�z�j:+MQxx��!�o���ȶF��@���ga��G��'/V�=��+G�a  3�����6���D��M@C�1� �P(� <z�����PQ#)��t�pPBZ��h~��|f	�Pz/�����u�9����˹�1^�������\�K���[i��-��!�M�_�I8��j�S�d��t�s�[%�q�zGy)]�Ɓ1��J�٨\���7 �:�T2�X�D�՚�G��s@�
��jH��m��$k*��sK��٦����1�����YqO ��:gD����
�2$Xuc�5^��n��dâ���沋���#0��;�<����)��/�Ͳ��Ab�њv��☦�����~����R�D*M��q�/㶁~�ZN���Z$¼/�Cc�s^�e���[̫��zU��i:��!�J8�V�yח �mU�nLQL�c��!���:�����)��56�&%��u-����cʳ�%��t�~��u��o瘣D)9N��9)`���j��X�0�/]fhZJ��p�M��-!DNVC��n�ߗ�dx )����>��Y ��O��͜ct�Ϩ�������e�CD�Y�s��>n��6@h�b涉&&7�*�{P� /���'UAW����ȝ�����ܢS�
Ky}b�������"x<_�.��`�STXS���;L��K(Q��=gP���1Gb��W����Ѷ��R!��}ň�ˋ��4\���v�+���^M�j�	�y���4�N����i�h#y��e=j���;'K(-m���Wql5��1C���j/\vM��ﱭnk�Ixo�R����^iWMDz�|(�1�+��e��T�wT�@��9��|-�F�xy�gD]Q��eL+Qy�^���z���R=�9��5�d��ۚxW�h?��:��L=g��ۣX����h�;�5l�����E�y�m��>:�`��
��&�N6���nΥ���������eyU��Gjt��W��U�	2O�����p�Ge��3�k?�Dͅ�Q�<��X|��)cþ��=�&~�q���%_���q\�����,4�MaFJEr�9���P:�&�ye^W���¢ҝ�����/n�A߸��Bݝ��|�����
��:��o������!�>C7%C\����y3gx�C���8��TQd��U�P�G�k�����W�$F��m�dxQ/���<X��r�,Ө������~��ɘ�E�z�F׃I2\2\��}յ{B
�����A��O)��0q�Np�3�x�قAOI��R�K��^s���:,i�e6kE��j���\9��͸"��>o��궛���@�T��	-dK6)�q�+����C8������j�6 �(��X�܃M�L�0e��q`O���8t��9~USćF�i+L���߽����t85kD)]� ��"�ҁn��>bQ�ep�#���N��ƣ��������T`����mɢ+Wb�
�&MD�tͼ��0�G���p5H�j��Y�\@X��GG ��ā�S�C��aa��Do����g�b+�1�����������oL��MNb�c?3�Zvj{u)}�&���/t��q/��~!�&�,,�Sy�{��v�����"�����}-j➔�39͂뱺�4��!�h�d/�R�Ȉnn��J�Lm�A���S�F�A$������$}�X,�I.hɪ�����z��S6G�9��c�T�P��r�E��C�~�v�������+hO�'���H0sJ�32I}��).Do.�"-/(4t�qGu����G?b���QmV��ZUοLX�D�m�QG�`�QP��l_�;���6,	� �^�wl��!t�����&Ŷ.���Y([#��
��&���W�J�چ���_c�Ae_ɕ���=9胨Ӊ��u%�6T��n�2e43�bQ�W��i2�vH�A�P��z?r���^��ElS�;O��vi���?�)� �T��~��N�Lw^7(�P8sS��و�I�?��
��٣��lkj ҡ����Y�Upe�<;!������=%D����d5ѩ��l�����5��7�Q�|\���\��-N^���)s���Wv@�gO��Z��[x��LFv��^*�I�)�*T{�7��(l��5�u
�vB�<	��e���ji��)e�N���ƒ�S�!)�K���^J(���0 ��t�}�M��Et���'�+��o��l�=�{�b�#��s=3"!�8���[�Ւ�`ڱ�zh�05�7�F�������\��s0�����F%��Yj�(���A�0� �K@G1j�'ז�ì�1��e\ �K����r؟���^�)�BÞ?�,������=j~��h����MUpC��Ur�e$Q!�-�y0��lu��bO �q�Ih̺QL|7^��%L:��q��T�&�z��-�����/!1�
��A?*��&��߸�_���o�����)x~�!�#[�ŧ�灜�s�ȗ��#��
B�R�*'���߾�	@e7�0MNĶ���
��ĺD��E��,��S24��B�0���V�(B��4d�_��Mr�T�a�+ON�����J2�hF^�=D:a����.h�Q�"H=a)�X�N�l��B-�i��At^�6-��~<M �b���K�� �X�m�ٙ[oɑLr߫�3�m�!dؗ��vj(�DVR}� G�:)�
(Tވu���rC҉v#������m�:��뉽���* �!�����B�z���5���8��V�#l�{��Ip��m����_w��{\���CҫN�{���rK�������Y�@��_��0/��QrA�|���@ʕ�������p��� �bz�Q���<'T�d�`�c�H�*A����eF��%ܪp
aKK�X���E� �I%xT��W�
���6д��a�Э��؅g�,���-dV���O +�S���.+eɝ��_�C�s]s�C��`��k���e�h]�h�-���O�`*3/^�i,_�ɏ��Ǵw&)�]��F2)���j�Ơ8!_2	|@�!���2���'���z����]N����c�
����-�͈Ҙ�n�"P �{S( ƿ��dG��/��.��� �g�3�*\|�sT:��`�����H��2��͢J���x�xm��D��N�}����OP\	.N��+��g��U0EM����r�Z]#sw���n�9�;��%PZWR�3`��������`l��rB��b�δ/\T\P�o�r`%�C�������R��"rO]ĕ�e�A��D�!��_���\[w�3�"��V�;3&�"4*���ܑ��
��w�OI$����Yi�`4Q�ە�o�+m�o�f٥S��-�F#RL9���������>'��gm#{F�H�&D(������'M�D"��so��?j�9p/|ų�4�ٳs����km���RQ���(x��r��5�7FD�r/�Ȧ���2qH��/�0N���l�j������'�J�`|<����
hn�r6;�H�^u\D���
��V�x����=<���s�����7;T�̰1�hi����6�i,oU;e�ӃB�[�'}��'Y�c��l��KT��y�b�ވ�*~ޔ�4�_?k��z��u���t��6�ŗN���s�+F��� ��C"d�|��Ұ=�4��m>��r;��4&�H����c���Ս���G����ڮ
,����p�1����R6;�`?��7����(�T7�bH��ޤ����o��v;l�Y�y�O�� ��7��x#�XWc��C�<$��W%�����xˤW��璩{�3������YB:�V����~4��F��݊��WV[��pf�)�d������"��@T�!�{>��xn�Kr=��Gk��/kUnB��8�+My ��ፙ�ͅ\��v���?A�N �!ŉf]���76�������v��� �+��~w-��]߅�	���J˶����*1�W��] q����f���.uI�ZX��d����7}�ޥ�h��G�n4��gu�?/���2�פ�J�=��Mj]j�m��3`�6�累���<Y/S�V��u[�zd��?�/Y�ޮ����?Ȱ�ŢN`Ve���|�H~�S=|�ʣq<D@��~B�?C��[�ʃ�u�|��'Y|��٩�y�����v<A���t�M�2�M�t���9*�x|u�����1������s�|1�����#��%vq�t[����2ۘ\z����xeqĿ�+���ؾr`�kl�6�s��d��>�,̧�gzK-k��4m��3zo%^�B9�`�6.����iY7o0�V�ߴ�G1�WmX�ӈ�l�wi�:�P�{�=�3�6��V��?V��_�iϱ��HܘN@��*Cellu��DA����*��ҡ+ͼ�M(\��ׯRf>7+�ޓi
0�U�"&��y|A
�`���ny�,���H��g�%��Z-C��Dy�LB�/��_\Âx��&-LԋW�%��C��rJm�ť�`0B����i'�!ZByr��H���#�����j��:)��~��z�/-��h��4del}]i"U"Sf�H
x[%��S�8l;t6�95��46ʬ�icb���ۇ%��ˢ�u����T.���v���7��v��t�����"'�ޣ���aH�S����]���W�sd��	��(S;ʡ7d��^���f�Vʡ]�-O/��5�7��}d*��9���q��}�s#�|G�w�
� 6?�G���e�����5.�>>de��Ώ��n�`�*�w�Z�*�e?���B]���Z*�4�5\�`�r��X�J�[4�L�Υ��&.	��88�FN%��a��:�L�������:��D�2�Ӥ�=�K}z�}x�X8�7˿X���#�y��:>u�!"p٘����_c���yיꀄ9F�g\15H�].�)�N����K���������9�L₢OU'��F�BQl�C�X~���x�P?�r���mS.���Ƌ(v�/]�@>С븱V��>.jWw衲<.���f�c{.�k��$�n��p!em�>�`���۾Ĥ�-���'Y}<��T!�VE^�u_�	0ܑ�O����.]`�q];
���j���.�^�����"7^�!�(-u=w������h�`�z���d�l۔� �y���\�wbIX�J�S�}��W�t�Pn���[�z�0	��zSP�T7���Bi�Ś�&�ٸh
U)	�b8����3(�e��2c.�j�L��Y����QmG��G������
�Jh>@_zI����3��Z��Hv�Lh��t�ܜ��?gX
�:�^��{���8!�t�!aAz*�[?+^�\{�h��g��6��|v��Ճ�b :����"��nl�6��l!\��%��q�;�.|^s���t�u��́V�ֲ��5�lg����}�t��k(d��0~F�]���|I`���a��t{�`�7�1Eu6{&\_�-P �4Q�X����e�hƶ��L"T(�f�Z����oه�e�����!��Zf�>�J�"3D^5�K���o��bE-EB%uSK�y�i��6{�o1��Y�9��J�:��?S��lp]ص�.�2��Dt#���Ƨ�ao��Q�޳�DQ���o/:D����׿k �m�c�Q�J�#s��u��f#Fy��x�8"������u��~${�R�1 �qt?h��)qdެ��V	��Q]�{k��~^��q�jTx�.�C6�u�����t��:�:���m�W|��g�=�he�8������o[o0��oӶ�!���*��^�[�]�Q�+�&��H.vH������xN��'A�Ǟ��\b˛+�_��m�F��##�f����9lՒ�o]�:r��p�����|l�W�1_c�Ɠ֞s�a�pnڄwJT�k��h��,�~=6�]��ka�y-�ܰ9�!�q��f�ʃ�Y�0�R\�;�5�Sbo/3�k�F�����(�Y�:��ᗖ�W��"T����69d��?��sO����C��a��3�BK�1n\
X�x��͠m4̌ކ�Z\���#�u��/g�����:B�[��}��1#~����p��D�s���v7�^���ɪ� ���ư�JNބ	k�о�}l��1Gxc`U�IjճV��	h����S���V@0{(�PiP��D�ݬitq���4| �$�d�M��sv�A���3҂0����}iLXЖC�a+�ͺ���\f����P�%���SC�l�$1��@����w��ĵ��(�zJ�������I9|�+��
��G�<�o�s �C�Nnj�à����|�P��n=��2.�I�����������Q-G��t9��	��@���@3���W��]S�x�P4E��6�2>1���zU�K)���!<��~U�|Tc�������hg��a*s���n�t�LrͶ�FA������/kw�BWh]�-˸��񓅽��n�Ç��j��D�OK$}�9:�$���b��*�XB�G}E�<>�ԟ�7��Ð;�Ϧ���S��(��Z�'��GC�&��dVi��kR�
�M��J3?�ּ$��m�CM�� �ն{��f�3e�j->1�v�P�f�;D?HXg~ �����g��/�b~�)-琝���l<K��e����l�\��[c3l�^6�˪h@ �������}t`@���A�(���5��������#���:�����:�1ޢx}��|M��o�P�����
��$2��x;��o�c��j����N1��+Cs	�:ciAmҤ��f3����R�>�]����i�K�aoQp��!���>J�N���.;V�9��?�v�=f�o����{�;�A���C�E/bh_�E�|������iD�G� k�)��h� ��ra�6�'�� b�q!E�:�ʹ5;�q�s���8]��@��;�9G�R%�+��L�ݱi6E0��]lv<#�K(�W�r�}p_
����%�8�%�I|0�r�;�A� h���TԦ�-�kh�O&`������k
���cS�޸�ɝ����J`ڛ���TaaTș�Z�"@=�@�����Tr}��{n�(�\�A�܄��/��i�K4��Q}��qj�Ya�b��|WV���k\|�a�]�
�Q\Y�[ѭ�c���)g�\:��د�/"�9� O��+s`�"�hR5|w��ߚ~���/���{��kRK�@#')҇�=��g9�!;�o_J�ЏB��AᲭ�H��g���z!L��$�|T/�a��gw�ye�B̋خ6�@3��hؕ���=���\_�m�jRV�#ԥ�%Ij4�Կ�<�b:RA�B�LALY��h����+7Ҕ!�&;b7��TSϪ�v�
??�8�C�ᡤ3�5 ݥcb�c�M��6�0�0���;{G��'�WQ����.���QPG�)W�Oy��4����=�{�~KU<v���#̮�!=�?ſ���]X���Zz����O1�a�U@�H�Z����+e>/!�ܲi�S=J�{���"��H��|C�(�qs�N�Ʊ�h�־P�؝4�'�����W1��e{�����+�i����Wԣ��|X#�:�O��bmu��e'X��� �v��cb�nv���
�U��j������� ��D�Jn�7�G��0���i��>�r
C�Δ��G�]�զ۔KgIvѬ>5e7�u!Y9�U��8&�A�Z2ƪ�2+��Qvf�~�`j����\��tczꠖM����҄0�t|M�UW�>�XaLm��W2$:ɚ���b�O$��?!�rVWç�:��Ȼ��Y�(+\��7\�^cփW��֥��#����\�UC��e!�>�	 "�����Vf�FR%�'}z�cȡU�0�������\1c�����p�5hf(D�W��7�#0	��~�k�r�?��9�W�[�*ɟOx����j�@��������nDN��i �B�7�WHDκ<z���M����]'A�L?�n�O��m�������_�j�S<m1��e�����84�ߓ:����|d�\ 'u�4cDW6:������{��\���;9q+��,�r0�d~��栖�U��h�{�/���OЛ#��P;�Z�6��
�]g�o��IkV]ݻ bs8 �M[{� ���t�*e�C���+aԬ��Q(�����ŃI1��oO���!@���<=��x8�@��T���V��}�1�������ĴSDl���?��j���`�>�&�˷������[��ۺ�I�˛�I᩠��z�B����ޢ�L��Z��b�p��E��V��zмO@i��2�p�毒�6�&��3ؐ!#�M�VnaީU�KL�Z�b����� 1ؗ
�ra����0��Y���{B�U}f���7�%z����e9C4(�r�����B/"��4��OH56/2�Y[��9u��O��Z!��^�@_ѿ�P�ݰ`�*��	��J�]�C� C8�t>�{q�R1��IYyj��,�c��>{������(��m��I����R}x�9*O.�l@d*F������I���$�ELB�;�ޗv�yG�y�k�C�Yˊ5/���S��H�f55ۍ5�e�H=���'�s!)�j��[u�����N9p$u_eN�D��i_c��E�Q��
��:��F0��J��;�M���Lx�����s� D�Vn�E-�+p3�1Yn���לgj	;/�φ
*y�X�\�[#�5:;g��l��ҥ�`�P+_�oG��a҃]$��r3�,�D�kw�Ip"����Ծ�r��Y��8�#L%M�]C�U�V`ߤF�:
<�|�������=�f�I��A�"'م�;!Y��(�iKv4 ����lo���G��e;^�����8�	{5r��7�A�V�:A���D�% ����Ĝ���k@ߠRH�g\-���Ʃ"ښ�C5�=:-�R�����1?�5���'z���r
=8�j�N7�{i������u�_�;5�[ٮ+��ˌ涁�!$�Q�߱�B6����?�_)SRMhtZ; 4��KY��*Ƒ�״:�z�uP��~Tb��j���趹����E��M?�K���9��f���&��n���Q�)j~�cc	!���(� y��`ς
*u��a�4>���6����h��;��#2l?rCW��"X�^y{��T���P�V7��'���� +}��B=�1��p��N��}Z�\�l��
"$tU�����U*�[�V�P��^�ڀ���.cUD�c��چ{}���٘�ȯ�{�3�X������>i�
��"��H�?v@n�0�#0�T���|��C�����ȑ�#B��7IΖd��K�ʹ���
ղ�?���4z���hœt��jQ{��l�:��ؕR�"L�~�&TK\ 9�g�G�v���')�Ӛ���z�h2��dpk��y�G<%�5���j�E]a�z�q��	�ᧉ������\5<��k�1�3|�y�m�_k<�Vkp�(bugx��W^<\�O�xO�h g�ۼ#��RdR�,m:q����#T	��uP�ƪ�4#!��`����&J�O�|�)�s�Nv����(V
VNj&���~�Ax[E5�d����5-�<���iT}�>	Ġ��Ą�qW3.����2�D 
g�@��<�;�;�!b�9W�j~s��p�C��۾�&t����M������*�v`(ɡ4[:�$̖�&L�l����vV]�IX,�����z����X96��S��FL����>�:�t�C,�)aˁ��`��gK#pÏ�n������.��iB�?8Y�i�M�W��ph�;<��(i-�o�H^P�����N���߹ͷ����>����ml��|$d�R	�_�x�(�6��XM(�m�v~GpR�5 ��g�d�M�D@�7'��=g�l�7yq(T�oY����#�y�i-Ƹ��W����W�v��t�1�D�Ҧi���e�Z��y ��_�����h����Ӿ�h%�i�s�ur��y�/l�ҏ���	t�Yj�Y�3��5/^Y/ԜV�n��Òu�Һ����T4�W�QL��)���Nc]��ү�d��O�PY��=XH�Ms�>�\��8�Ztq�rכ=l�2QfgQA���u����&��xX��'�Z��|�����w��t}Ux�A+����C�5� U�ʋ�+��h�1.�"bO�$f��Jv� ƦmWƱ����,Q��>�q��x�:�a|w���h���α
IDK�~�Ԧ�͆r]��^k�,���`)$�����fU��1ۑ���E9��X({���i4v�6�߽�-���-�٤�ȡI�s� Pd^.��s�:[Y��+f�$2$�v� �����F��I��3�:���h�G�K��vN�ch���1��if�6`����.�����º'�'Y�e���E�&���g��/�І�|E�&���­W�����X� �����U�& ���t>�@�S���vjt�2R� ����h+��h��Y���4�.�1�>�iH��g`���k U�\�28ݶ�T�>*m2����Ù\f���+��mg����`d�L8'��1]%
�a�t�MB�ˎ�MH��7��hPG4X���!�p'�P��*1h��2�oĸ^=�"�[�`��Dgc��-�j!	�邬˸Pl�5�-��8�!m�{�?�^pko�w6ڎ��.v�5=��o%�㜼�?�& �=��WXIn�k튧%�3hPxT1�oU���iֽ�>c� �$��X�^y@Gcˏ.�F-�F!kaϪ�H���A/*�*O��Z�YgU\V)�\�y���e˷�ض��J��1a�s<�/�g��� �����T:+pg�LtvĻmq�2�3���K[��g���!�8�sOe��3|+M&�Hu������ca���,\f�|g���a�����M	��ᒽR��%^SJx�iI1�:nx3�̖Z��(��K�5�qٵa���U���n�s��#Ʒ��w�-�c%����W_�G�*r�XE��gd�8��Q2"쓂&؟����s�����ꅛ�~
�1_mI�1�o=*��O�7��5F�����^���.3�b�y9�.�pנ�S���(l�o����o8Gפ���Rc�3>� ;e
�{cŐz��4Y�X��i��xWfS�Ea!��EC��b�%���:�q���ȴ�-=�����Έ�'g�� \��#a�ؙ��%M�̟��Ĭ�z0�6s�?c��CR!i�?��$
�N-B��5��uwh�Jgz�3�B%V�9�g]jF?}O�Ž X{׎I��"���"3�Q����3P�빒ϯI!��Ӏ����
%P-���ұDS[)&_G�n��iG��O�n�?���'���p0S>;4c�|��f���e��8���߇._]��:����f_�TB�|�#k�Yɋ������l��9����"�@�#��w!��w�f�������te���p�H�&2��������]>
W���	�+�:I�0Ґe�Y��uF�1���w�!�h�qPMd`�˞4���d�rFk��Y2�T�x���S=T�;p�La8<�9}T6�~���h2��%�ǫy�`�Ψ"k%t���N�"��\�*�A���>�Q���U�*��:m$�E���S�E�$l��hx;[���;+�"|p)1���H��1�x�/��U�{[{y����dV�i}�HA�[������l#��]��Vi�X?�t��T�j�#@�.E�Њ���3$O, E�&Dֆ��|sN�~�X8>��Zd�����~C+�\Wi6DSz�Yx��nr�kW��
�cyTylw����(\�^wh�k?�����2)�sEms��ͽ'�wǅ�.�)$�Fs�%D�������H��B�D�v�����c,���i�t��ja5���5� ���~��-�s��þ�]06I����|SX�[<}�u�R��	�	tI!pD'^�t]�6̏ߖ����wB�8��g�]b�O�"?c�+sv0w�2�L�a��R�7��N�>�Jg���C%t�<UG�?�Ӹ�"X<���W�U�
2�����c7���s����n9����O�_����#D�5��bbx�9�K�G�N��cKT�.�!m`z 2^�c愪i�&�M&���<�A��|���
*��4yH� H��G����9�X�3L�7�{���4��o`��ޞ��Km�uF���a���H�\.��8Ug��#��'2��.��G�}Ê�(0]���3��~jC	#�D۔-ɜP�X҇�N+��l�E����ʸ%bj�C��)���2�`��Z���ᆩ�wGa�r,����o��安e-1�'ڋP��59�^��%V�c���w��n�]�D���]����(D?��paK1�ƓW��Jn�'C���"����g~�NCL��aUc�0e���y��\<a����&�I>���}�� ����u2zC�fr�e�4����k~��"gf��*�� �V�<
�JR��v��c��&������	��b	mD-s��n1��m��(���a#Irk�ݕ >�U=��Ӈ�8��$�c��G7;��, {"7���~��6%>.��)YnW��(���� ,�an�&;����H�A�K}HE+$ӊ��ؿ�z�.�;�l-�p�i$�M���Y�Oq�sC:t��Wdqlj2���5��e����^~Q�ŁE�V��P�9�#��Z*���i��u�lPj���N��cR-����?���XsvC�Q��w���q��e�鼯�fZ�;�����e���;k>�7�t�x�7����"���qj"#�ѶO�[F�����<��;scnE�������Z $��5��骡TM�Jw�7/��E��7�g��\5�Z-ZG�_B�Q�>|v���c����!���&(�6o8%*�eO� r���X�1$���$�
{Zȍ��$.,H{bl�/:m���y佀O�E�ŹRAZr���0�VH�կ߬��_�9��|��Ż���4i�U����*�;�qQ����u�\��k���&���m�.S4���������Qw;��KZ�c��[�9 ��bp)#f�6p���V~{����z��ȫ�q�B�x�s��gLW�z3�v�=���-U��<�/�	D�r͕�*��!>c�Ar� v�)�y�8���٭EE�i��I�?��r%vfᲐI�d���xR�ș'X^��}/��%	HP@~�C���O�١�sgp�؊�N�Q�IF�t�?d�h��b8��F��Yùa�2@�:sMKer�E�^��@a�߂(���2N�r�ޗ�i���g/���}�4�/$�DϽ�|�����>�H���>�F��W!8ŒOp͔y}񊡂Y��Φ�"̢I �J^�#Oߚ��9G꺁+�*/b�P�N�#�ML���X��7�y�j���t"o����@������hƲW��&4�u���=��z��&ls�to���ꚁ��>`��:?��л�+1FE�jRU�u1���AMU-�~�����k��0^~ ��@�]e9e���d�7	df�v�3}�O��r�bߟ
����EO��rKl�/�ó�uͶs]&�X\�r'j͉���;�\�XC-��z���S;�~��^��@} ˘�섵f���F��e�	3y�
�&�"����p���,O[������7�N��c�^ >����b['!�jּ�H�j�=�8����ħ�?N\lI cџkD/���g���ǉ]y3C�o�EpENH!44�]&7��3�S�N�������?����f�Nk����&�X�:XÑg�dl]���mF��D����������=ӷ3�ѧ��"V7̲����0�ٮj�TK�uڜ��c�`r�;�쬁U���}h1�Р���?�li-�\}���A�jl�i�+�'�Δ�bD;]�� �r�(
ya������R?i<w�L��:>��x�I�����B<����0C��+���*u^��+F���@�DBo��� ���'bp.��b&_�+���V.?�)݆p�#C8����la
5,�����B�5����!��[�m����׋,�1�=�����/�Ww�a:�p7#'��z�ut�'-%���X�.7�ٞ��ߑӌ�ޤ����j�o�!���R �a ��2oԂ|�Եe���0���i7�����韕�m�Z�m �Y����KN�K��`mv "�|�X���6k���/n���ǉn����
@˵�����H�fy�K�gk ����B�s����Q��K�8�dl�XeS=����pD�fF��BpF$��á�搩/p3N�K��g���ۧ��|�ĉ!�cT;`Z�O� o �6�u�8��tʇH�@�o��	�3c0��P�.��̲� (���mlI3'eR6��m!`&��+廏yX)��7��T�A^�W��
|����v�GL�UÇ܉)��k�~@[I�gˋr���g�c�5B�u��K����ޥT�l�چnM��a���4�<?�C�u�ɥ���z��df���D0y���0g��B�+�ӡ-AӕUƭ�)M�Ð�+�m��X�!�<s��]"��, κה;B o�R���v^�׾8L��,�.�,_��Ac˸�ySÌs��s�T��6{�n8�6��M��`B�Dp�+r���'O�	Q����oˑh��I��*�a�{�a֭��Ŋ?��.���e��g���Q���0�E�0{���ʤ�eگ�s,�������,G�Ԕ>W8���d�	mv+9�@�__�u��.��#��I{Ӆ��;�
�R�qwn��p2��tf5�$�Sm����J?�eYd�ۧ��-�h�KUS6֦�ɒ�)c����V��ߨ��Ԧ��H�M�E.b�#���;n�mv�nl|L��#�x��߈{���d���KSэ\�*��<�:wW�򿖩���hpA���Ob+Ό9��x��[)y�j��p��&��(!�_���&�G/P��"���5d�E�"+K�`G�ۑfx��FQ"�[����%���Ie]���$D{�6��|�Q�����uؑ7�[B�E�0�n}�_!le�]x�4��+����BONу8^�ϩ��L\f��k�9wá��h�#j�L�3�$�> QAޤD�,NH�+{=&Z���մI�;caC�O��Yr;�y}e���Lܪe)(sY6#��p�Ի#�Nh��kF,n�i\S4ro��#�l��Uf.�H��Kw��z���Q�
�E�&+�-ӽLMŉA������^Xp�;��� � f$�~��)�83��v�đ�(��P����xz��{�C �)�T혅�{m�@9jJ�죜'<sM��b�(��lz�LO����?g��������x��ᱱ%�*���$�A'��b¨����G_SR���[
���@�N�|7oя���Gǯ^7uB��(��c���eu��)�\U�-�3xۏI��U���f�hcMr��Cf'J�~��H;P��M�I�S�\a�+e�Ghq���"��	�'|;]Ec��)`y��J�_1�s_��K�Q�UJ�w���l��0}���rD$?�v$�U��&�n	�{�{�0�5�@��$��S~�j����pɋg��K���/e4����d�᜜9�.�S��G�W�^�G�o~��?�Q��� ���~0��s�R�NBb~}��X��//��F���.�v��$?o���E;�E�����Y��y����n±[�:]Ы�j9��U��7����O���=Ⱦ���V������:����%�J]U<[���4+�l|���X��@,(�k?]��]�5�G�1�L���˺^U�ewƷ�sr����p��"�bBL��"�C��kkB�~8jN:ĳ87uN���ԅ"�U*̓���]fC�!_��`,������	��7]D�
���)*Uk��s��}����>���KIs�t3H����w�?L�	��A;�I��
��N�8͟N_�k�]U��d�ᥲ��Q0v���������]�V�5%j)�6�0^ 9�x+h�%3hn�c����~�?V��-��GM�i�f.́|�..1ƏJ_�\#i�ut���1X�m�g������)%���?i��g����/��R"�y5Pa���劉R�d�$�Tĉ5��AYM��K܏,�L��6# �l������殜�@���h��o����/�
��6���M��?����!NR��z�f���'�31�����L��96l(�h2U^l���iM�<𢇛�����)m�g`��+
���[b�M]Z�PEM��
�`�	�l�qN�	����+W�%6��䋬�ڳڹ]1�Toj@�T����e��}Q�+� ;�a��O��?�{���W���Pa���un���m�Ư��ݿ��o�}*&G/�CtqHb�(@�k`O�T�t;�]])�	�� ޅ��5�ճ�rR���
,��9U��Due/��uԇ}}g��(��o[Ʊ���vw��>$&>��I/F�%9v��>Mɪ6��O��:�l�Z:�_g��]�΁�1�L#��Jx���0��#����P;C2�iq�6������@�CfNc�Jf�����O^����Lޞ�3ۯ���,��-0Tt���u�?��+�;�J��y[��8ؕ��M�w����K�XAx���7�}�y��T�As�0	dJ�k�$�X��#\�.&*��VE`Bq*+a�qF�?�t�خ�����0Jd�$v���l=��ͩf�g���A�䫫0V0V��"��5��maC�t ;��2a��O�.�Z��n������{�B�A@JQX�W�X�<� �oc�e�o�bq1�b���tZ�f����ř��v0y�:�<��3���_���VH��(����XT�[��Q�.��������r,����|^6}�R� 'J�a}���E��:���y����k)TMgz�E��θCOGh�Eް��Y�{6*�� z�F�@�R���2�	E�ޟ�#f.Z*����<&iv�M".$QYg�FT�jǙ���:��o�/��M�Zލ�����}�.ok�ӯ� �m�p���7�Z'�Ywɹ��y�~��_Hx�m���5ok�M�]�*�VoB��f{�$J���*P�*��6��"lC�E�Ҩ�m�K̜?K���}�ܬgz�R�cb��s_l��-aHq���X���)Dp`��{�ގ�D!
�GTy��k6G�{	�.�x��J�+��-i�Ǘ	�[ry�{()�-Φ�"Kes*���ak_�<l@�!}�$��@�V˵��YҔy<�l��Wt�:�Hx�R(thJLR��(n�s�-f4�8�]�D"�,
�:F����\N0{M�}���r��a:W�ZX���ߜ�
�XYwڣy�V{�ff�\u���¼e�Sպ���>�+��&8`!���Pa��&�I���pqg���C��7��|�W.���k,��f�!����G��'E[3�YF����$z�Uąk�[�8�P��s�?�V	8��5	�{:�E��?q��+kbp�p�'�	d�x��Q�zr}HV��B���JGf�k��NG1�S�K����gSh[d�8\�RZú�l�����~�'�J��5'�K�2K�%��R�i�y �D��_����a�6����Sio`�v�om��k�ag���f�c��˅
7���C��l,�i?�ND.�X���g>���	��c�ǮձF�6#���\ŕ5Id�s�3� �A�o�u��MW���tz޾Cג��v~l̅�X�
$�wL��&�����\:d�T5eW�������6�}[
�S2]&)Miw>�J-FG���J!��M�� v���If%ԓ�Q�%}J������u)?��fo�
l����:B�ILV����A�R��x����v��߫q<�<�ۧ���.,/��+�1� n�T��QYn(_<��P��ad%�ԩ=�&�C��Y���-���c�9w6i͒�#X����*F �C~��8�-k��Z� G�@��z�H��V,2C����$��,^Tǩ��L��O�E��lk�6�M��A�Dhwsa�)bh�j��YX��E�������0�g�:R����]��/XCSƼOYM&8.��3�6Z;e[�����VY��CEs���[|����f+�-��~�f`C����By�~Ԋ�7ۓXAtP*���ս��%�=#4F�u��� _�Bܲ˅�OΊ!F��?c�U̇��Ӆ��C��ʄ5�':�ހe��8_�%��1#b�0���Q�]=� �&2/��.g�G5��r��7&�'k���tߍ�G�����~�g,ɿݪs5��oj���.���:���v~o�sMI��g�5�%�mt������/�Z�i'x�,�"��B��ć��Y�=f?�>$*e�G;�UK,Ҙ#Z�я�6_AHwl�U_�	��	נ�+Io.^����m�K�2!�6�`7�&%��_3�_��k�0���"�&��F�J����l�EJ�&���J�ڼ�SN��/$��������Q�ψQ_�L��WjL5[
�߶S=��O?҂���P�;�/�ϝ�oC�e������[G�n�@K�a�hJmp�z��w>xẉrƮ�cR*���||C꨼'zWf��nﲧ��g-o�[k��=V&V�"�y�Xhn_&��
4zL�	ǘE�[��ԇ���$O=�Yy#����Qm?��	1�%Έt��>�21�l���9��$Lm� d���RǢ��4��~_ u|'��{8�T�d�c~+(�=�(%���d�I1��8�7�8��g���Blߚ��+
����H�T��~��R��V�	�n��c8]�����I���(8*��M�L\m	�C��M��i\���`�}�A^7$��~��?�?�$�����h+BD���H8�v  Z/Uz��+|�V[IF �L&�_,`�X��u����5�(
���	#6v�Bq͝�,U��E����P���k&!D*��)�(���j���+�%��1m6�K/�T'� 2ؑV�+�U��p��y�=NkudP�f5ǌ׈"���m�W��l4���k��&��#M�^�b@�[]�3�^�U$��s�b�^��������{���r�
��*�P�������h��/1�P�ThE|*���u}�
3��*o	-����8��[�Jf����5�?�1WW]��n�Ȼ�4=����2�0��r"��V�����/Ǝ/냱Y��V���_�I���/X��D�,��P� Z���������s̻�����sWt���h��\�����p^<o�\}pJ�%��W1�EcL�w�ɧ�z3g����q������/�*x�������CL�Z���}tcu��F�}{rϟ��@dL�H8x�����|2)�}H���m��T���yB� ���	��.��¢q���^�N�2ߙ���7�b,�C;;���uF���$P��=Ʃ�����`�@���/$�UF���*��S�L7�eǷ��U���W�a��˩�W�I���h\H��le&�=QJ-��կ9���Lbc�����D���X�G�_§Zg��nzoLxeU ���ﵪaϏ���Q������B�]}qXu�]}��E����@��{�U�Xz������Aj�y��F�юf�b�"�?�QG�3��jx����=���g��R��5#�ؠ��+u\�b��\R�r�!7ߣ+9��\A������^�����|�y����3�!%��i�����Y��o�JSph��F$x��F��"~��rBU�N��y��y��^�F��Ӹ��ub��-=�[Vn U��x�ϖa�$�~?!<����FF�p�m[ɕU~>h��∨���F�x)�Oګ�Pǟd��^u�˜�(r��415�c�< BXsz��A����+O�&���ÎNĨ����ey.S��T>�엡�O|~?�S?�i�g2�&e"M2�iy1���O��M�U�%
���t���"�n��e�F ��]�� v���+SُSuG��CC�����C�Ե�	F�݇�Ǫ aOy'l�j������R&�<�G����������9n�������7�"Y�Z%&�#�Pc�����x&֥�-�H�Opԉ�ʫ�q�a�F~s(\�ʶ�fɅ���y�ڴ�y-�-SDҹj��PEk�ͱҩ��K`;��2���P��߶��<j�oe7�Gu��s?b,4K]M�t�hT�m��$4U��Ď_䊭O9Hf>_((
c�M��7�Q���k>����ԝV(�|9k�������K��^�SRi�E���~�[�ge��X֑9t��D"�7�ڙ�cU��uu,�ls !R{~���� /��?0�k�B���d�l?��}g�W�/���w��s�I��VQ���l��|�+��3�'�d�uV]�8��r��e?��۷]�����e�n"5����K� UI��lǒ+YR	K�ݟ�cs�hBj�&���d"�H�4���F)6o�����b&�R갦�#{���n�V�d�+�C��O�MO �H�/�����P��,j����t3"#&a�Je�\X�!:�"9���j�6�5<J�V�����a߼�"q\`[w�����$`n=���i�?���k�_��e`��)Q�����i����d �hP
(ǳ���ܧp#�9рy�di��bI}�t=�D�aXφ�P�[7�m�;�Hގtj#���y���Ь�6�2�M�_���T���i;c�`�j�G��5�����;��+>x~:�θf;��a,06Q	�u`3�3�ؾur@(x����ޠ�}5jT��6���~P� ۧ� �n�h�Y؜q�T\��	���A�R�7�c�!z0���;9V����ꌀS�)��C�03�A^P|�I1��K���d�9	P�E��Ed��6� ���
���茻��V�QZ���k���|�M�>H��:-�(�zU�s7rPgs�Gh��c��s�볈�(){/����X^��2��0��f4g�fˌG��g��P�/�K�����s��LlO�����;�U8	xq�U\U'^gJ&�i݊��9��]�Ya��[z��N]}ޔn%�W�֩�;-<�q�b��@���;���3w��v�*z����'�XO|�i7�y����ˁ��R�~�=(,������΃��C_Ӻ1w��u���[`����AAy����	њЕs��Zoj'�1(�J�6N��4�#)�����'�ɪR��T�Z��nH�*BC7(�_�޽�����Ь�G=�SN�Y�� � Iɀؙ���>����Cv�I�m�}���M�#m�%?���cn芣N�p<���>��&�����zV�G2�i�CHXU�a�ߪ�����$=�5�?��J�(	�P4cH8~9$0\q�j�=8P�_L��奈Zl��pX]ݷ�Q�uL�ٽx�'���ϖ��+� ���H�q� �>t$���y*��\��t�,*X-���L��B=D�9��!�x���IM��t'���F�&�s3i�XA[Q���*z_��͊�a71Q�G�P��R��1?ɵSl➐�֬wk��r1:�)�.ˁx�M�,�k;���6N�n/v�h�!-<�y:�	 �!¡�}������s��4���?ݠ��h���MZ��X�D*��(ḁ�D�@\��Y}ba�U�|�i(��}� T3�}��ijb��2�_��y� ���O��8N�:��j����*}�U�''�����~j9��.,�55⬔.C��T/��L�֙�n�<�.e#a6ř%v����9*���̴.�����A�p6Ԑ��x�m����g4mH-��#WPsr�@��De�~�j�c�EM�Y��mkLJT�q^	x���»�ƶʻO�0qo��'��I|�D��׬�^�ӷ��|��*�rO���@��.�{b�h{cl��g���e@"��>��.��n�+��Y�����j�Ր���Y�[��rK_�n���m.Q�~Z�7.֔��ʵ�o�Mjᾁ'�+���
B;�����ը�?�N���[�_bKe1z� �}�������z��	J�+g��������&I�5c۬ �F���pO+9�����Ϟ&�28�}����(s���V��*ҋ��]��QOi�\Q�� ���Q�/��jQ3�=0�E�m�p�1ѕ
�J�p��u�'�24h������cI�}�8���ɱ&�n�b/�o�Î�� �}���Ĵ|�1Y�%1�՜�H��o]�� M@��>[�eD<!-��JHt�T�����^�JZ���g�΢���3������r��$"nuP����O>����q53�&�&�˚a�~Z��<�q�>V��n�ye��ι�uoG���e�D��/Z��C�ѥMt3aI̼�BZ-�.Z����*�g�[��Y�8pv�]�W�3Y5R�m�@]���l5�ɇ��$X��y���a��3@�	s8i`9����ԍ/X!���B�>T-��m7߹��eU�i���Y��2*t��OP,��2s.�#�&6�Fn]\����C'F������s��xg�5���V~��?���!
L���}�B�L��MP�	&ag�L<����t"Q��X��d�re�ylU%>0׮��#`�>��f�P�B-fpz*/�[�h�.�2�(�B*.���HA|f+I�`,Ks��wP���|�H��k�`1jGڽ�2-bS�6����r��K;%����g_�隮���U�=;�+��6��&�,#�y���wC>w��SH�O�Z����x	e�����#�`�͕�h�Qt����S�ơ��{��*��P�+Y|0�Z�ͫW-��-��1����#���&	zh��=꘱V�'$_�d�{	��Q-.!OBr���s�d톞�r g#E����=y,���)����?,�S�Kf�$7v���7�ʗ��������;��:�|/7�m���.�Ӂ���&\�?v�]� ���
䭆(�G X���W���җ���]b��f�
qը��,��_���]�u�F(^���_�C��H܊��cs	����u�g�O��ܑm�y3��{��Cŉ�#�E�Ý	��ө{z�8��e-\�l7yv�ԕ����J���X�qG\$Joo��*��bET��I�� �5(<��)�8�2*���Mg�c��zQ�ԇ�@��\@�s�	���t�@=��	BЯH|�V���?[83��q/�]V�#~����
�����d��7٢/LiPB[Q���EQ��{�H�u�����c![�+#c��I��'�goc��sȩ�c���?7�Rx�H0J=���L)d�Y/+F���i��s����������u���¥�*/�;���V�ΞP�C�/?|>�s�L��:R��.�0����r�0��� ��z�Q}a׽����ͥ'o<�ߝ��V��ecW��Um���ͼ�B�v4f�ưz=��$�'t����c:I<,�UVˋJ���3aV���Qvgq(m�
�����h+����0�ܟ]Ǳ�8Q�F�dу�2|�?���Y����Wئ0��!tͫ���U¨^V�k�Zz�	�lXnß����#9��+'Q<�`oo��`9�]���_pK���5�Ã��f�(νj'��}��9��A%���u�{��_i%�6ޫh=�|F��qI��Ƨ� ���v���Yރ���Ya�Gj��J�iL������b�0�,-<k�*��4�ǓQ��7�꼣1R��x�ؙ�=�Q@E�XP{aWR Z�㴯\[�@�a�͝�?{i�'a:r����<�����v�	0�ӷα�ַyҨ���A|�[��;k�7��i�6�W9c
�?��򸺾�e?��������ΫR��w� ~�
���'c�,�G�	���Z@����_d���u򍍓j���)��Ҫ��T?%o�[i�XW3��ͦG�B�K�B�Nɓ4&��Y�����:��r��_O�r�ΟT�{Hp���r�1�γ A`V�<��F�k�6����.��l���}\o�/�}Y$6��{|ǣ�I��EԤ�J�t@�4��"VHh�3�3,�ǲ�~�/��ˆӴ�*�k�b|�է�_�	�N��rV�-��)F��?�z���E�^ j b��Ce��,�8�H��K�����'��GI\@�����f��և���W[��[=���w�D&^���ٵx���9Lk'`ҪT�7�^�c������B���^-L�z���������'6}I�Q��F��k�"�=��%�h��܁�P�,��6�3��nj����]���U��`�IY�{��0㮣� �]��DC~L�^e��d#�bP�l^�*��,��p�߇ҕ��` ��V]哌����7=���p��v"&��c/����#6��MQT�+� 07���R�ya]r��9�>��r�n��φ�J԰T���ɋ�>}�����I����r���ȋt&G�?�����^A{؂N�:������2)
y�F�q��c< ۠������&x�P&�|�}�|־���	��G"ĝ��/%�9�bx������,G2��T02��S�Q�s���:�J0R~����dL���D&*h�o��N����yiY,x��׊��>�b�Z�I8����-�$(f�8�j��}�T��+@�P��*���� ��j�߹E�@ȅ��7�Xv>R�T�J��?����2���*����`G�>߻�2ת!�m�/���0^��U�D*5#�l"v^@X�ڵkN ��@yT~��TS#�����x��v2��_�7i�%�0��x�2Vٜ��B�{X\�m����݂��w"=(�X���؅S���U`+�����;���Ыo;0��������BY��Ll�3 ����O/��\P�bF)����$fY#�г�iS7nÙ�����o]
����g6n��0Do���
V*�h�)�9��sG�tj���}G�nI�M�T�G��t(�^�u�)�O!�$���@m��=n�[sR2Ogr`D�G���4����qx����bh�#r���זÒ����BJd�\P������rL1Ml0è�eL�]f����)�9o>����*��O�$ 7,�����2Q��ح��4�����1uI�Z����4MŲ�θQV���?
29���#}�4�ܗ���,�}M���0Y�=?��Xe�	i���7N"tE�3��<.��׹��-B*��p�t�S��:�E�@坘� I��������G�C�)�{�(P���:v'��{�� �d��TT��~,4.�dϦ��ԣ�eTz7L�1l-l~�W�����8��2Fe�L��@[2ӱ8�p�>AZ�N���>I��+_�{]�0`�CqQ�K}W9�L{�}ޤ/��a��e�A݄!�~�:W{�,�����=������1s?��_x��f��|�\(>{��T�ؒo��s��I1�˩D��\�%��>�{��h�?�<�Æ&-�����`A�)�=�VB��S[��W��s�(tL�3o���#�����X��O鏨Ӵ���)�h1֋Ɩ�N�k��a���z
|{p���R�_��9��f��	W�|}2�8��74ճ�g�: <ذ����g_r�m���2䱤qw: Z�2jg���X��#��9�p��Ys�B���m���aʩ�B�ٙ8G�]p+�Z�ٲxU�ΰ�B��w�D-;��Y8+2�����U :J�������5�u�{lar�ġ�t{ޮ�jƄ�y�2!��C�G��NB�@���`۹H34��d���њ��qdF�4a��SqT�ږ)T��n��Y�#�~�4å0���%��>K����ز�zTGU����{���(�4s���XdQ-�h��t^�m}+��5���s@[!�"�DH@� w	$
w�QP)�ў�->�Ա�c]�(�5����ҝ7�|���ӂ��֎���G�$6�|�T����`Nx�B� -��F�������Z��.�F[C�;�Mf�M����%Oha}�９4a��x��������fy�G�J���B�։A��f1S��"g��2����_�����m�@��^ej-�7ڨ�0w�8LG aC��&sc}$w�����k����,[��a�L�V<�&�dФ��꘠��X&��`�'���[A��c�
��{G��5&Դ�^�0�*�V�y-���}o��.�piioX�Q�?��O����_�bAt8e�u3"<|_c,�%�9'�73M�:ղmu��<�j�NY��C���lsC:��/G�b�׫q��\�n�EdA�4�c�� <EA�� Q�N�����>��e'�C�$�@����m�ǚJ�5�w��4z�B�_K���ұx�����ſ���F,�|�/5��HImS����	.xw� v$�[!HKX���R�ɢ~���+����PR" ?.���3QF��S~	�~9w�m0o	b{�nu��k��X-�(��b��I�κۑ�1�L��j�V�i�����n���)p����$��XsQfP�u&� ���|�D��򼧽R�X%2bz�\`��!pX9]���҇�f��C��HqY}l��.H����D?�շ�c��$�m��PLWA|>M�Z�����34*�ڭ�UW薑�v�Ҁ�	���HS��KW��wQ�1���=�ڛ�٬T#�
�n_��`7y���e?�Y:r����r�r�~��gU�C�J��+)L��\ŉ���cƊ�R���m����偬ɼg�H�iCL�Jȿę->Kw�
\���-@�,3���j��z)X������fK���7�2����rjG*��8.�_�KT[3�)�;D�P��|J��_��f�r����Z�����N��z�� �زtrUf�RpQ����SuS2̪�9�����q���/�*�Z0���y�Mh�W��3�?ה5���5���s�钓}�H�����Fa@Bߴ2�q��>Gd"��WGc�gx+@����;�-���(�>J�.g���B�6��� 8Y�<z��~���d�~��wۈ4��*�c�9u�8
�K��� zBt�J��`��p���8�/y�+��L�2ݪ6:����)���ܒ�G[�ċJ�����a:ܦS��!��XKG��=1�ȂY��u#G��v��!�H�x�0���J��y� �[�����Z��>��$B�n7;�b����4��ɶ��`��B�)�`��5�����#���1�Z҇̌��7a�J�[�M	OC�+]ȋ��M� �t���.?F�H727^Ԅф����2c>;�t���X<,��32~��U*�$W�c��n3��	�aHC?�_D�������~]�ü�@��&̷�����W���BDR��_�B�N��.�	r8�P����O}���ȺO������f9 �]��=��������w.�_k�~5����
���
t�W�� ����c��@]�D�܁�?������ֵ�/����V�z�,��X4F`$��5N�ә0��htK�c�ٙ�6��R�pӟr��"L��� �{Fa,h�䆐	���8F�R7�;�+W�Cu�B�ڿ3J�(i�7"�a���Jl���_:>p����預���.|kCs��������'�-�r�]ۯ�:o�y�����浍��&h!zo��K���/��鰥fƌ��qʹ]QL6ǃ�g�ۑ)��>��Ǣ�q^*Z�A\�iq��ⵟ@�1�1!����r�e�_><|�#����ϺSq��Y�E���Z/����2?�:�'�����H��*�pGE�K6�ӻ�湙�W!$���Oc%)&'��p��x]����u��H{����?����'��Oh���Ѭ���|�'��C��!֗|��*�J��Z��02�ػM�yo��WQ��΅�J"����<@dH�4'��ۨ�^?&�58�T�r�ƣ^z�.�l��dd����Շ�d FO	�k�m��~yr�yWX-PQ���Ͽ96�:} ���D�~M�ZG��_#����թZROӔ/���$N2������
5�/%��R#��w��	��(�ݐ<0�A�k��3��ô��'�A���1�H!����%ZN�ǫD�l�����1����p���ˋ&d�E��ǧޛ�7�Ըd蚡�.Z�j�u�D����G�����"y���RU�I}�����3�I�Gx��ElO;���*}��p��x�Z�E��)�,�:��,�f�{����=#K��rt���2O� o����ƬL�P$��\ j����48�N���H ��ǁ�.��0Md�O/F���.�"�vf��$���V�=)z�v�&&p]=�*@1�P2jv
�\\y:�	*���\b/��� �{�IW���A���QzL���U����\L/PәJtV��q�
n�ǧ5��][�cI�S�\ę�+C��r�g�z�O})�-(?ɣ�?R<��K�d��_�#���i�aԖ���>Y|��.���'��N���W��TA�JLu[z>��n��yx�A�®w|n#���r_�m3�G�e}�N����_�YIp��(��6�S+6Z�ū�%�*c�<_Z���֧1�&C��?�<I|�z(��^1+R��٫�w�7=衏�@��9Nr��=��/�B݄�S	[�d�ٍ8��8�F���LWKa£��z_�[�'ݳF�<�jM����������0ȷMb7�0�#�y�D���]��-x�[�ݾ��H��;Q�����a�h�G�Kb�W��^'8�G�Ρ�|�6�YjpK�\�l��ߑ{�F e&Ӣ:�7t��7��%A>w0A����x��6�1����1�]���'�O
Z-�GE`�p]������z�����\�bϓ7���f�Yiw���i��o���O�"�i������������4	�NF3�Q���Ly���o��gc�#%[���;[����|Q���Ep�Jٟ�c��$7P��F���*^i�e����E���F���u ���i+��c�����dJ�&ě�_�l��J��Z�NƦ���\uTJ Jju�I5�?u1��ٚ<0L����>h3�)��B�\���U7��������1sn?���1q��O�g��Y�o�@��W#��㶑U�ͷ_%�%��0)lDS�$4f��r.Qm��e!l�K��
�����Q�'��C�M���&,p���qK�C�k~����5�~�<��q�c�tdޱoO����Z+�p���_#=�U��ګ�>�2�J����@JJE�>��-8ݬ����?720���)u�}$&��x;��BS��O�;Z5����L�,�_�,��$(.�򍕡�=�E�2��u
mx��Vlﮠ�*�6X)���{D8�ʚ�ME����E�tW��yq��	v%�v�uR��'��P���G�3�KDGzANNt�׆��!袢vB�`�(�%#�rT)��^�	z��i\�3�^2�N@�����3�6uGq pŃ&d�ih�k)U�ws[�������k	Ɖ�-��4�Um{7��߱�|�p����p]�:��A���4R��#���j��#>�ڷ��Ii����z��4"cJ� ���{LAda[������!���-a*�Wi&�k&?�&�YV����M�N��f,Шd����58�D5��4����]K;}��v��߳�b4���[�Є.-
>j�uQ�@.�X��`~Zd����@	�����h,DhN&D�@�9���=�|���Os)С_T�ϣ+��T}�dJ�bCmMm�z{h4��x- w�M�0��J�)ء��L�֩����B�����fQ�d��N��n���J� *x?b���������l����?�F�, N�τ���{�� �I��⸤n���MgnM����։Ɠr���e �XO�0q��'����������:]/����}i�\*c�SP��A�W��X�.�[��m��и�D�B�H�q]9�/���t������)<�?��'��Ob���.P����<�o�����آ�^,z���%��9�_�1��p8ԯ,M�R�
���3�⥦'�9���+w��~t3��� �rv�Imh��,�`����c�|M�S��/&�{�P^�}�C}�)��ͷ�����G����/�S%K�����L*T{�F�Y�ۛ-���M�?�����U%0�I�Ҳ����f�����KGQy%��e�5��Z�3��]LP�ջ=TAY̛)uGͥ�/�]��Zt�B
1Š3���J^;�,���!Ue�avֱ<��_u�X���������)4�ϥ��6��92%����Gp�X<P�4OwH#"��i�3�ǛJԬ�n9�*fm�ێ�|��Us�rI�k\?ԡ�O���WԽ���@˼��@��k��5����Ҵ�`�]���Kc?�����9�= �{��ן�b)�O�OҴ#F����䂰�A�Gϊ��b�f�3�ۼ~���OЙ�:Av<@ox�^hcRIpWfNk�6��&�z陏/h5�4��,���G֐��l���(Ғ}��'eA���.g�&��?lm4�w3�
�H��~��yȏ'�/�?R��~s�粂W�'�!�S%,�z7:����j ��w�Q��lg��#�g�p�� Ԁ����]�j�e��6/Ya�"�s�ך}��}�o�7��G&��v�O5,Hʳ�F\�L�Xk���x5��9Km �Xs�q�����~:�UǱ��n���>0�ǲ������'��.�WK�"�䖤����tRͻ�e^��t�������N`>c�6�D����`3�q�-�!��~���^(-�n����<q�[�Z���:"`H�QV���>0���l菜$���7K��T_	[~k�*�VV����G�X�\t�*�\/>��[��p��|�Z�ܸ��=6B���rˏ�~�o����b�bn�ʦ�}���o�L�׹@M�@�/�
f%3��t��Ȑ�kd���*[* G�{*g��ّ�Sd�ԗ6�֡7��3=���BpeGێU����⚗�������	ޜa���yT�8�J�כd�	�C�����@���}oݔ�.�܌�^����MT;�ǉ4�ÓuUә��c:Z�n��1����t��q�p΀��5r���U,�g�ۙ�MHM:ԙ���y��9h�-FU����	���D��^@]�T)J�;/���t咣���bM��:q��C=���Љ����F1�VP6��wV�����Lr]�X�gE��8�q ���c�������|�,��d�^�p�ˣ�ԃ��|�ΨkU��/)&�����3p�~x�_��</0p�㏡R�JY�&�餺yX�D�W,�b�/�Gi���`y�<E��QK	<-"3�� �_\��@�3�J=�Ue{*������C)� ��������q),@I�f0w&I7(�Gݵ!��gғ������/P>O| �%�9�ͯ='��ݸ�U1�s�
�L!�)����<x0�w	P�
������j���[2��e�RK��v��v)�ܣ�X25�[z��2B	�%��M1�υBZ�U��]ٵv���֙�Yf���h�'zF]	�m58�˹x�3EfӜ���}Bb/�㏁��ad�:�4|>M1=z�<������Q΋��_S�L핌���rDB���d\\)C�W�1i�͍�_��#;SDM���V�H)j����S�qx/K-������.6�� ܑ#��cx�;	I��P%�� ���2N���3_J@���o8�yC�)1�\�V1��[�'�k69J%N�	����z1�]
���9^����'g�&r+��ᩏ�u �1�LҦq�*�~U5&C����YT�t�����0�l�9�Ʌ�0��rY����s�lI{��;_w�%���	~i��?ҍ!�w�k9����S2F9c(sY�zS��S��!��j�f]hʗ�-�񹱷'�{U�ٚ���0%���	�̖�l#��pQ� i~k���*�DI���@����λa��o���!*�S�h��Ձ㽤i�v����r_�C�+��@|��2������!��*"�jҘ��\JZ���bMR�
h���#�͏y���D���_���4����R��k�0_�6�K��SE�-�,e|1��3����0
��䦛�Y[C$h��y�7k���?�gQ������E	[��{Ѕ��c����Z2J8Dw�x�{�����_�����zD�u�;R�k9�1�I0�u舃=Y~VFI��.R:+W�ԅ�,��Yr��[!2��	:�WF�5d��9s�UIOHJ�َ��z������tP�K���|��c�V��>�z�����HyN'/�l���7V�;ӧ�a<��-��J���-�"�є���W�9 �v�Zf�qF�r�C�� �����Ç�"V�W[����X����K�ߚx6��T�h�|c���q�c�"�! e��k6��BB��7�[h��ӳ���+W���Qٶq)��u!q�h�v�.5,)=����$T�!d%*�=��m/U<�&��7┮�c�t��_�"˾5V�����2�H&�R��j"@D�4���m�k9a�V���d�O�]��Z��v	}])x�ڏ��l��[��=��h���A��U���o<W���C��(�Q~Xs\��_�!�8H���tk�6��@z��l˞�KI:{v3�ޤ^� ��Y����i<y�Su@�~��[�і�R=��6v�H_��vJ����0<̵��A�VU�8���VN��}�X����+2T�h_�$�V��Kf�U�_�m�Ds.;�*r��i��pTF�={���QF8xxy����Cg%y�Vؠ1ZL����0���ib���@e���1zG�I�2Gݍ�Z0юیXC��.V�i��6�BrP����M:��~���Emҭ�@��3��)�
���H��ܖl���!.���gf��'��ݴ�D
[���#R�!Y��֞@8R�5_C��*<0�K\'�WȲ􎢄��^�c�7�:L�./d�羍��92p��
�짔����ֺ*Wz�L�l�,q�Y����![$9A�jp��ޑ�M���;�d�K�A��-ږ��#\��؀�� �tTƤ�7��=��T��.��X�fC(�ץO��_�j9Y �]V5'���r�E��˅#P������Y�/�������z,�AQ�q��ÚV(�Uq5���-&�Ϋ���s�����9F��;'f�|{��XD���,žt�~N���h�g.Ǥ�PM$'>[b��a�,H�~�W5^
E��Kh���>�����³DnD9+Dd��l@�l�b����_��1v�)I���/a���*�a���I�.����(�Q0��Z�E���Á���˨N_;��mF�h4d���[,�ZE��I��j�O�`Ox�Eآ�9�&o�������A햧_�`P�8��@HK1�*@�{H	2R]�^S2��hR!�i@�${���5��w�*�[� �cK�aC�8�����zv)�u�%���	����wuٸ����.�������Չ�y��
�!�|/*H�1��wz*H�'Ւ#aW'I��Ѱ�u�YxW<	�t4'���CS}B�M�L��M��g$�����M���R��O�<N�UQC@��)O�(��zW�e��Py2�8,�����x�;)-/�0k�4��F1`���_tm6i���^�l5�L�|@w�-����K��ZL񜄶��l��������L�rυ*�p\�`�7)�5!��1`��\Ͷ���G+%���ͮ�?'��W`%�WhpL"��9�z,
�U�J����$dwz�	|�����F�^Yw���r���^x�
׳��	�	����D�Y�������$����t1@$~�*�l�Ap�p��6y�^��>����q���p�N%��rw�,�A�s�m,��EKLЮLl6��"��i���2D�� P�N������6Y1>C����6Va��x@�l��$���*E�!TցN�q!�B�i������>�^Ѭ�g�A��T���E�C5�
o�)Y�+��64ɢq�QWh6�$��X�^F1�+#�r��:/V��鏸_����"�1Ť�V��;�^ʯT���YA=�[���M�{,��z!�2MC�E�	8���ԅe�}���I�u2�l�b�,������w߇5Y�{\��Uu�� �UMV��b'�5�*8^�pu�z���,�l�IzE���`�u]!����z乥�1�G�{�ֽ��ɋQ�0ɦ��#�Գm ��Č��V��*�@O���}�y��Yű0�k���K�f}����L�o�bŸ:���Y[�Z$̞)O4��/�^I��R@L�v����`)�e����	#Kbo�+h��x���>.�m��wR��/pn�� I� ,�#��Ƶ�	����栉;}��&DP��,�����7��>}�G�����xY�?2:�|��%"��%BD̗�L��Vj�r'�`��0��+�6���ʸ���&���/1oi'���,� 8v��e�.*�xX*�4u��!]o�&SL����8���꣎�~��Ġ�Evs#>`K��	JI5��w6&���Yߠ�]1g'��у�����`8ֵ�!I�����]@K${T��xٯC�ΐ20�s|�½�_�I?HB���f%O���/\�E3()E 82�
���a���Kcr�o4-�]�:����1E0�+��gޏ�H��T�f���������A��,D�Bώv����% �V��0s�l�O|R���	��ǒ/�j�p�u+�����1@�Ҍwe�<\3`�ˇ�{�I."��Z�N"�GI��ܡ?R�����ԏa'�`g��}*��<�ƺ�K ՠ�j�+EP� �R]�6�?T�<$Dt�t[�DtK��Y�SM���$-����ҹYo�r����-ڎ��+���B����_�JP��'3U�j�R&����h)����'oy�����AyI"��iǳ<�>�J��SmH@"��_�κiQ���k��������hD��'X|.b�y��r�9��d �6�=�=����kKM�23�M�����/{�[�d��Ö��x�Nu��&J�j*#%�H6����AXw\L�~�*q�U��\��ӽ<օՊԺ�(�(�q�:%��7׋���}��8+�b�� ��6�dx�O��f.�
�*NP�4-�U ���A���1�t�$�vV���v��PA��e��[,+�DX�����)ClJ}�%`BX��oꬵ�'��|���n�悦"��9��@�˫ܳt��G�g��};�Oo� 5���JYǈy�I ��Bk8��9��["n�E<W���2�R�o@��u������_;����z�h������W�hm
�$�ٔ�jS{�S�7a�g�S)�:��w*��aV���I�jI�!�T&k�O�^���+�+�}�k���[�{�����s�֗���y� *��~�sޕƦ`/�,%�$�@P�Q�&v����oVΎX���j@"���2ܲ�Lw�1RI����zy�ơK}��	�a<J�y��� �Z�v��U\K�&^=:	ϥ��lq�_3��2�H�[%D�$�0�+�����`I!P/�T1�i:�7��rj?�Բa/v���)�5�s�b��B��þQ�	� ���!�c�I�+�y��*���G��C{�.��o�t��i�6�wXQp�6��㶅<k�e*l�Yh?!�8q@D�U�u��37�s��k���Ik3��lc� "�򞒕�|��}cA�����`yH�7����u�%~-��"��g�t��.R�Ø�7�x�&�xǖ]:J����e���e&��h��z��w��晢��AMU6dsMYBP�}3�k!�â�����G}tQ��	C���$;�WD�6�ҭ���e�����ߜ���{�TQsY�#!�A�8%�v�i��>��X���2 ����l��~���#U�&�,��:I\y�dgU�K�����v=m�n����!����W��?�:��>�=�d
��q���̐�V�*�|-�E�ڂ�	��ĸ`������	Ӏ���1��b�sۀ���~���F��G�������x�1%���9�nm�D�\�ܮ��7�q �O��+Z=��N�~ﴎ��{cC_zFKI����%J��wl~���7d�Q�m7�;1�{gW�ĭ΄"�)[��M��4�+�3���}r� Y6	U�KH%䰹w%&>ӂ_�gޞm�U�>g;Be7"�`e�-��ӱ�n|��r;����%��/�����M�$���|�L�������da���R�y�sΥ5������o�~!�)��Z�6.3c�N��ǰ�*��.��
@�8��C����s�qG�̟�>��|��Κ=A؛f�<����+4Fh���;
����u���u��!^�Ax8�����ǻ�����|_7���T]0	;��Wz�42:��Z��.����u�ީ_*Ƽ%��#
=�����Ɖ�
&l�^"�{�5F�(��U�1=�U+�q4E~��|����8�kuK|�|�
�>�Z����#V=0G�pEu��@Jk
����S���s��~®�Q�*���7D��_瘿\��ӣ� ǦɎ(*��{b�$�yl�q���� 9�̎��_|�����.;9f�jg����+0��s�Jj?���(�*�ĔM	�:��Gqe>@�k�m�KDmͷx���J��uH<e��V;c����������� n�Z��?��܋(4h4��o��F�/
�ޑ���'wW_H�f�_�s� �KT���X�i�f@��s����p��"$LirPV*�MDLnu}���U��λ2��>��-Y��,r�O5��f�/�p�3�s�Ӹ"�3�gO}���Tu�i$0P&3:���N?Y��s��p��8�V3�DFC*��MmU.~��+3� �K24vTs��Ǚ1���^�R�Kvj%iu[��\���SC���G�__�(�i�1��g`K-��ڿF�Ӓ�	!��-aK��,�V���wrmhג��S�~i'��%4q9%~3d�#�6Z����fƘ%Ǧ#f��{��ɗk�	|ǥ"i�4^eV�K��������� ���&��K��r	K	(�� �e���7쑣~/[%!�@��2˩��έ�zҗ������QJ*��d���J
�&3��4������eĆ]R5��0iT��|��N�[����[�!/��;/t,S�"���R�X�}���3�g��?�L�R��n�x�Z嬜~7WM��b��id��/��L�i?|W|ѐ��ɡ�	 
0km��b�"~�ּ@�,��H�f��M&�m������hjQ1C�H5C冓J1S����w�� �=�C�p���@I
�*U�V�@1z�FUk��(RmE06؃���47�p�u��u"w�ڡ&R̍�H��ƚ9/]lPP��HUj��.X�v7��>c�ܚ��-?*���D�}����m3L�Teƍ������q]�~������Nգ:Ȃ�#��܅cj���z��:� �[R� Z(�_%�zn.w������6�fG���,�R���5���/�Ey4�!�5I�������`Պ&zRz#®��5s<0���H�vN��E�	ij#���=�N�z��R�%����V
M+�y'�LRW�d���ݯGa�9|<EB� �Ƨ�x� O1�X�T���������@qK'\}SV?��]�I#]�-9B��P �S��sYá!��J�t���˫��0�A�_mOt.>����-�� �E�p�Q�0������d�����1w�7�Rn�Yx=_>G�i��h�}L��@<<*������ww���>_���E��)�{�}��H�1�A� dhI�T�d�h-�Mz��WИ74
aע�&Q�2	
��C�;A�Vj3�n��=(e��؈�]�ks�䖊r����IG��we2�I@��e'i�LPbN�B	sb��0_������~*�r�E�����gA�%{��,�^$ -�_ -�Xh�(�w̟z�z��E�����������X�et�����b��гr�i���6������.���l��kI������^$LsE� s�nu��Jz�s�q�9��g"Qr�W�Ӽ��.�4_�;^(5X�n�n#���U��a۾i�r1S���~���K�-w!�nONY�~��(Y�B�4x����C�
�P�U�4@��4��#��GZ�E�*�z�P��'2�a2��r)J�}\a��٧����,S�fm?Cc�f��|�~��`�	���rXY���
����6A��P���0 ��i��~,���0�3y�T(:Fd+�Ȼ���sof��k�cH���b��P!�{HC�_إ:f��͔�}����z�vgN�u�0lF���k�>]�U�ܽ}t�W;F�ʅk�"e�� R����Y$7�l�����ƞ��^���zv�~�)֐�_	~���E�mʓ9�]�	�i�P�� ��bH�����R��K�sxYؚ��6K֔�6�vf�Q��%p�`̦yp/���OF,�W��ԇm�se]Yy��+�rc�m���(��GbS�N�>4q�d+ֆWt����7�%�-fEǚ��
�Er�K&H�[ԫ�{eP�v��1Z�S��rh�O�t�:^^��O�j�].�i�oA�JȆG���'aq���[Dx;�[�+�
�����A	���;�/8Wz������i[ƣ�!#<���/��ş
2���h��حM~?�d� ���Ui>m�H���Z"��L�T��S-�=�&��c/��l�wvɰ�Z��o��'S
f	�� �;؅���.����g�y_�M���}pZH�ޓWd�Xl�D.��(��<��m���|0Z��?n�4#�).dM���n���n;͕�$ح�iQ�;ǰ�]�B�ٙ'{�˼�2Wǳ
���������������V3N�ݛ�p힢f5y�����P��/-w��ψ�0i�)]~o�ڇ��R�w�����o���p"���U��p�[,a�y~﵄j�yC��'�w�\i'���*�"b!^أ�����XY(��%���A��%�+�	}�81`g�̫\���$̶1����_�v��e���'���Ѫ 8w����nq~)���]Q��S�e����K�0�:���EP<=�j&!�d�ڰ�/�5��j#ᾛ&)��!9O4������D�m�8�|� S����{���p�Y4~6m���@c!��F�Z�{���Qݸ�U�-�����n��
ޏ�a�q�#{ق����Х��hk���\:�N��V�ޮ&6��/ay���R����j�L�~��/�Wt(ܚ���|LJD�EL�z�*�Ä0H��@4���l�e��X���=Y�#��P�.W��bNw�����.Y�\?|��U-�\Hca�V׮�*톯.�l��e̐WNV�e�п��G�e�;��Ik@�����U��}^���s�oզ,"mT����m��3���hn:��Рv48�2�Z�w�}�j�ۗ�I�M��jY�p#ʢ��>�:ǟ��S�f�]� �i��rME;	�<��ǵ6_gP���S!w�e��0)$D+��|��T��B=�+hHK=z�LĸRg.+4w2:%�#�>�S��]�<y���Ŏ+��b���ȷ뤈I��1��L
^�� �~�+�i����7@iH�7�$D�b�$� �����6|���H�*J����b�K!���4�]�
���IEez��Ba����hHq'elb�r�(��au!�Ck�����kO�Sl]�e��������uQ�I�=?9�/��:�KI*��N��$y��.	�|s�>�Q1^����#ϩ��j�k�24p�?�D߸�V$�qC�z��A��Fvw�۩�A�/S���.o	����JF��l�.��F�u�T{vLC*��������d��~�<N�G_Z�ݱ]���tg�oD�n$t# ���可Ŕ;�� .&�"�+��cguff"mw�+���U�EA�����#��ޯ�,_aO����M�X!���"���}32G�V&(?��'q�M��{�����Uo`pF����h7����1k.m��#1�j^���m=d9�6X!yT�����
 gb"�㐓{�Rµ�RJ���7�OͶ�{\{�x�G�2$���$�������z��?cIvY�h-3��Qj��g}���]�i��1y��T��:�|x����H�u̵�/[/?y3#.��ͳ3�Z���3G��s��"MJx�����1���*lR��}��ܴ�!nva�8�g
%>�^8�3�0�ْ��1�Ǜ���j���'�$��s�A >�CD�/�|��_��0Q��e��:��L��x֚=}=��VL���0Д��M��uJv	�U~�	?����gM��u�x+���/s�^����h�z��w�>�� �/3�AgA�'��a�{�:`dc9c�Q��?f�]�G�U�a�"�-�kyK�R��O�����5j��wm~�u����c��h���^����bv<C �#h�R�C��=|~8�됀J����P/C]��t�����[��ڜ܋��<���/k�q�\��p�V��=�yG�n��E�R�IwΡ}{3u�iHH���p��$�y�38��WQ^����~�����q�H7̷���P�	o�g8n��ߦ����%�P��G[�*ӹ�����[QLԋ�~��E*j ��r�x�$�j`�����O�>u��ZbKV��������ھ�A'��\�o���&��� �?���'!p��=�U��4���M�%��[Ú�i�i..�|�)~+�re��U(��5����Fm�I��\50��ksk���BU�Fb.p� �4��ZT�
�x��Wς��d�~�Ej볡��]�,��t^ψ����/��:�K�g����9�O�upЉg�
.� 1L�S�t��9��R���/�P��7�?Z�0���M�l��X4(����v"�C���~�(�U��e��0�K���(E3hjT�E� ���dP�?7�֔h�X��ܭ��S��v�;7/�*��o<��{p?�&�1�e���D4�q�e��{v��Zse��Fd,��l	�XL�4�>�3b���fْw�e�8�G�\�=i�J�H ���c��>�?�a;���w�i�������.������ � �%|ʖD�����>��Mb2Be��C�n�0��J�3��Q�v�����+�Sԥa��	!v��_��ngҞ���r!>�JSH.n�ZB]	��!�.��4z�c�k)�f���W�r�CW�c�)Z��dh&��o�G��S�:�Q���6�5�{ڑ�!Z��oa��S�얂vı+4	�n���[s��0��P��f�}=�=�Q��
8Q�T�L�M�S�M3ZM�Ǵ�\[\�xe�֓�����o����o�#�)�&����a�v`lI�ƃ ��-势&��A��Xs�A|�����6D��>����F�s�iG�R'��uQ y)��c�="zC����Ҡ�b+�LBod�����e��zY�{��.� *�z�bM&�}T(����!�dڣ0��|��tH"�w�~��j��k�b��s�S��%˾˕��!X��Yl+�:dM��;�#vr�PdΖ|�i���ށ�y���t<�ۊfn眪~[ �P����J�W��`��u-�D9��$Ϻ'j}}@.�6��_f%>�+#�Zė'м��"<�弧Q��n��	w��������^���(g��E���G�쭹Ί�3]��<�