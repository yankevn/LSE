��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��?�I�J��p<E?<�)��J�b�s��e��/�G�H��d������-��WM`\8�sz10�V�ꍌ�-R�-�bE&g�Z�;������{Z��R\��ؙnF[=
�w�?�FF���>T �gz���4VJ�r^A5<�&±�sPiw��W7���ĉ!��~[_�ͱ���2�V:�Fe3ݔ�9�G���T܌c^z2C䓗��j$'0N?��
ar��K�Xk�E�'�l[Z�Ѱw���#��j����RUY�b;����I�<���_��C��Y��<�	��4�I����+#4�ia�nd3u"8�TMֶ���!d��V~��N��q��2����w�����y�k���\Oy��� �� + 's���1�G�z��|��+�;n�F�Dq+
d��V��;)i+�;$�*`҂�5TYT��yI,��aql�_ x��d4H�m�6��5Q%��j|ʵ�޹zr_w&�Κ�7i���1C���K�7EoGߓ�ke�k�@1�i�;�x��K��+�ߠH��j����ռ��?r?DG���obg�2�r3F�.$�$rlq�|M�r¸�;���!�.C|of�mDC����� R0�l�.��}���ר��'���zF��_F�������o.��&��T��y.��l/Z��*��p�JH�.Yh�ˏ����t�C+BQH�V��0] {�@0�՝�w=�ia��$ĕ�l���Vdc�ǵ�����\�>�̧L5L{?7 �@ޕY��x��j	��p�
�B�: �^��&R��'d����*���%���޿���r��B;K�eJ�)�S�Ȧ%���������k�ߕ �7�7D`Qڀe���y���AZ�:J T�
\�D��q4��;�dsadˡ���Q��د�g}��SuI�����X��ԅ��d�d���� ؂�A$��?N�����Lt�чl�|C�sm��<m�C�~w���dH�3`�o�OG�l*@�p��Oq��RF6��ŗ��۲�i|��~mfpU�>�gu"�?��]�+�<{�����hB5|~�� c���<�V�s���l���l���b��0��F�
駯p�P��SW�11�U�k��L��Q�K�_���R#Vf����bZ}��5��w[�W�MͪID<p�}��ar��t��,Ad���i�E%Xm;�aе=��9d~�c��a{��bn�.�s� �
�r�u���?t�#�XP�7�i��>���C<�qR҇�1� L��wa͔������G%�m2R���;儮����``��z3�1'��c�Ȥ��ra$j<نZ�ͼz`ZQ�/[J!�,�A��My�`M9e���3w���wh'��:X&��<�I�\���k+!ɿ{����V�1x���}���;?�x�(�ؔ�r֜-RSX�%9H?�>SG�� #��הX��m�1�ڹ���4t���=��d�^Z=��.,�b/#\��W����GòO�Jq{��oP��̧s�U���UG�μ7�br����G�2�Ke�CDꑪla�{
���)sM���0��SЬ���z`�l�>�{$��pRu&y+	]����a+�Ek{>�v�v!ۇ�#�]��j��v�7� 9&'9�vbc� S D�Rg��sx��M<���D���M�N�Ȕ'�:i��, �_̉��u�|?yo���$Ǘ �&����V ���5N��� {����+]W�[$�����!H'�6xp��1#9uh�]��]�(%�����z[�I��޴R��4���RB�g��<#���tC��`���ō��V�N+������*�a�L�k��'3�SC��D��5�,-���u�d�kj�E����ĖE��S�$+��烔X�27<f�N}!�ڭ9�U=E?�̝\>��D�:}eX��x��ԓ���'���[��r���|��	�+�x�ܡR��o�v��
����.R4��I�i-h�ʯS�:1�ٵg��	�鲨��p����ͷ�����ð/��?�Pv��'~����|'�ɸ�ǛpuB���ӹ{�hj~wk1f����
Q�T,u��Q6"?GX]@~,�u�Gg�{�\�1c��݀c'�����*v�n�'/�Dq	�;Ђ!j���^���r����&?9�1��+�!奈M+w(;S r���#��<�%v�cM1���$����k��[�.�PH���ܣ���9YY6ќRW�I�$�V���#GS@Ӝ���7�b/�P�j�v����)1����egB�����osm�;�iu�^������o�a\$�U��=�2�� ����T�w�FΪ���*w�+q�����s�F���j�9|�}E�й��sD��xn�[�~;�kX*�ޯ����zo@)��?l�"v}�ڦ;��������Բ��3�x�k��e�f�L�B�sO��p��"� ?7����K=~u9o�wj�tk��d�����yi`�;��)�Ě�6R�n���	�m@;�^2��I3`{Q�J,:�f��;��^���+�C~j�X/�����8T��m�%'1t�'��=�m��l4<i����_��ʾ�֝�3ݹm�ppX3��V
�P��[F�&P�&�_G粿��3�$�d3�rΜ��|��n�[\�$I��t���EW�콤���:��c��2"��$�m�΍���˕��,��{;�E�-���F��y��<�+e
_�Љ1�7�9乔mH
�dQQ��
��X����B�C*��쫖u�XooR`݄���ȸ��I7�L�/~�!h�a�������
�����F{t��s�������v���/ڶ�J����%�9�8uc#A?<:��	E�'2�d�����ҷ���E��yPo��p��co�*���
�R��`��y�xnU�.��,a�*?/LZ:�)�D�EI��F������5������đ{X�'U�te&�:&�z�⤟��^9t�jR�YBh�J�(����z>����ki}<�=r���0,�ĩ��{x��KB�R|K�T-r:ī�d��'rYʎmhG��"��Q���)%�JЛ�VXv�o�ک�#�fL�\(J�k%��`�Q��Et_HE�o��8�����zXɎ��nv�S�e�<9�"���3f�)c<r7.�Z4���yE�����J]@1|t������I���[Pĵn�E�?�����r�47q�w �
��F����|NN�q�~]!�Z�l��j�P^�����ᣡ1���"��uȏ�����9���}��[su�seE�G�S�P���ܰ��0�8eR�JjM,v%&��{mi7�����8h�}}U p�f$rF{�х���b�����r�	%N�j����,M�F��<o����M��89�*afò$�9���?=����YŞ�y/kp��&�DQ����E�|z�#���ԥ���h�A�:����"�QM���V�f��S�7 6�j;�xA0���g���,��Tse���Λ�4�[�1���#jX��L��q&)g��=1��T�/��#�~;?�s�������#��Zߤ�?�5�����eT��PrN�N�1��A����w��Ǿ��W��[^�#�S��ɤ|j6�	uc��2V��m8f�u�*e4���ն��+���cS?�`�1hM�9�5w;�ɣN\V!��kR�=�H!�1��M9��3�[�l��)cZ-q��{��я���8����7��Y.�Y�x�a��͟��%��"�����!� J����p��z��}L��]꿇� �
�U;d�����p��`I��@���ą&����v��O}���Ũ�y/:-g]��w}ˆ��J����8��6+APS`�>]5nM��+���|�� �brr��&�e��ek��Q�i2z�#���� ��d���X\�5G��4�F9�جw��������R֦���",��ِP��VX�Bg7жh��Q�|Z����7+?W�o)�!���z�ӹt�}�G^r�W��ׅ.��~J�'��aʬʨ�K=��$U,d}�������iK�[鞄��f'
��Azo�����S�X6�_�Y�z��Mud�[�Q>�,�H�c}�(���LN�=��)m*4������2��'�� ��~9`��0=TE7�l�E��$�4{u���ґ���=^gP��4�*�PN�ô2�gH�C�a�g)C��+s�y�Dܤ;���k�S�o!(5	���#~pp�!&%FɊ �LkOPL"�$��)�#��=����U͘��Pݶ^^�]�yу�P�J'3J�:C*B7��lVdB�L�3�P�p�?	L� 3��� �۞�)6ɼ��X+���r�ꍂ��3`�ֿjv��3�����8'd.C.E�=��� �%��~�m~�\��e�4�J�E�<�9P� ͞������L����8�Q��b�~?9B$��E�Q.�x[Eşf�=V��	��oH}�Ȉńjc�YsR磷l3�?*A�ʪ	wO{?s��|W��"?(�pOB� ��z��ɸ� �Z݇(���lI�'9�(GH�h�ÞK+���@��k��Ε�cbgy��?�TW�T9�@M���|@��PQ�6K�Gk+?�k?$s�Fz�"���;ZE�Y��|��g���~3/Y�D%,������S(%m<�n�X.=��_*v�x���LeQSWS��x�-b:���i$��9����^����ز�2#���D1����j����D��K�8
g}-������^�]H���9�z��[�I׽2�:�D�>�"��ڲ*�W�г2&���%x�XةeHy���P����օNA�= I�L��LOF1-�t+W��"(T>E����-����|�OY
�S�R;1��DA־�)������é�[�cpD��n*��/�YH\w�V����L`F֕���e�c颊��M�� j�O�n�$����S���
iT3v�@{݇���k��9��������Sx�@���.���!l.��y����mU@��9@f���9x��%�Vl�#ԑ0Ԟ�Ch��K����b�r�(��W'�.�ď"�8Q��/��fw���f?�AV��]1g����O���/+��|*A`�1�7t�taϫuH�r4I�}����-���*{���+;��T����2K5b�F��Bb��
���Ce�O�-?����B�#�jyj���{����y)���g�� �4�h�v��13T��O-e�A��H�OV g0;/���	�����R��{���S!��G��5�8��}�w�If�f�f�k�X$�Eq�g#ؖ�;xV�4%E4��y�1mtޑ+�f +�C7�� F���`�&e��u����ɍ�wg��l��u$*8*��I��<w)*�}�)�cQ�1U,�=��j)���~z#�"J�ݢ&�0�v���G]y`Ьq��g�oՋH���4_&�9/C�-�i��IY��&�U������lF���d;"j���_��v��^�AcHGg�;8�Z�:������̼�ܼ�W\��z���[@�p���@�ą�'ڭ�^��A���E��\i���Stγ���<���@�l �G�E���{�L�h�/A3C��|��4L5x���Y�(�L�Jl�Ga B=�U�/F�����/��3��:���Q�'�a
�Ha>+ ��Գ[DT_��3#�*�$�Ee�HW#����q=5Q���(���>�Z�2j$g�s���X$�Ւ*��RR,�4����Db��vG���>�#��eM~%���������P�ʞ�AAׯ��>�&�4�M�)�]ST�0&� ��a~8M5�#i&主�Ə�AJO�Q7yD}���Rڀj�妮�R|�m�ό���	�-�D��ҽ����S� �����U"�d1t�'����:���!�q$<������ �j�=-��x��b�y�	
���V�&��?�^$"��9¹�!"_@X��	�u��u�뛹��@�8��9B�� ��pb(����Y�W)��9���p�$�0�����@	�E�y���IP��Ϸd���>I
-��+L�T+��e��j��o6�&��`7c�(PBE%���<���aN�&-)5�_E�AG@#IM���l���1���*1�(�wZ�fN�����S42��F��T�5�ׅ��dc2AF���Ԍ����Uq�/e�`gp����
w�?��#��������h��u��pT�t��V�҈J�xW#��d��ҵ�+c��R�)M�(H���_x�����@�"�WB���(Q �Ļ�8\���i��'VF�>�*@_a��0dA�j��3w��\��C9�qɵh�zܗ���,�W�q-�yف?�D%ȫ��ƥ�+uV
��	8�T��-�����c7�.���l���e�M鵙ܣ���u�I� �G��
�)+�����l�,Q^�{m��k!�̰+�g��}�Ŋ�0��S�Op(�M-��N�	���|m���I0�T̇3����:4��t�=I�rPyzE0]X�t�ebO.i�ud:��Ś�	3)_��J#�W�3�p���FصL��O�pf	�^t�c+�-ڭ���Ö���o��^�E���wm�4�]t#�-gO�����G�H:ԋS'|���|��g~P{E.8悽�t�LD�sڶ��F
壘5<��0s�U,&�t���]B_���d|*�ݷǽ@v����@s�m�8���z�:�>���/�d�.�E�Eh�HEbD�e�k�{��(�F�8���SA��I���ͿkS�)��e?��>|%"��d�mjs>Y9(��`:�7ַb+!���l����F���J��6��R��)I�Ye�A'9>����O��x�.�>~���f�/� H���=Vŕ��ʇ��I�#���=�FuG&�D������ �t�����?=��b�,�ːՍ1rS��9!)zK��->Ls�i���o�b �����PP�\�T��X,��@[�Ddȗ��/zl�����JO[j����۽D�O7"�I��q��t��s;� ȩ��"B��zk�������t?�Q����̷Gk�]��L�F�o�o<��4c<6��������^�:�1�[@=g�q��A�C�>��ե���}�^a敬"���=h���-t
�	 �gV��&�k���>�L����ك9���
�MMog�%�M�����ʳ�368�ߔi%^��,�ڟ�t�|��p�;���K�\:��j�7�P�T��?a��`�eB�C��x�y�L�\L`}h�ڐ��fQ-�$�Ԃ5��#�*�^��}i`�@U�k��KHދ
�m!�:RE��+���b8.Wp��k�ˋ���^S1Qm ���7Y��� �߆
u�5%�z�V�t��*�z�҈�=�����۲gނ/󽽯�����b'��"U+��GCv꘩�K�}��� .�� @��	����3�Hu�Z	ޱ��S�p�; ��cU�V΅Q��)v��B`�{��k�{2SV�����P��8z )G9b �w�6O~<l�;�2���G�ueg?y�~�q4<��L�S���j��;�:e���ɧ>�OyHu�t3�B���<[�x\a&w�j4��<��LcNJ���R��ʹ^��N>��g���X��-�Ή�n]����O�nj�s�޽'>�p� �h��C>DluT�DYt���b���kn�c�Y��5xCP�9"��]��$p�IL{KZ���v���.�T��b���� ���Z�B� %�&�x=�ޞ܌�}�E�q��m��T��ma�֖���F�S��۟��C�,�8#?:ȴ��.x?Kp��ރ(>ߺ0NƐ�G^���A'nWg
�i��}�����^�	���a]=x�
��<t��<ʦ���,y�J�௷�*�3�8��*�g�������Ԧu�U��1J�q��ǔL��O�(�I��H.���H�=�;a9ߔ�.#�� 
�^�|��$%�?JuKK�Á��_���X×|e��
m�v�����p'����p����jz���-X������@�4''���OM������K>��B1��rh0۹TX�"�DT�B�zZ�D�*X{��K�~�!���|F��� ��!?G�oX��Q<*��LF����M./6mY%����%��4�Z�!ᥳ�eH�7c�i���E8	����(��?<���谆C��D�l'�ӭ	�M^A�U,�"�!S��e��*4��#W����lF�~/7����S�L��5��T�=$eo7F�]��{,s�J`+�;�B��#�\�'3D�\�_>�ɀ��'   rw�vS�_��H�K�B�0� nl������ñ�� t�Ҍ#�d������m\�߼�!{4Ȟ@cF����6�H�O�/������o�s$�x��-=��f
�����1�����1��V�Y�9`qY]�y���ʼ{"]��k�����F|0(pi5ɹ+�8���J�p�����^j���^�=ϣT/�H�]	����] Q�I
o�q��xz'�	ޑ'p��3�M0�I+Dt�^wx�n��X �V��t�ѵ�u#\Ka�r)�|��`��a�
�ژ,�x���mIy�š���+�Z|���[#�M�W��U�B�
��گ��;#��F��g�ѷ�7�dhe&d�x2�u0\[�snP�z�,�ŕ!�J��&�,����G%���G��a��Q�6� �P0�<�W���.HR{��M	�nS��rG_ʌ�A��&d�8��ϙ3�&��������ߋ�����Ǻx�ᬄ��?L�w5P��}�Τ&R+���Z��9~�>�͡�+���l|�fBO|V|v:utU���{��t����^hB"ą�Y;M�o��j��ew5'
ܕ�p_;.�w>��9έ��X"w$�xIvE�(42U.M���&s�YBX�~�]�Tq�U�j�YHm���7\�B����1��\����=�G���"�V�<�1�;0�ID꯼X*P�Q