��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�.��ܗ��"Ä\�e�E{��#�B����+�8�~z����.৫I��e�SM�,���}8��	\���wJ�jp��L8f��͓*ܡ��X&�hqW1-a|��^�q' /ڻ�<fA�SG9��d4�*��;��\�2��ˏ+������G��	�5���8�D�c_�)`�#�1c>G�loo`G���MBڞ���-�ڭ�?ӹ��xʫ�Q��E�ӪAPh;7��O/ʨت3�М_3�J62a-9e�Hdظ6��W~�݀U�su��%�ni����;MY��6�'Қ�zG��q�ŤV5�Q#`B����q����$[#��'O�r���WGfĤ��&J���M�e]�e6;Ztc��������""�/���CvLK��%���n)����Ö���%������i�;�w�]՝������� ���<�uzB�@�q�5˂O���������s�����bS�B���y�bW1�:�N�X2y1�?bQ��J���\���I�/����(��'Jx�_:�+�6U0�j�,�0��Xt9������g0�)��,N����Y�<g���D�ؘW���ʿ�{3Q�k+��Ad��=�V�B���8�/0��� fp�7$֕�C@�B��tS�і�p}�+"�R֊\o�>!�H=	��G{w��@I�?((�x��Ox�F7~o	VRpt�]��U��"pl�/�b`7�A\���zn�G�Y~�yՊj'X��¤���ߒ8O�Fm�ӔK*`�J��~�Ӓ�/elkH!�����|7c�3�5�/>������2"3��nL0C0��5J7�8��`AYg���z�8D���`/����p���E��x��m7��
ښ���x��B`Da���n�l[�s��'�[�1�തq7ȝ�Bi����O�&���Np���7�����vzRM�_>*�����m���=�.��x�T'�]�Ѕn+�<����˧z��N9��Z��q3����|�b��0��xV��~��a����`�'���⻨��?8��o=�x ��e*\l���N�v�=S�~�z� ���F}�����D�'��0G�{��{F�� ��HL�IsS�U����O*Gh��դ�\+i�X>���*�G����H#:yxtץ�N�%�n�~�*j���lX���[��_W|+w�\����C�g��zCT�����O����+[v	��V�7��5T��O36���!�1�bһ��%3?�w�!�C)/��r�
׃IC@�0
�e�%����_L/�p8�y�q�A�����d�_u�B�f��p���P��2�ߡf.��\L�̚;�/a�2��j$i�a�Ҩ�/�ĭ�E@�`�2�7���+��ZN�}�������f��)gNX�@�E��Uv�jf[�}\$����+��.�B�s�tEfs����xm�pT�^�|�%�"�A�%!7�]��!B[Y���~�\�,��(�'uM��a�A¼&�����1�a��K����W�L�\ſ��iYMIW�Ĝr����'f����=z����҄����xG�L�m�b���cA=����Ϩh�=��M�-'k�q����[*�]�A�%�G����VPD?ťJF�4����pgiN�{$9�Od����->�A��v��e�!揢�ѽ��+���D��?I����8���P=;�^^5���Jܝ���S`�kʯ���mbeN�B������J�j�b�؈cr�<�ȝ-��.��4-������1�X�;s=��B�W���'D��@mD���`Ҽؗ2(�4�*ehwx76�PCS6���eW�L	��_���S��~Ꮽ6����5�����\t����.#���x	O����%r_0.�����:2٦u��� '�-��)�&�[�����Ot�Yt%���&KQj!�~X���a�Q,ʪ~����@F��=V�.�g#!�ʲLX_I�M�������S�� �m�����r
��H���N\�q�ID���L��c)ȿ���y�܀􎃅7�?� ���
)O9D�-�ޚo�l
��so�xX�OmN+�,�w ������?�{�f�\R��m��p+��^����=��"4�Q��O���嚟%�2�h+����u�r�(Z��`.����� m�.kZУ����J-���ڮ�������bJ%��F��{�!t�Q�����ߤSǨ�������H��8��u�D9U%$�����)*���냮�}60�(��xU���Zf@��B�o��1���n�*9��DoBY�� )HS�c�]CR^����ׂ}��,�>�}��:FKU�l��uR���,y���Q��,���>��OtDDhP�1��.&�f��\��n�ӻ�:9H����D��a7��ɪ��|Ή���>f��>�OFu@�CƗ��	'�N�%�������.��?�����0!yt���1:�/������T;I'��������c#2��s�=Ma��Is��6+��7��
�J�~�<��1��j�"'|��q�	��%�C2��zQ����#�^)����PMU=0N�I3��&�Q�*��`��k:$��%��U��������!�q �u�}�}�!6#��|=ݎ)�h�9�!�RL���:QUd�뭍�4 �a'pR���b���m�f�8�<D�Č�h8���DDi�DzY���V���&�i���D>�[���h}Ϧ��j�K��ۓ��"����� ����>
"�4�`�N=���7v�{��	���&���D��ij���]\�]�<8�ݞ$WB��7�Gא�R�>+|�\���B�@S �茟��q���(/I�l#Ω����HFJ&!Mq�l|mG,�<�^[��<��j����w�.P��;
�4�4��"����,������gJ�g
s;�*Q�
�|00�H�2��!<*�v�}�m�HP�X,<ζP���N3� Kɼ��L��E�В#V�V�+��PQ�#i
'�T��!���GA�v���M����d
����9K�k}{vyd�L�,TĽ宠�et�D
�dP%�8�Jr�܄��\�ϦF��:��R�BeM�EβrUV�-�T���t���we_s!�,��o�7�8K�#���wL6��X��f�Y8Z��M����1!��xzZ4�)��8Q��F x.�|�&˨p9��~�e��.1=zh_fLL�V��$�/+��B�
k��y�tQ�ѕ����bW�yNA�mW��ڴq�Z�l��Gx4@w�+h�"9`��z*P)�4�ՓkϮ�/�?/W2C�U�EPS�q�&���Y����<~D�c�X��G��Is��l_i�L��h����9E���T��	��m1��}�{Ln��Xsw�ٹ�C�v����y�ջ'8뒟8���u�/"y]o�ߴ�r�Ie�QWd,��9�ɫ���߽��Ȗv`�~_ ���gѧ��D�.�Ʀ���ʭ+�Xl5X��	��Z#V�亝2c�1� ���g��ʽ�Х����
����^([7��͐Z�u/�f6#��I�?Aw�bT�� �FD'm\�<��`w��]�|��ʈ�L6
� �b�{��;�q�](�i�poV|�.�����2���~�*�"5�#���go�]�����f�Z�� }JPP柽�#��̚XAV�r�.Z�J�f!{���C��al���<�/�M�\�%ːhw�J���X�3�6�X�O���Z�V��"��v�9'�����nۓ��rk �n��O�9!��T�D	F�{��������"��t�i�T�#�ő��E�6�U�|���3sT��^�7ľl f�i�9�l�e��}��ݓ5?�>��;F���y��������ZdF��6�d�ŝ~�?y����U�1����m�?��{�T��٣�j_g�NF ��ș����N����J|���0.$��m�Y��
��c��B�@�_a�Q�l"�Р���}DKw�@U1r}1ɣ��ğ�aj+���8 ��~u��BH$w�e)v(o����4D��xU+�4#��������槑��a_R���2R����n^|Ԝ�l���T����~wd�GR5���	�e����$�}8=;�D�˟zj�8o/߇�X�{���� ���6sBE��l`� ��G͸4�K���`����4Ո�K);����@����p�T�(C1f�{0O�Z��h�p� LI�a�9�����#�������T?њ��C�{ȂdFQ�Xu���[�7���b��]2��_�M%�]'�Db�:rQ3HL������j��\���1��s�e���R�H��_�����
��"����b!��Ӈ"GFx�?\�� �#>��cz�l_�fS;�mψW�	��
���NFʵ|z�`�w���y�p����Eb�|�Pّ	�� D������\.�M�mz6��f��}RD~��#��0�9dX���;௓{w�o����0
}5=�J����p	@���������\']�(i3���0�V�V�w}k�P�*?Q�Ƨ���ސ�j����p�͆��g��v��۬��J��$���/4�-IDM)���ᵶ#���z�6���p��V�ߓ��Re759�N���
~�6���
��;�\��ˋ��`����]���G=�~i	�3��Y�~�����V����18���f�)�~Q������N����®r�&A�o���|�0���5V�rk#�:j����G�E�xxa�%�0����������n��R�(wo�m�>{�q�!Xȴf��2�KBO��uiǯB��r~�%NH��J�|��a�F�/��ʓ��S��|��K� ��#�lSO�}����l����^��a3�nj�n~�͏�W�zd/�����ԓ���^<������ ~0�A-�xC�1i�&�Y�����Xm�L��z��
��u�0j����G���^�Am�ƾ�,Yѓ�~ɍ�A���~.=߷gCD� �1��ko���s5M�E0me����q�1�iZ�9Պ�76�v�e������du��oM�����e���roǌ��;�hS�1�� �"X
j2�	�[�+ Z��Y�'���?(�@�hĀ�1O������$a�.UWu��N�|s�*��C�UXM��/��
�G
q2��I�PE�h�дLJ����G�+�}=AU��f��r�L|��z�EL��-ɧ�8դ�d�u�gS��J��Z��p��Y����d��5	,���f�ς�F��2�/z��#�^�u�⍗r����$��<]���`���߉�#Iu^
�j���bEș�8i���7�VS���橠����o�Eik/p�Y|�Mr��!58���8��W�5�QL/mdk���5q�<�f��/ˆ�ۖ(��<�h�XC�>X~�B�Ɇ X�_\��������|����3��e�:���=?�y��8bH�^\��"o��8��6,��_B"�rR��q6�|=�<�nMy~��{������K�����p S����+�J�B��M	t�`�f�ˢ:�ơ�nLu���]*��f�-������R�.�93�0j�c/:�F)}��L��*��^<�j�e}��l�pHw��rz�9�q��{P�:�2DG�7��c�i�⣙��Кm7��Q�/X�}�W�g�q�!<�a-�pe��,�h�G�h'b��v]w�AAW�)z�����yku �)+��[��릆�y�"���I��?˶���$e�����%�͵�.��Ȑ�`�E��j��EV���� ��!�N?��[0��K�2���L��7�~?9��6�_>
�*D-VP|��6����̋������I9a=:#g-��%І�0X��Ƶ���O@��6L3{��v�w�	����7���X|�
�H��@a/����4aI������'�u���o�#�~��TB���<qvh�`їu��B ��8cj�OG@g,���mkR V�փU�O�J�M�D�{&-��._Y�1l����Y��1\�6�D>]a
rMwg,H��#a����b�"_w���[d@���Ϻʋ��PV��(N�^]�����U��U�������*����ŏQe"bQ�#�5��_ۨ�0�%����_}�������@���l�(P<�#��Mt%ה���o�~̱e���D�5���U�2��=