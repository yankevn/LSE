��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���ORwǌ��{`�E;l5�/�|b�Fige=�@��.j���\�6w��b�ʘ�}2�7��G���d�V�%rh��u�9��i�E5�g�LL��*L]�¹���0��7��}�;�۫��hE2g1��$nG��~��4CD�$�0�Ӑ7XA��C��� ���Y����n��Q֏��z�͗����
�Pd��&����ء���c�TG�N��~陂������c)Qq-/����B!p�,��8�e�o��u��<���\c���ި�2�Z�I^��f��w�7�����=�h�O`��� :��~�r�K���D���n�4��h\�/�ȓ�\`:a���6w���vn�����q�r����^+�$k���5|�*�-u�EG���|J�ÐyX�ѥ��1h3`]��զ#�\'hm�_[�r��!O��'?�~ذ7-�;9�=r��{.�$�ݱ�����Q���o�~$N�����R6������o�Ak:��׬α�Y=��\���k��Z�(�0Vgfd�?��W�V~��1�E����*���s���kQ�y����VC3�w�n�J�`�W�b��j9�F��*o��74�m��bY*� ���#�i���pt�b`6�dRb�i)�o�pHB�S��;Q��U�L��vfX�\�N�s���d��U��|��͂lVxaf6k��F��2�ÔKqe.r���K�s�Sd���P�!�9r����N�*���Ͳ;�5؛�q��t���IF�XEn�C�ݲ��=��2��ְ�R��c̢I�Р�_��� sU��|>ל܃�/8dA���5�G&�*�� ��R����a@v�$�'S�ž���
�?���XM3�m����<�eBx�w�q'�R��f��l2#�3�8��@9��a��Qe ��U�@��yR�H����rC��,6���.f�4�Q�<E!4��4PF�}��(L��k[<c)��$�m�P��{��燰�\D?�3BM_���Ӵa��a��a���dC��PX�M��;�7�/��O5�Y��#p���'�h,9G	9�Xa[q�9='4�c����S�VUn��O�&i�[�ZF����ڜRd7f� ī������hI�L�nMlO����i��Mw�A�J����+w:p%,`ɑf.;=R�5�+)!�l��ry��R�Ze�j�|S� ����;�k�����E�����Oc����6��r#���|p�Na`'z䤫����R���_'���ȝ��P*�N]�K���0�H��7�;.E���yu�Ѓ�����N���5|����X2-1�uy��)^ԗ0�P�\].B�÷d��-���bZF���B�%�+?���B�]Nx����Re�YP@���{Ӎ��rL	�#�.=@����4�ˍ�`Y���'�^�0!�`ϣ�p�!t�=P�
SFQ1�,g��_HP]	 �?���@I��qư�P�CLg��z��:���m�g��^���SZ	Q��a�?���2FW2z��;��~��v9�'�l�\`��<ϙ�3ͱh�{V9���\ľ�����Y�����uע��~��yk �%�cB��:dgѩ��l�i���D����e/!U�51�$�
dTa����&�/�~"�#�����\d�R0{K�RYC�xD�Wj�Ǯ:�)�?M����@4qʤc�:8sp��P�IjS�a�f>B��n_J@p�T��x:���Q��������_�������ݏ��h�T�V�e�p�����׃6a��`&���
�5kA�&6�;-x�?y/G!w���cKBE7@�\�����:�F����/5'�d�(���;�5���E�efh$���U~
�+����Z�Ͷvz�����)[�I��ȧ�_��&?^�o��{��7~����G�L^�P�������W���������^�,zA���d�F���� ����,.�Y��>[�4��� �u���w�NxC�A/�x��{뀇"0;��� �F�%�-2|�41�~qf#�TJ��)^���=����D[c.�{����v��OQV�5�rxZ�_)��ܲ�jj<AO�[�v�����'� Y7��|!���8N<�R��2�0����\�e� ��1�Xa��x4�)��H��vjr���`(g�p�#0�`�����o)���M@E(PI/Fk��6g�"��l����^fdj�l�WA>MM{��BKڕ��.-y}�h^�����E xձ
�F��x���.�p|H%_+?�3��Q����0>a��xk�|��_��o[�1od����E�;yU�0>��o ׌{ڲ��/~�0�@����/�����}�� ��2�Q�(�Y��vhG�y�(KiY����N��x�{�Ϸ�ft|0���)-�q���m������T��h<���mr3����jE���"����g�����䵱��m��%[���y(Z��tD�'��Y"L��#ep�����5���V$�ǩ�y5 �CN]V/���7C�����>kס�2��ߍS������"VB,������H�|kz�?���)�bL����Iq����*�&���Lq�{��0�H�~��ʏ����^�����2�B=��i[��p�ט�����P{�	�(��x���d���|߫dR��n7���a�wHJ�L��b��ܷ�D���u��O�|Y�v�&|�U���P���!�]a��xdH�}�x�=�b;7�IN����k���Ċ�ƃ���Ȁ�h*?��g[��=)p&��c���,�&ᄕ]mc�?�!0
G�m�Ū�8�N�(	��L-�)������F���՞�k�]��E�� �c/��|��]����V�4V����5��ϛ&ݾ�_��1��I�e�fL�duJ�%��L���6-��)n��˵�
X�Y�pt���8+�������i��)A�m`:N��`�R#=-��wcT�U��hY!�{`�O+����5;�12��%3I��2G~o2'|X>A s2�_��(�(�%��J�H놷�=�*7�I����SMe�Q���ö��M��A�V���Ag�����I���S!��|���{�5�`:zO�+|�d�lx�����ڶ�Ðꋼds^_G��Y���6��ᱷᾟD� 1��ȉ����	��~�^ܱ��X`e�_O3ց/���%SD�▤l%p}(F��J�� � � �*?����KIP�-�ll��=-Z�P��bA��X���oy*��Nqɒ(x���9�\����:�թ&q%�����t�7Z��0���9C Β���I܀�"�E3p_��C}m'꼿̳C�C�6x/���O?oe��I5�"�>��%z��|h�[��08{�TE޶���N�cDU��&e
���9ޠ`~U(p��nVY�O�"+�1�m�}����j4�#�����]�&0k>�Ja-���ؖ��I����Ǭp�~�m�� ̛H�)�K�A:�4K�N(sϫX&�ڙ�
=���tb�vEd���q�}�ܱ��	E�q����Vu�/s.�7���M�SD�.qz*(�g�%�Zj�Ҙ�x��X�($�ɿi�@��x?���à�	�Kk��oќ&���P�1�&������b����W�m�ҭ;�A�}�0�|%�sq�1��G�ru`VT<���ʁS�'K�K4�Q���]��f���"<�[�Q���@oDf������In�v&po��U��ڠ�E��m��3�����4�fፃ�/��^�������PtEsʤ���'a"(�`g��Z���A�譭��e��b����A~����^�-z��VE�G�1q���'��eӝ��X�׆�`����獀�v�5%쎌e����p��32'w��m�˶:)�����au[9�Iύ93��N�Zd����̸^CA�uվ����D���>�5 =��Ϳ����T�Z�4�pW���ĵ�%}�cǰ0]�/$�� �+��V�yګê�2��ݹ 9ط��z�$6{-�1p	&a0��tp��7�vqb�C���e��|���
3��k��8�5�8�˞��f��"^��rh��'o���H���:�J��G"1�}��@[�5����2�viʠ��	D^sД�NZ� ��{�M�� �/9��s3����l!�ȩŎ;�L�E��&�Y�>���������h8�R�mw�<2�PX`-�
{�
��B�6X��)?\������{u�k�~�n�f�i����Ȥ�N�f�/��]C6Ah=\�$�N��K�n>C_����Yy���Hu�V2�:=��AN�q�kj�&�Ύ���J$��fN��/�;f߹J�
d'a���{�PW�o�\+LK�٦|1����#�|4�X"���$�v2�켴�N�E��o�l$Y/@����X��!�a0p%˟3�vݱa?9k:SYZo�������	�\9q������l�:�܎>Z��M1���๼��=����r�a�n�}�rP ўA���*�N�Y����˰����,@����W�9O�IV)sP �[x�o���Ư �L�؅���,���~��A�(se|.��r�3�/Z"	̦��f������V��g���.���j�1�C���k�..w�9��0�CȌh��숂�8�v���Pq��=k��'�KBe�!����r��}�����ה��Gtr\ߣ���32��� ��oJZmN��p��C�;���(�����Y#�}��q��O�� 1�<�2���i4ڸ�M}��y����>�0�~T��(u(0Q���l��
8X�>l��`��H�	k�a������@��aa��ٝ=�w֯;�-j�M�+�c$��<܅��q�#��g�F�5�b��T� &��N�O���EB�mb�[p�"p�ucej��C��h�h�r_�x���$.?����^�D��c���O�X{l2��ᛓ�wk�Yay=�=U���7����G#s)�ܿ�2.�DVg�I��0?�V���~����v(���Zf�]�IvL"����gN���FǰQ�5O��io��'��U��.���-�9b�ec��B�g��Ы㍎��X�{�]~Z��.m_��;��KTK��`��j�o�����l~� �ُ !uӣz<�]	L̯{>7�c:O��>IБ1N3 c���T(ٸ~��Q<*�-���F�������l��*/�u������c�D�23Z���D�2�H(F{�%pFuF"o�J&���Q����$]ߡ�;���]��>��9563����J�e�枃�3 ������T��1	�Pl�׏Ǚ��r`j~�z�W�)��1��D����Rx�a��	��&ڲ
ܚ(�sn@�m�?4��D,c�n%�����q3��8���7�*��Ů���G���E�
z���S��h���� �5�|p�j9N�S��1�N޿�`��!��/�\�=�O�Z�h�Uc���Uv��1a_4�iޭ��+E�P� U��`q��z��3U	R�ʿ� �7F%&��r��\����L|q�Fɝ��;J���s��/�M=d��8Y�f���z��vqNa�(�A �l>ʉ���2��@75f�zpe�dP�2�i��y����N����Hn�S�J���B��G��dܾ�,"�q67�އ�Z�b�U�*�~MƤ�y���n!���z�����EH2�A��N !
���n�l��0x�����ڛ�!��_>��$ 0� f�������#腵�-��z�F�{;{�h�lw�D�VB$�_t<�2#��|=��?+����V%���ѕ�_�scd�ĭ6[�_���w�V�#�&x=y��G�o�3N�4��nwzb8�:ZȫD�
���V&١q֟�h�ØS8@��ׅ�S��R��%��amN���Z2<S=�Pph���k���hT�2F���"[R�X��g��|n����hq��Z#)ed��)	4��|A��=����;����2;G��������K���Ї�� �[g6���GK�]�c��bI`�����:�t9u�P%�#��3���j	��p�� �x��$$r^�fVp�E��7&%�_:�X�y3f{�f +|�� �j�K�<5���F���'�ċ�E���ȉ���Œ�HJH�&���+[�Y�.��m�N�n�?̗�������go�M��d ��X�����|����ʄ]X���|�{r����ά��yɮ���R�,U��z��`i)&���nm��,��Wtʈ�?>�A����	jt�Y����mص�qw&�{�xLv�V�/7�"��+���u�I��n��f\zo�r��ƨv�da��#žX42��	�R����_̌��t�V}n��{�sԘ�_v��������lb>�[PG8N,uI#z�H�}��<6�J���dI�
	�pX��3�~�m�Yuty`,�<��/���5��s�R�.4z�2��[eTM����G��Q%�/EoA5I%x����"���L�]�-Of���ypW�]����[H�n>��ZM��[ዻ}V*����6�N�;&���whl�?8.D/�`$o�ك��F�|��b�L���̋Y�n�� [Z���)��Q؅�{Y
�1��ӂ�K�;�>�����,��ح��Sn���T���������=%�J��7�[̘xW�|_�(>���E
�	�]iq>��V<l�!�e�X[���y"�=U��������]s�2~;{��M�Z���74́jqy�2���T�S�ndt�.d�C��cj�)�� �����
ci���G�.0�Q�cI$\�F ����Wz ��"�ޔ�Ň0�1���,��d�����?KQ�Fև5�����ۘv���8��ﯵ��@w��yн�ҏ���8�[�˭�r��g��v��N��vɬ���'j�2���ˎ�8Q��F���1z �|+�i��9f�k��x�)1_(z�'�F��z����/���7��'���e|�{v-���I�P�N�q~����{�,S �#��
�".l+s�)���۹�~h�]���ΉAl�ie�+q_ɪ���Tt������O�UW!6�̡L�Ƨ��g�/���j��\��pt��7i���Qz�>f�9<�X�AG�� [#un/:���"�3I�-4��N�~)!q��8���%�>�P�
jz�}�f���`21H��MEh�}�o�sF�2@�������N4�eI	���bj�S
b%����V�_3&*�,1G�DFf�e+Br�\n�[�'h��k6� 9z�:,���C�Ō�Y+�ks��MP�.��`��&<q���Ƙ���s�M��p�<�'W���M��|��#����D�$�����6_z���A�J�
iN��:�1�W���)2�.��ū�1�A�W���<��+{@D��-�4 �9��]d�;x�#�;��Zc|E�2�\�jo]�0+g�!����r'4ȇ�ê�ז�G�Ր�S���4ǽ\�Vhk��b���Þ��^����#~L�r��	����aok	��B��55��֕e���I������B��K���ot�R�G���dT�ې��	?9?����N��ʜ||���*0d�8�����_B�aGT�U���a�,�n���ɓ%��Rڹ����Lf=�TU#�/�Z�^��:Wf>�o����tQe.�\9��8�&��M'B��<'s!�R�b-I�y����x=���ߝ��L���g�vs]���	�u�G��;Ϟ���:?�_�S5�{�M�6ȡ���C�ƘJ��L�,����^����@�v
��D�ɟ�č���8J�$�t����}�4^BR��1���&�����P�KgyfD���l9�������Mȥ����m����d�,)�8m����z�m��$kLs�"�v�l�n3.�����F�i���=6=�۪�"ۑ�#,������L�G}�I�$�	%f}�wMk]:g���:A�ϫ�fG>�:>�s^��Q��ĪXgM�4ߛ�I.�]=ѿ��9���\jr�|$º7�,gQϟ|��2:���X⭻���5�=���EL�a��7��z\�jf�{u���l�4�a��һ,�R��4?!��#0�̹���%� %�Y�Cv<o�x����U�o�¨��dT���y��L~N#�j�։��DZ{���TFJ���ʌ۠&T��xQd1$r�6�*����!�����='����%am��g��&�BQ��2���r��љ�]�v���vgKI�?�D�g�J�ږ��h20�lӽ��6q|_(��ٟ�Uý9`��￿��-ϭ���(;"8}�?s?��f#nS���g�#�3���U�^����fjaZ���Đ|����-r�P�fr/}����dM�s�
�Eb%�1��/sފ�m?�G�D�O�q�_+0\�#= ��Hj� {.zYB��"�DzI�Vu����[uzz��^ҳ|���=�\��Q�C���>����I��sO���/ �
RIqa״�+,HӗЩ����Ȉ�_����;�N8nr3���\O�tb<���x.���G��h�Ę�)Q�X!+�� x��6���EģK�����hșd�����N�7�eH�6�; �w֣]�Ɲ�ٸ��|�����5cjxќ�\�� ���W��h�D����oS'�/)XvrE~�#̮�(��ӎ�v0-H�kD�t6C,3v/�D$sp�R����_�T�-`���3�ՄK�2~&;�$m/������Y�a�'O������H�_�b��kC�̩��X&g�ʞ��ކ_��?�i�˻��߀��<\]]O�
���'�!O(h�>,6�����m�����4x|��6U�H%���P�����U��5�Zq�o'�:@�?�4Bƨ�8��4�[��v�t�P��/Q���sRqlצVRiBk�-ֹp�1A�3�2|*�2� 0_˕<��=y�ɹO ��\$Т��u��H1Z���2�u&Z��4����i	0t�f��:ϣ�c�u����sfr�|9�Vu���f(��S�5�z��a.����mn#y�����=���1�CB�7�n� �&-�Zګ6CUZ�Cd�TK�%�(Q=`�,,��@ݜ��@����{�I���Հ��u�`	�y��G b�B��)t)�)*�{?T2�QP��<I0�p0�#���������4�Ã�w�ZD���5񵐫/@��/�����X��&\b�����C�� O�R�7P�P�Q��1�iV;~&}���g��ѡ~Ѐ<X��_�X3_��*ܰ�����;k	�l�P	���	���}�]��Vg2C�P��d6'}�Z����c�Ҹ�IL���7�[Zq��)� �&�4E0�Tn&F�5{lϢO��a���7%���l���G�W9� �5���f�\�N�,��M�R�W;�>�n�rL�z ��H�rb�wR�ٜ��k�E'� ˓f;�EM0O(�;D)[B8��M/o���k����9�	���l�Q���R�"�Z���7"��9�5M���������
���J��Y&���u9��>ȧ�]v׫�Ϋ`�W�]�t%���2�ڥ��@��d��p��r��]���F3P_�y�x�E����.�@˧���y+/W��l��3J���*���R�K�h�`&yc}���/U'prrV���k�KZ����
1��#*��Tk�Qz,A�瀡�Ͻ����:$h����چ�P���F�'�[��+[P<��V�\d.�;���%t�j.�����?���V�P���7��W�ފϢt���m�&�6����&w�}�8��ݭ��٬����r&�O�i��m�n�XY�u��YR�s�>1��T���_��׼yGXZ
ki��\%�7�&E�d�nr��D4�M�7	B���s����D��t0ļ���Bb&�N�z��Y��B~� �9��b/����`��u٢�����R��������k��K]]s%�C�2��84���k@��������-����h� p/�t�i3[���2u7�W��$G��0���g9�vMg��F��Q�f�=6%U^�J�4�� ��@����|�)ӷL"���=�F�+���~��[Jݍ��7Y��6}H���AF�iJ$��p���%/����^��0��N�j!*5����޳[�J��@~�M��zq�al��%����W��S}b�p��?�f�����:	f. v�e��d[�2�8�KX4ݴN�1���pT5P27C:�}��+�ꭗ�cuX����h��tk|qNͽC�Mk0s��ZU���Խ��$8di
�b��T�Ix)��c���mC3�Z)DE��zRW��n�}'׷Sg���]k%]���f���w��Zm�yX�w��&�֒��R���9�&eb�kı
��f��`���t��,��n�Dɮ�p�f�8�l#vk/��,zO��mʆҐ&j���@h"��D���l�XL>jy�Ss̗�	k��{�ƥ�D ��]A�1�02>E�=��4CHk�z�W��>G?����?�P��8ƭn[�]��$�K��Y:��>ι>׏t�dCU �/j���?�/�>W01����y�I�����]Y�G���;�����?��3�O���������ң���G�A�|���u�M8��!���FK�*�-�CЏ�ks�D����ړ�"h�l�"��]�5�2٨E{�ޑ�6����~p;>a�P؝�Q�O�|-k�	� []��5~�3�̻��G+���XVY��/F��1
����3c� ���v�q��2nBLX����H4�c�Wv�A�N�P����,��γ��j��)��n�"C��4������ںi�ܾ��$i����ݩ�F�@;�K+F�h(���<�$^N�»�%}KԽ��2Fj�����&on�@��V���7�X�>�� 0��
eW~������o/��$r��q���w2���G[Ȕ����v�cW�����=�>����o��=u�/���㽛ST������i./����:>)�	M���_6��cZ�xMٚ�cV���X:�Z���F�8��S�^5���(GE���;����4D7c^���@@�]���W��������f���|�F�ò|���PH�c�s$V'�j7P�h#<�&��5��#A|z��Ê:s��ui(���fu?�?�Fi�����I~�����(��z/~�X���^�2t�h�-�T�H�C�nx�s4 Ѫ��.D���D�S!ޑ\�-�3|�X�T�lUĮB�U���A�4�8[���Fi^HD"��Q#����P�B7���9����p៨���M�e#���S�"�8̤��d�tՅƙ��c��u]H�����V���erF���mQ��i��>������G�Uך�H���)|�yv�\0�m��0�+��[��������e��ܺ3�в���Jٯֹ��/�$��bƾ�]��ņ��p��X��6NwP���^����Tcn���4�D&���xQ��15\�q�F�6����e	n7SO�X�d�n�K�"�w��|xL�0���!-8D3h2?�QJ�B��5/���,K��;��C-��xۀvKyRp��Xw��;�~o�>�c���oyh!
�:�V�v2v��I���4�:K�,��})�۪�{W\\	F)�����6D�@"sf�$�P���vQ�����)�Q;�9=��I��U�k��y�we�S� w�yh<����J���j�\C��P���1 S�����y��"�"���T=��>������F_*������+�0�m' C� ����Q����`� 87�!$���dы��gA��0}����y���#N��{䉞��_#���>��g.F�O��u�ܛ������	s����/&lI������v�0�#��X�v��SədZ�j�a���v�*�kp��qƿj����*�w���RcJ�;[1�T����艈pf��i5����{I�1� � �L S�e�� i��ƇK��xE� ��mm l�,H ;4 �QN�Ԏ��M�q��9�]�S���Q��d|SuU��R���\�r��g�aG�;�͘�� �f��V��%NZ�%��1���������4���GXE�;)0�-���<�ȧ��,���:W����V��C��1Ϙ���j"
��{u��8�0����Y�g6ӧ҉ d�E6)N��&�]�5��U ��b/��y�輜	�&�����b�ɓɽ!�[�L��͸��KgZ<�Y�^�T�ԯ�! �1%���'%L�{�sR!Haq|�c�c�f�D"�W�-�lF�dx�p-�:�fc�n��5o�!�-���������X��KCN�~�o�2��k�(E������Hȟl�	nz-�F`nF6��*�8�O��*<��B{Հ�~2խ��A <��pO[���M�5P$�]�"���	�sK��.�ŝ+;��_��ߜ����W���IT�f?��֬�QyJs+�G�#��(���Z�y8F�3_�֐>��'Υy���Ř�_�s�)ɉ��fz}�H ^Ԁ�PX�W�h���V-;��bT���)UT�L ���і�S'4ў �g`Yz�t'D/�|�޺��{T�і
'/�
����~�q?~�O�[yB>�J�bq�3��8�gѮ[�yfm�ez¢���\�o���Y�q��[���VTEGb�"&5{.F#$������w[��.V}	��m@�N�p����ev 5	M���%~�j���x���5�c�J~��h[���H�T�%�
�qk��x��ϒ��E��Bϵ���_���{D(�9z�D�ϒ�.E��[�W�ۻ<j��b����m�� J�A~B����y�"�}CV3�B�X�$��v1��w�ۚb` omp0��ɽ����(�Xn��`�5��[5���`{��Կ�ILSDS�*�(�<Ƶs��( ��t��j����Q�2����R��+1=��s�D]w��tN�k6��
�O)z�D+�J�l���j�����K����s窴��b(�d��P�O�H�(�4)=b�������	?I~Os:��._��s�£Z"�ǀi��V�/؆�쇕�C-s���.�h�D�(L:�����Ĭ���i@�G������I����Fy.����OP�<Ԇɤj\�����*��Q>|�'!� m\�� r�z�|8;�>Mf�Aڤ��[U�w-��rkS���4��l�����J2/���Ln��J3Aje�]sr�LK�!.�X�~�]�ɫx���#[�w8&�._��h{�hQ[���ط��Ͻ�'g�{�����H�/w�a35������Ht��#��٥T�Cͽ�毞|ӧ�6��Wf_ڤ��k��;�d�q��q�
	{y�<�>+�z����~�(e�s��Fq@|[�d�q�ME��l�T��ڶO������4ks�</\b%�-�r�����8�r_��!���P�V!��6ȝ?�V��n'���d��<����F�T������Sf�\�eY��c[��ӗ�n��WN�Uhb�wpJ��������tk����M��+�����J	�A$�^Ws~���
B3@2Þ>�9v�=����l]L�)�J����ؿ)q��%J'�Hp`�	c��q���O2���P0��A��U���O~����SyЃ�8�#|�L���U���24&��&� �3@O��W|�����Ih��W
lNF�jO=�5 �{*�M� �b�ը�<�ؠО%'D!`MN�N.{�ŉT� ���U[h�nl�y��d��%��4�I�Jzb��Bu��G6R��#�&��-�<�>�e��AA�t�X��gB��g�JA�q�j�9�aD'V���3���Iq��Mw4+p��MhS(së��=�&��wV��E(gE�PNw�b�kٽ����}t4c��b���<�+��&��*@'�J-�����b�>��l�۪5�oب�gI��X�"˔K�j�7��%M�w��M|v��[3��d�P�}+hB��z΅�M3�_c�����|G 1G�+Z�o�|�	���vL�h���)�4��w����MCj@+y�q����b�\�[�(JtL�����UC�:v�:7�
��]s|��)[�*����9��1������u1�}�&$�,u�pFA|��DY���o8l�\�����m��V�~�T��ޝ4��aFJR��ץ��6��N_�k[$Ʃy'pSק��Q����`>k8�y�b,�DiP�$�V�!�*BK�OF���Ru��Ĩ�D�}���]������T�w�,�E���h�5���E%�+w� �l.��7F�,j7u)O�TJ�h��|�C��kRu���*ae�����w=��3y4	ʹ���@�{R/z����s��}Q�����pS�'|(Z0���8�� j=� 1&d��2S@��z�&_g��H��Z��c�sL$�KQ�1Q�G��B�oz����Oa��]�R��כ@I�`2��{օ���}��̖���C���<����D��`鳱Ƕb*�����c({�i�����>�.sw�m���Pe�\�Z�V�"$�R�봘����c��!�S_�L��f�T͒Y�h�2a#$5;����2�چF�����H�0W�o8�}=��HP���p��dAȡ��П������pd�ja#$�뭰ưȖ{ڵGoo1�ֳ�Nh�6��~�)8(S#�AA���-��;(\5�S�y%�:B��IȀa\���� �qP<��\��q���*��S<q��,2E�S����B���0�E���
P�Ӫu�{Q�(����Fs������ҹW5wG��b:xա�eT���ja���m%�'9;�I���V��?Z������j�pS�nQ���<�dR��n�/5W@����*T��U�	�CY2s8Z�X�Vz�y�<�Ү�-��g�)������n#azxkkD���>� Ut�u$�dn�SR(�"�۶Ȕ,���	�È���cR	���i�㒍���r�L2|�󳞀P�����L�Op9|q��kcPmJ�*U�Aa�(n��pI��
�ӎE^E��C�����\:ȋ�+�Ώ�uE�hpf~2,��X���'x<�h��.�V����� �T<|U|�D�L�N3��/���92W}��˳���k�^�2�:{W�`�Oݾ@-L��}��퓃��RU�t���7��o��~�)����&:mn�<�.����M#�t��:��1�3M�a;esC9>�(���V!�<�`'�������:����=��p�<�c����h�I�:���R��j#��"e��]Vf�UTh1�G�* ar�E
P�M�ʩ�3ٱ���}F����`�iH�X�I6��C��M=�G�=*�,��B-�YĳVet��o~P��9�m�a2�d��B����:µ��Bkl����q�W���Rc���䲎;�#��'A���&4�c���מ�K�<Pe��^�,�o�ӕ�گx�+ᾚҗ�R"��D5�¼�����a(�F���,� �N;�����G�,����˴��,��qL�Q�Gȿ!C��/��Ռ��p�ϙX��uS����"<
���)/��ڃ�_u)(��t�q��n[�i�۬�����BG>�y>��!��1�=��ge���)Q:�H#`
���(5r���b~2Jr
�u���p���}�|�(ܹ>"�+�)c���tNR:ﾡi��Z��'�#�S�5�'5D�'@۾�.;hAY*:�b��p�O����&����8�d�W�y�&��vc<ke�T/�����h:��(p�������<ؿ�Γ�T)���ft�S�s�l6p%�-�;Zk��W�����n{vX�7�ه���,BcɀrO�V󫕜�E��"/*�� �2O�#\���Ú��Y��Z܍�a㙛��H�~��d5��;�oc�nR���`N�(�d[��n�#��po�n��r��	m� �?q�=�S�k�x����<aż�aB��0��>f�_�
�>�Ȭ9�� �|�`���H����+���2�Q�.�۝v[o�|d�<�'(���A�����U ��*� ƋfqnG��)�U���� G�=���
y�B8O|�iS��#3�ǜ��cX�h��w�ǩ�p[�@(ߚM��6�J4��"i�$(�m�p�V�j[�mT»W3U�����a4����7������������)����$x4F��\e�c�emDb�3�7&(Re��^���+.��l�#�T),|M�BB¬ԊA�?�9I��N�<u��c��Ĭ��|:������$M�P����@^��{W.�d��< �7�$Hՠ:��C��Y���-eA`0�-֦{K�W|5�`��r���Z���a)�N���n�m�L��� ���Mm�� � �k;J%�2L(�`2��pD\o����,��<u��ih����V�ʂ���Dć����O=��!
[����1�E2)�ͿB�?�ܿ��]���	)B��c_p�h�[����~,���z�Md���+��*[	q��:�C����r�ȼ�;���^$=~I��;7{@���Kv��@F�s7[V�ިR�﷮��X�1ؾ]��]�cG�����x1�G�	�GYO/2��O. 5���n��[s �j�l��.���)<H��f� �J�����"����F1.�����9S&��XgH1\J��|<�_��5F#{	�7&�]��S���$��gu0$ِ�N��B~���^�Q��4�c�PQ�H��U�I�\*����d#���P����8����ҍ�޹�~x�"m��P�KyT��t���}�3�i������2���8���5���	}���^������G��0 %t����V�i��Äeh�3���«4���Lj�C5A�aR;��'���n�%9�� �J���o� )�~�>���g�`�xJ��֝)w|���y0p��m5�B���zj�/Կ:O��I�_�O�.���s��E�vb:�p�R�$M����Q\��޴\�>V0��Mu��@�{'e5`΃ϰ�����˳4�7q�� �
XtAV�=Z�VK0����z{EJ�\t]k�O��O�濿��5q��}��쇧�w�˨p���8f
��P<�b G����@�e�sz���.�Q#�o.Xě��Dچ���÷�
�1�&]�$(���L�b�� �p��)��_�l��7[9���K(�;�G������!\ȶ�΂]����ޘ{��{���Z��HÍK]��0@�F��&��9�XӴ=?+r����gv,�z��^�h� í7m�LB���?D��,����\7�zx���+��U?`�v�,����mWǳ�$�ǹ��gg������OO)0�	}�?r⫽�m�\��{ϧ�0im*�Q�CjR�3i�w����u���#�C�iw#���Z���u�?�M�%	�1b g�G��
-�	L߫(�3Ol���<�a	-I��jx�D!��	>��6<��%�9ܔ9��nH@zT�Qk�ƍ9�4�vg�����}�t���q�Q�ǁ~��@w����ӱ�N����Z�k�]�'r�[�w;��gϱ)���R�����ǎ/{ȣEMo�g!�����>��/R�r%�L5�错�s���8{K�n��[�i�DP*�f!s�\��iV��'��)����et�t|� ������;�����7 ��W�qf<���b-��A���.��PHh�QkP�3�v���n��;4n�"�Y'���2�� @�y�X*�)�����k��:�Ff����@謁F���|T#�~˾�ٞG�b=�}��>���� 4J3��bv���v�*��]���b*M�%�u�:;Zqy�������~���1�ȼޔ"��:֠��Bk�w��gN�z�tĺy�!eA]��H`"��fynm-~F
�M"�5���ޟL����u���Po[aJZ�6A��-إ`|�����!��O.�E塀�m}�Z�.���u��j�U���,�B�:se�΁�|�X���p*ף5�d����T�z�{�4��BU̥��^a>�"��={��8}O��0%�ʃ�H�	�>sm#��k;B��k
>��M�~�`7p���a�-��c�Y/>�[�� ��{�0�[�?&dW�� ^��t��"Dp&�n*���ݲכj����ՠRC9f��;>9砞XsL�N�����O��Lb�*�Q����D~R^FEj��|�B���^�����a��� �h}=��:)���^�yiͶFp� ��'V��x�����������m��;T�3a��v� ����oF1f�d,� �>af��,T��H�zNb�b���T�}!����疎����A�������5��]Ϣ1aV��*�׌�LJ���zJ�G��_FΈ���rib��Au	AVX9��[r����a�Һgf��r� H��Q"���	����Z�^��ix�+�n�OP�u�B���}�ίr�T��#d��]�z+`����A���	K$�6�/���Q6�����1��Y�Η�/e�>������jj��@U�_54{?z�p�}9���0���'7�P�$u��&J�M�I�4�|���5W�RARMq6)�Q�������S8w �Mt�m�����x��|0k�y�6!�"�F��uS�S'�1�@hi�2�٪I���LW� _�.�����BA1W�+��\�������*�����{I[z���
U�h2i��x��P�Y��2L:���E����?/�t ������qQ�m�p�bQ�bz��g ����lR��I�_-&��Ғ�g���v���N�1_[}n��u{<���M�fo,�;�k�ڷ�1
��A_/d$��
Hcr��G��gq1H���� ��ص��L׆,�HE��/Ɍ�ڬA��,��ѣ��l+4�&tc,O����~����YO}[��&2/�m��e�<�_&}v�!�� F�k��!=��$�+,�d��8-�u	�/uI�v��u�ge�~�Vz�.G�e�_�$�}�>�g�|��B>J���Ql���q�h�[��)��d|�����"�o�H�����+����__�!��qY����G���% ��� ���j���}=�������Jk�iY!�r���U"7<�%l��iM<D��|�[d�Ӥ,�T3q�G�;�L����?�2u����
%��/���y�@Bc,Q&�ٛ����?��%yA	���\(ܭ�Sế�n�h4ͥ���C*������p��	��j؎Ӿ�-�p�,��Ff��+viԙ(m��곓�)9���G����5���0r]!�,���0���`���f<Iac��-�C���>��[��t��;������V\9[�}\�/[���1H��M/�1ތVw����X �~|��<l�\09�,bl3��#��C�
�o"��Bt��<��ω g��̝���E8YL��	�c��c%���O�A�/0ˁ��5m��Z8C1-�|��a�4���(��>[��x^�z"M ���^��QEiJ���Ф\�6�6���w }ʎ/~���t�]4���M@V�9��tJ���^s�d#�h���ӝ�[M&���f�ʅ�E�{[2���,^龔���i?�1k�;GX%k�kM6ȶ}�n�E�G�l��PTk�m{lC 4��s郹C�d��Vn�_'0T~�^������F�L���ĻB�Z�jU� 5d����Aѐ��?+���irg�I&#�� =՘2_�����)�2�N�GL"ܞ��G��h��ow>�S��F��fk3ɩ�ݐ�|_�\�����/F@�HV�-�&� a�4��!0���r��mo�M���(F)�pu�h[~#���ظԮɞ��سjksr�6����.'s�!/\
�)[}^���r2����;�����%O��*���3�ktv 6�x3f ����/���x�0 �b�er2Q�����0[K�snA
�$��o4���7�%��3�p)ҿA�>ԫ�H��qޏ[:�fǴm����7���R/������;�����))4�?f�"
�6��&�dgy�-��*�i�'��D�]{*�bC���̹��:�[ t�,A[\x@ȝ�)ȇ�oP*՝�5�RIԟ�K���՛�.�n{'Mx��O�MI,k~�t4'��cR��[{��3�vx�-�n�m������F9�H�TîP�ql׵���G�R�-�D��e�X:S}�}�N���+"+�C�[mV��7]hn/错�ދ��O��5xC���ݰ4u���_g5�̺�������̻)<A����Ü���kN��M@Jo��W�S� N��5�ޣIW'�����96��e%P"��4��:,��� Nvu��pH��X�uW��i�E+)��� �?��np�����BI=��q��d<uQ�w��i52�<h��C�*�~Ǩ,�D��ރK[h{�5���Z,��4[]a��b��YM	
H����d�1�qFx�xڝ<PV��a���們�(Z�L�I1,|�5�YҴ{�Y֪7�;�������^u0��M���Ч�p��R��Y��"ɉ�}Α��t�,��&�N�WG�`; �M9�g�4~�����H���[�:��lͧ����< ]�{�d�]�������4Oə�?4��aw]��r�G�e;q�7��]�����_���h������+��m��������*�#��j��=&Ņ�WJ�ޯ��W�,��D�5^�͆9��uaL���lOTA�ˣ?ph�LK4��3�:�m�"s���և�#V���%x	U&O��ۥ .)�� YdS�T4C�	��d9Ka��E9E�-2Q�9���hZ�#kRgI�Ϣ�B���c5���p���t��׉h�[��bȩ�c1���jhl�q��8B"��Ѣf����㻃7��O���E�>�����~[�2��*�3}p� .T'�&�G
��^������.�����?���C��h����EFB���u�B�(��_��>��R:Ȏ���>ճ&��/�b,Q�Ll�����"�&\^ɛ	+�⊱w��V獔����u�1;-
jM#�ϝ��l�1}\0���p�3z��7��s_*b� �/���	:F��d?��}���w�d~��!t"¹�4�Lp�e���"}�>R�H�K5i��͘
H.�0n3GyR�SZ۸D��Fa�zr����_�<��*���-Ȭ��u�Z��VJ��0�������C���gk����S���`t���zգj$��}��g�~?�H��B��JV2q�g��ki���?	pNZ#u��scmL�G���q^�z�i���`�"�d�h�٭��0��'/&�V��20�[&�6Ň�R���)���2�Qĳ�ѧ���� U!9�c�+�+2+<��C50���LǺh�f��.{�]���*V�riz���J|I5S"Ӗ�Q�^b0�����\�0F4�L��P�닝�T�����jUmp+�|��7͵�����Y���̯�b�;�"\�(��Q95ma�6o��i��Q���!"%d�]��܁��a�.j�$f�AH��L�B��b9#��C^z�y��,�6�җ����<x�;U�uj�d| *��k��?��b�b����|�G�r#�pʉ��h�Jr�ll��������H!7K�Ԧ�s�OHB3~༎��C�>l]?y����P2��Cb��>Q�H�҂�O���Q�-��d�{#G�D�xL�f@ .�����S�0�G��egW�)qU�~�EXȸ`�O��U�TC:�n��̚���&}��pI�	��շuy����������3��b�TS3+YP�p4�؅m��������^*㍽���_�K��~�#-^�zLN�S��D�t�+/3+V��T�Ġ%�G*����,Ԃ����G݈[�;��hy)f9�}.ٵ�¾1z@�~v/���25��Q��Y��f�ŗ�ա�I����9�l� ��/�Yx`���@C�����u8�� ��U������ս�58Xj_S��(�buڽM|8+ܴo����~{R& ��{I�meһ��{��I��k�iW�l�@s̀����+��:��c�B���+���P�
�FN�a�Ԋ���1�F�{ ��'�T�h����T��;��M^�X���yw�v��]#�'!�^�غP�,��M�����>���"6�<��mm�x���� 9CC��0s�m��b���Y��r�q0` 4etװV����xTG��,��+�z���m�<E�N�X8�ٞ����e���^�x(a�<W��i�?k�_���sq�@t�$�՘�v)��+��q��$��@��O�.�d����:��,��=L��ưL�YR�;�jK��	�!��0���;���BaF}��vD���,x�>\�jlhN�3FC\ٟ��qc$�ZB�Tm7���w��s{-]���M멌Z;۟�?k��U���>>�T�:󀚯��'��ZȻ�є/v̬���c����lsn^�^M�T&/�|
 ��%�R������/[]�mB�ν>솗cn8�XQJ,U�.�}�f[;M&�	����!�.���2�F`�0��ޤA{��7�"L0�P�0X��]#8���3�z��9���p���0%k��s����,�͉l �Y��.���@�Bۜ1Cp�TwFc��}�e^�KN�����e,��vD�f��^�w�!(F%GT6m����]1{�p��w�{����P�؇:�3$�ʺ~2��9�r���gi��6�W����J�}����'R<V2\�|]���eǥ{�%���>L���A_UR�6�Z�C��h7X]�m��	���E���� �?(�?P�Nn<�+N/ņ��	��9]��S�t�o��'��}��H~�[ItT��xByK��J� (���/}.z�3�9Sˀ"�c��d�wL�]���3�UZ�|��|���,������uq����s��会�K�!?���_�(2�{s9������&N��U�S_g_a���&g���o����Ӝ�E�� (ä��vFQ�.ܕ�X���ع�vE�����PnuK-i�&�Η4���	~�n�1�$<�x|T���z��!���(�Ͼƞ���`��]��=p%t��uZ�'%A�h�"��v����Z
��
�%"��G�K���~>x��枛F�ipy�1Ű)_G^$�888L���b�s���BO��K���[����8+��� �ob��'\���)��Tֻ6�E���4)�{3�Kl�	�|0Y���[�f�]���lQ�І�l_iO��i(�Z;�Ac���o	���"�أ$ekB���<l@2��Z�K���{,&���yF�lv�4��
�b諸א��8���ĪU=e��]?Q�]Q.�b�*0`��2������UjTs�1�R2�"6v�X���zV�	O��k8*��w��w�B?�cX���m��ĉ��d���T�i�*�M:��q�?��C���9���Gx���l��=�F	��ն��)#��=�#�M���,gS� �*�8�opqn	�ù��)���ͦ�ԃdI�No��w/�!�]�v���b�`_�
�������`�PCͬ�^�u=�=ԍ���҈�l)�	���r���l~(�y"��ɧ��ѻ��y��4K-z����'�_�O���R�L8�+�p1Oƴb������o[F�ɦ)�C�ww�u����g�T��!�Lz��ʼ�����ˏ��(��֦7��J
�j�g����>��HO�K����<Oy{����8��Z7��|��A���[��>��,����n]����Ғ�\��<"�4�2�D�F>�,<�k������?���J�$^���k�ޅ�F�,�`��c���w��M�r]:⾙��0���FЮ���H�W�/	5ȒX�����0�֒z�i��*a�W��&�22�D��V�]��k��j߱xb(q�*��Q���b���!fw��̀}ߴN�����I�EC��>ė�:�ǯ~|���)`"���`�W�n�&��3XO��ݢg&�[�h%.��~�X��|�� �?�M�fw_�%��I�ժٚ[�9�ˌ�C�tD�ȫu������,Qwf:�%k�qu={��A���^�5L�<'Y*"�3�_�A$ �ņ�g'.��+��`a�,\�:[�Ќ��*UFWc�����σxui��be:���O����-/�� �veMaa$�N��u�4=��)T�8Ԅ��w̜Jo��<&���	�j�v#��h��b��Ǩ-�"z�������WIfq���>���Z&�*���J={�a#(Ǔ���_�W�炝c���oL��ve�F6�b�i�GZ��ۣ�+x���ϒ��p�#D�[�y:3_MHq���'ѧ�!ʖ�C�C���Oby��G�.��֛��عvr��F�������Y>�
&��hr0�Yh/���2�oL�n����B�0�яQ�~1��u� �?!5���
��!�-��-�����V�(k��I�[:g�~O+�<a1ɭ����Q��nK8��5Q�ӂ��ͼບ���,��3�8���	�L}��'
 �&(a}^�{
*&���(��f2�xFV'6M���t��-@��C/1�Xdw�p��a V�l@i�Q�)i�#X��u'������8rEw_��������3VH�M�qҒ' lOC�D���!�8S3�2�Uh��	0L��O�ܛ~p��I�+���8S�!5�=�}��!�޳1?^s�n_VB���π%r�<�����=9��чơVv^NaSiV)'͍�q��P���s|L�|�Rj�q�6�<��PK��E_�bZpb;���l���^���̄���϶��%["�}.ZiQfw������՞��<}�B���^�)T��J��?�+�����9}���ܥ;�Y̍�����V,��Q��Ól�2�����"���,<�K����k 71����� �Α�Hcs���~M۬���
�(���jx��k��n���'7�YS�G($��dKo�u$ĸ�������H��"���"Xi�|��X�e�)KuY#�j�!�����ՙ�掟�1����c����rQ���WɅ�d��6�2&th�8z=6�\��|��x�ڨ9�ǘ�A𙙾H�
�GDWK}hJO�u�"A	���n��X���oسF$�pqi�R�'��qQ5��ߞ�#�!$ػ��Y����*rY�e�*	��^e����/,*G���$�K����"�4�T�� ��b}m�㴉�{&M���	%N\���ob�ԁ��5Q�;��AJ��H��ٮ}�Wy�a����`w<���_��Ӎ��>� #�������
\`q$P�i�@:��F�)g�����x�&V���z�����/ ����+��de��pт���6�� �m�$��J��s?��o�X�ф������(�K|�;���18���R�`�ᶸ�@���Akh���d�dty1�"�N���Σ2q�_��8{��D.x0�"��O攋]�D��b���vΕ��O�$��ѿ8�MYk��X�-@	y��Ao4@�15*�����\��L
�2�oA:c���>��Ah� �J�/�&Ͳr�
��+�|���I�}Y<�1����A4���߳���5��CWг�<��pN
}eY���8�����1��Ħ<��͙�}���:�"Ti� )�L�a�����؉�'���+�8>F��x�|2���
�^�����q��fa��vn'�w��D2	���Pd��|��D~��?�R&;�X�o���3���NN���#E�f��3é`���q��$�;V��5�����8��z�^�=��/������ ��5�' Fm?��V@d��`Ϧ����^_gX�q?x$ ��k�XmT�A�1�V����y�X�R�u-�H���zV��l�z�}�bՠ���ͨ{��~xץ89�:ͦ���B#33bޝ�-9RB_�*�Ţz����%�K~���h^S,$��ÿ�^�*�3g�"G}�Z>��/�J�7:ӝ;U~�����j��u?��UGѱ
7���T�qx6��u��c����u^˧_I8��b�āp�T5h�i=0��]K~B�BTюkBsj��.(V��&�E��ک0�3=xj�	�����<����Ղu��K�Rл$(W���5ˏ��v��\o�v�o���HK��dHѴ-��$f�S8Q��l���u�ms�Yu�3Y"9�Lwx\�{	^��� *L�S�U>���p�Ĭo�Z�	lvLפ�so2��x��7ba���-h��O�ΙȠa�(>���MG��3Lo����`���_(}W�IS�캧����� �%',tA��]`��f���v��p&�o�L�3!�ib����y'�!�Ȼ�ص��"=��g7ĳ���qbV��D�{���ݛ��jR��	�0��Q@I6le^C��u�@ޑ�eQ�R�}���.{)�J��:����Д�)�B�o����:밂�)���d�`3+������(�u!��וr�N���E�f�!~o�\�X�`
2��ˎ�iM.H���?��gp%��rj��Ql��)�̴?�Z�Jy+4	pj�L�ON񧑀V�'�#���D�l�q#�=���Q�q��ۥ�+�������2K���{�����t�7!*�8�ʭ-�V�8t"y�A�Ұ~�"ȡJ�]�$���#�`�e>�XU٤.��4��)����|�n��V&�[W�ɻo�e���9�J�Syk0��ܦ�+�.�l︖�:�}]TUZثp��Y��F��FG�\h��9�K�����r�k��}o���ؚ�@��s�e�����t&��K���RA��� �.��2��a ��kݒ��A��;~�胶
`D`vȬ+^�tɔ���ګ��hl��6��l�zK8cľ��l �1K�X.S�z;�}�����	!P��K(�u�d�'f2b�}�h6{"3?m����Et�=������&��C���I�d� �6�R�O�*��G��7�5[&_�U�;�$��
��7�,�9J�%�������Z?�EwM���J(=r/aM�N���?֥x���gX�3���p&Z��i��yG�u8ĀL����w6Y7ߝp7G�y5�6l��
�</������ù�a��yKŰ�2�2��c@�?%�\�x����l��@�ihlV�r"�$�(��#���<=���++����y��j�k��\(F��p[.E�����,5���JK(-����]��;��k�?���p��(�`����/����#.��u7�r�&l���0�=^_���''��E�����3�p�o�Y
3���V� �����_Eރ�0�t��0�8|��ވ�;<g�٦Q���o�����~�Qt�"T��Gc�{7d�P�8?b�'*wrVD�/d�_����¢e��O�|&>��Ԕ$nu�L�Uȕ�/AF8q�r����ڲ��@�
p)|a���Q6�w����m�w�ۘ�w��!;y` 3�qsJP�	���`NfR�$U����xv�jQ�|
mr0�ȏ��C0��UWI�R{'�?P�z:U,qoq���ڢ������W��i��l�
RT��Ĉ��+n)�T|�=<|SZh�Ŵ/�?�p��?m�T�zZ7�Aa2�87bN֒:��؄�"N>u�R��@o��*>`(�V����J�D�4w�n�;3pC�}�K	T|�xr~B��6�U=0fQ�S����&��"u�O���n��R�h"�dY��������݊�0�17�;6ݕ�q�>8�}!�N�М�k�"Sf�}�5%f�t�#�O��0�:����>���ɜ(�wG9���(p�h��P�ɭ������/ܗa?$b�a�����3w�ѷ�y�Vx��

49�~d�¸�ED�T���om�.)����˲�1taL�c`����]ոD�?�}��,0�U�`I呂;m�c�A0@�