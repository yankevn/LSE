��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���}�C�s��9���1��	V&jCӒ�}�ȅ���^��7s#}+M��N0����JKq������E������n�=)��O�9!6�^,��}D h��+c��3�zχ+F&�jy��pЙ��%|�ԙL��V�A�mHO����_8/�B
�qBFԧ:����ͣUoY���\�zP��1}t����q�U��O|z�)'DLAh����ju+4��	Y1��[�Y�=rܒ+G���7f����Wf^e>խ���0ȅ~/~��d��ۀ���'��@1;�`�����~��XC)o�fU�
�-�ropO�%\RY κHe�==j������q��I�uɪ�&����0��s*�W�����[>*ӎ�؍)�x��&I�
�T��:qG�t��j�?^j%�x�J��l��?SPt��+�m0�%�*���|�%�_�~�:1���7z���z��V(	��:�L�<�ȅ3��w9p=�����ݜ9wA�?l�r��ڎ�p.>mBiY�1��R��)�x�����s��D7��"��·v�!/!Y�����n��S�jL��/יf-/HT�}���yj,Y�ۚ⾢XB��]:���]�b�����{փxHQ>u>ԕݕ����:wU	�@��OW~�s� b�vm�gH���e�"��Fɒ<�elD����l�h��^��x�J�L�mO�u�I�O��x�fC	h��$4���vx�Y���m��H��c��C7�|��*���o%d�L�ݢu��[��ZN��>s��#.�(>��~.\X��;�2��M�8�\��(�;ȸ�����G�����<c������'��\48��ź��تX򹄰z$���p�^ �m<)B/�}��3).�
r�L)�����ؽ��6Pg��h���^no�&I���V��)��J7C�Z�V�4����b��"�o��GI��'WF��M֟K�%�^�������Uٯ/�.����wi��}Jv�m x���������W�.��R������Ǣ�#����9%y�����_o�sL�.+��1��n;tY<{s�˟����`�{�UN�kv��7�<˥95s�k��Dv���fm 0�9/?o���="��/�3��'��Y����T��������G���3njb�qբ���*ԅ[�2M2� l�ro�{���/��&9hu�:����B�qU�:���PP'�/���-�ܴ�B�:��R\��
�T.�'k"�n�	�7�=f<�����~����u�m,P�!ʜ��n��x�����8��"�ȹ�s���&)�5c#���=R�,\�D"i�х�sQ0W����ׂc���,{���k�%�J�6�.y��x�4G�MR�'~��FY+? �Y-�Ś���^�)ٲ�c2�o�
Hm�\q�����Jy�c?萞D=P�'�1۽|�K��0e1���	lΗG[��u�[� 56��a	�U���a4�E�9E�����ͺ�t��9�D�����jen����H
b��Ɣ�mv<\}��`�>�<�p���D���q��^�JT�|Sq��u1�CҳפkT��Tl�r�֒M�\���ϢڴJ��!�*��"5f30�42�d��X��ĩ�N�ki���@���G/����p}�+�������Dۺ=�zm�&�k:����a�q�L������mK�⏓z	%�wY��!]�`ѢL���y�)�|Ͳ���G�Tr������)��Cwٟ>u�̲������Y;FQ=�'�����[�;�!1�^-��	sg�{�I��⩸��O֏���b���A�{�	�ʆ��W�^Լ��P{�F�1f,�<*2j���u�%mn�R�����t���f�S�O�`a��<?�%y4���@�P`-
`���fM봅.�+������C_da�L�vF�MO�=M��!��<�H|���c�,����<�Ws�_�a��ֵ��?�0�O/��,?}�1M�����j����2/�{��^�VϺ{��Ozz������[�W�	_�O����]�?
v��o�}�1t֩g_�u�`u��-͙��@T`�5I��=�|�_v�^Z��8�\����������s�5Z5���W	��y�D:,z�ɐ_b�UY���02��Ի�����8��2)
N���޼l,�N��w�<�55iR2Ѕw��'e�v��Exd��2I~��S|��A{!���g���޿�[�x��U�b�[<����~��l����,>�HI���>kIҩۃ	S,I��W�`�2r�m�,�"�s�P��M^RawE��3��N�6�x}M�Q�Fh�1�N~<۟���'�9�RA�\5���ͽ�HH��B��_������w�F�Cm|�4h ���n�R;�$j�VE&�F+A�T���3-]�8Z�Ve�O��V�D���
\K��A+�YQ�Z7�q%K��#!$�S�&���!yl�AU� Hƾ�5U��l1��T"�N�U���18�$�I�m��c��5�f�6Xffb�;�!�����wHC�gZ3��	��5ٞ0<�(�� S[�!w��Xn45�
wW ge8_� ���Q.Q�
u/ΰ�1����Cu�یUFQJ'���[�\�}o��w�� ���ɶ):7x�����EL�7�-
̳��,�学�2��jrK��cKǸ���k��B,vy�O��R(<mZn�[�<Z��U�@,�54�D(o��:��k�����V��i�C��L!݌X�ѩ�A�8�XA�aSc<�(֛ن�,n#Gq��@.eP�K����ʗ�$�. ���R���C���ӯW,4�T��8��q��a@J>���	��2�*L���ܗ�~���*)1ws]RG.i��s�-_�W򠭂���P}��y�&9�R�`�Y�o\ϼ����@|�nǳ���93��� 
?*3��z��!��X0&���TcE��g0%p�ofd�%N?�8pO��{����v�N+����`݉:q���B���ŝ�3�¹��Fm7���r��K}�k䃩���ޘ���tcZ�F��5l���H������ `�b`G�@�c׊e,��7����/lN��=h�˻p(3���f�M�g���JT"5�"���/T��h$ǋ�%������3�6������W�f���@�V�~�U���3�_��1Σ�¢�ʢm���8|�,a�� -S��Z;?b8Q��2#����d@���$���Ѣ�@z]~n���T�)g�|��4t����6E`��ɸ�#��of����1�[�����콼��k9�7��������b�}�6VU�X��Q⥄@&@y|�jT�=���*V$���y�F��(���mp��RI�%�)h�-�LQ���(�z0�;ھ���(u0�3�*�1�=K&v�x��2�7��;6��Mʳ�V��Ѽ\!�X�|�vjR�.&&9l�`�k�-�?f�>�ύ�������KS�1P�(���-姻�Hz\5Mtē�C��v���m�@t*�Ӱ�]�t��/�����]d�n�� ���x���@(��D,�pw�My}���r31�p`e��Wiw���Z���#d7Iu�Γ�ɴQ�iU�֏�N@��%z^
j��*�5*����؁�"4,���:�+}`C�.�ޙ������K^W
[���,�:�u�q�t��'Z{�]�.$���W�#���p��g1wbo�ZT��g��n2�ǩ��"ѣ�Z��Ϛ���oad��1e���¼Q�#dxd�~��ͅaOE�j�ɑB�fx�Z�0k�[bZ�\�v?��|钑���,m�� ��dc��Ӵ?/�����x]�=�����]�SD7:�N �M�OL,3����O}(��b�d��M#>]�����#'Op d0��M�lS�������9r|�=�R�%t����R�H�6�I昷������<c�i�K]�U�\H�������5�lX*�ig/B���.x��b��BO_�ޱ���������9[��g���������y�%��l-������%OU�bf�v�lle'EM��v1�l�^��F������Ѧ��kw��9e�}�������s�!n�'�Q�2ȫ�2 f�j�g2�]Z�+9��d:+p�{�p�lx�.4�q�߭�Ɂ�xMWO$����Ym�բs�����{��aZ'��\栔��x-�-\*�^wm�z�E�/;r�Ws� Q|&�t��r��lΓ�p���l*�AN����<�W�0~=Z �nI��
�����h"�6.�\�	��Ƈ���Ay�pd����H��!,��%e������5������	Z�vQ �?����&�ylc�h��?��u;�����_b�?�j���l��AϘ'�#����ǽ?���^sX.��JW$��&	����uZԌ�����8Z/��zo]}�/p�4�(?��`|ܪwV2��T��_�	�1�齔�JO��)�����:ڴ�`c{Af��
D�����C�Z��їC9�%�e��%'e#�Q�K����⚄�2aM�1�ڧT�K�8�o�,8��G�虉�����;�e�1�"�a�.���\QN5�ql��,=Җ�/��F�*H�	�6.3�/%�j����	�Ԁ�]��|������̡�\V�DY�*��18�� ���L��8S&�=c\]�"���[�~�!���_�M��P�jx�/����A�p������J] ��:�ȳ����
+�S�T�4u��r��)�5��m��~�g�Uy�gwk�D^.�]��X�4��ed��(���k��"':P�$ͰZ�n��D����:O+�j�f?��K$8P�"�y�߿0��0|X�̏kH��@�˓��ԩ��(Ѭ�f����N�ƌI���f9k���ݺ_?ɒ��d+�5���^��8��MzE���4Ƙ�*��$�D��/����]��"�a��]F����d�\+�oނ~��zi��&��P��_.���'vfn��vv�:�yͶ]�o����i��>�O;��ϦDMO*H���}%��{��3����m�Ѓ�A�Q-��xf��٬jD��r���<�5[QK��xy-����z�R7�'�I�a��-�����a����oÌ��PkLؽ\����ե]0h
�Y�t2{y"������80X������fP��x��b���-����m�F�����b���T���ª�iwFڋjBh��@<ԧTی�G�fm�7P���1#t���[��iV��=JJVe"�ό��(�,��zNL�"�!M�^����U/�AE9t:ʦ3E�i��0���T��z��� ���]ph���v�Rm�:�a�F�xlTjҥ�U
��"L���s��3�IZ�Em�������/��6\G���l�] �2H�/嫥N��<r{��I��`$/��6�>Н��¿��?q�!���6�R�̤]ތTp�pj�Ӏ��1����L�l0r�I�y.��e@ma�/�.?,S/�";Jk�s,�Q�JY��3��9�7��+�BY�-�I	��-�_�[��ĉ@X*��"�	���&R�zѤ �I�j� �T-}�e^ȇ,3� �����[ћ���5|Dk�T{y�l�3�t�lw[�/Z��8lv�CI����}jS��^DA��h���K)�_Y��]��0j�M����[ʐ�
���}���cw�e�N�'z��&S.[47�
e� [`(���^������:4��I���TVzܭ�Zgw	���M�OGQÝ��� �;����Y�3sq9j֒g�t��h�g����ߛs}��;/"r�{Œ�Y�%"y��V�)���n����gZ�����j�9<Kv���B{g��R�hU(t&,h�-��g������Yx��F����