��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~�����,So��un�w!��R�LQ���h�&]�\�Q��u�rF���P>� �����	=4�,Qn�r�p��u�rw?�-�+��'8;�V*Ƴ#�5}^��0b���G�1��P�fY�z/8"�3�����hp,7j�Ti�`�a�1�O��n0��ښ ;�i9�%!w�-g�(�_b~����g���b�r��?t�%Hɂ�?�J>S���0����?L��ϖ<Z���9)�	W{fW�9n�NA�K��B8�u����.��z�)Zi���ӳ	���,ۥ�-D�Ӑ�#J� %�s���M�����L�Ć���Q+x���Y�!C.�9�q��G4�=ڢ����NEj�Q�6��q��ߞ}/�|w(4�0C�E��ۑ�ν� �X*l���_�^D��O8�Gw%{�2����^횻��ds*~µzo���_Q�"q��*�
kR�M�^F�NI=F�D� �g�ꍀ/9X��Rɜ}�!��6o7�]!�8oBl$��arke$��Ö^y�܏-��������x=z���0�'4`\'���Z��g�m��|���ܓx��it~X�J� q.��}��6��V���0�����;WC��@�d��;�X�5����,�@g�
��&����KT�!�c�窇~�k�rg7�}��N��p
\t�<#c����Ŷ�X��0B�#v��>Z��k���M��d���g{�Ү�#U����Fx��ql�/����Y�g� �7�j)=��	m2���+P!^�(A^��G��g������w'T ��2��U��_�}c>h�G��u�v�r��Y˔Sce'^4
:dCX٤��Յ�K۬n74T�p���[��GF_�ӄ��fo������1���=�W��>%�Q���a��0D9"�N�����L��AO��gh,��<��Ӥ�сd���d!�%l~v���Ɂ�M�>�����Q&��y@�k�y�F�W"�W��3�Ύ8X�va$��c6g�#W
����yh+ѓ��X��p�	�cpN�w��Ê���0%��l����Z��c\�o��[��� �9��HV=aϯ��q�%���'����ߵb�-�}N�M?S�L;ȶX<��WǶ
���HkcE��K'X�N��q_�
/�ʔ�8�_X����o���!b�M��to&D|��1��6���̄��v��Ν
9_����`�X�Ob˫;>�>iY��fu�WٝjA��V�V�m��O�IG�9�Z��6-t��O�rT���DlԫB��'�_��yԘI�6M|�������L 9�D�����RSR��B�h����XF�ӵ(;k,?�2+��m6<I���(��f�����dD�'W�����U���V������!-�J����i�� Qx�Pք��q�����^��-t�*�t��i��#��Ɂ~���XS6=X��φ��K<�j+~�E��B5(��)�E�d{Qj6c,�D�l�.��p;��ooB%*�`�k�I17����ܖ��u�D}�ag<��S���\ ٫n{ AV�Y�%|����-�9�:����q[;��ڔ�~�o�g�i��P���?�-��T/AK>��y"�/��Ӣ��:��EݳވEj��y��6��~�z�`�v@�ƏFT%p�P	b��E��,�o��T�����9�)C���Ƃ��0�5=�Z��œ`Q|8H]��Vj���Հh���(��U�,%Ŵ�vty�Ί	5׽sì�����Yo� M'�&xd�j�.Hg�87��fW�&�VtȲ�vE�\�5�k��r�< \�K%r\�p��uJ�B��Ԣ:}aG��ua�f� ���D��|^���~L;�У&��N# ;�+Xto�B	Q�Tö�tx��v˲�G"���S?B���8�B)����V����\�������G��c�5^|,猩[&�4Q�I��7gF�[`>�ZqOU���'�<g������[]��R��[�R��'!�XS7�^��ͨG�E���Đ�p�m�o>`m���a�nsG�`y�鮒&��( ޖ��y�v��/G�8q�Mê�,��ܟ&IH��l��݇�ao1�bM��&~<Ʈ�\_C��B������>���J���t	6%��-/��D4�&�_�0�鞊	-�?�D�OB*�m惆��3qX��A�@~cJv��D!Ay:e�ap7�'�2��2D4���}?�o�^7�I�S/��={��d��H�2�`<#XK*~on��.$W}�g53�G��dG�����@|�����J��y��(j�$��C�y麊�s����KD���(}���8A��C�}�q"��wvj5j(���Qs[�(�FX-P���e�`[�y��^0s����b��*���@��ұ���zM(%��"��g�\2<��3������xٮ��gz��Bj�Y���w
\���~?���i�a�v9��3���Y��/9\.����O�μR�ua����j$�׆px���+�匸t<�%.T4g�*q�db`�PM�A�{ܖ�~$�,��c�$�'z�J�=���L���	�F��ƩLQ�A�E�ڌ����u5t�{8��ޒ��0ag%nIҪ��-����PC�	-������Z'�'�E��Fg1W�`�n��@tu���\�~������ȝR'�R���?P�ǮF�Ǖ�Y�C�6Q��9��G��K��1��/�6�����nǻ}:�)]s�W��7P"XCJ�T�	�>����{sU���E����[�RA��1 �6!~��%������G|.�S�w���?}����O�9�`g->���z���9�l5��㛶[<�� �0
$��3��ѭZ2J�-]-�H �#�# 8ؗ�KI^��2���������f�,�f�ǆ c'P����.q�B���C�*�'�Gj�f��x���/����
^�O�͡$��N��Dg@��eZH��v���FjFGY���_5muw�.��PK`�j�%���a�/
}��vA-�i��~��;,��D.bd����86���&��d����o�b_2�n���T�`L�!K���T=>���u~�C����>٣��Ԥ�53�.N�l�y4�Aўu�}����ɹim@u�Z�7�㙭�xF��:(>��~_���/(ȣ��j�㛶��.�T_�a\IMm`룴�,<����Zs2���2��Z*	�`�� y�}��\���ԁ��:}��1�*[��;*%��\  kq��bэ��!����A�͉ADs(X�Wy�2Kn�.Tg6��=B�2m��R����@)��0L�E�>]A���4��P���Ϊ���S��UW뚃�hL�ya[y������|�ς��&b6��&�@���6͏1m���:�<����˚82�ʛ8-�_g�!���һ�S]���P���xɺ"g���oINU|=y|̊`z-
Z�P3s�Zd.�6�w�fv1f��.�q�&��ꍐf�)D�х`1*DJ�0�llV�QT��|^V��T���'hPKq�H�� �J9����i��m��sgti-�\_
(��g�LM���J|�_�3Ū����F�`��_�),��q���L[��-���_�Gb�_1���?���+[��f|����ۥ��H戏�v���D�_�/�n�z��v&[�����9��c�$�#�^�����5�I� �C����_D�,WC�g�j��~�)z)(}�*:���H���^C�l4 "1 �D����#� J��EeE�MxO��c"�������;,��F�8�JI�*�2��s/Ҭg T����,�Y�9}t��?�k�p�g�6��j-��z���.)=��۶��LhDA@[���=��Z�?W�?��e_V&�r������|}!�$E�K���"�1�;h\=�[۴Ӽ�Yp����^���~	�]%���8�|�|}�D��c��m&���l�G��Y����35i}����S�1O���@�V\B��czܑ��b4[�mb����^��뾵<31�Vx��s韜2{�+/QmC�D֋�ɚ)���ˆ1�`kՉ�vq�j���ud�ܨB�|Z���Y�e�����׉Ѹwk�)���ЦX��'H�:Ya�\��7��c�>���pN�}��!���@	�D��1cR~_?���P��0ä���7s���^��~^3ђ��rjc�B�78�;nN`��,"�xsPN-��)��z&�!�"�	9�*��攧?H����"{P�E;��}���H����{+faޭ����~�s��u4>��PÊ��`���9E`'7M�A~�·=�!БH�_��g!"�}{�;y�=g�@�*��xE~Y�;L�;K����B�zk	!(Wz��lQ�Uś��0�$�~�:Q}�w�"���`V�п��4lc ���K4X���|,ėkߕ��I.^)щb5���Ȥ�_zm����=��/����I�h�Ma�&�;u|u��A�7�3��IC=��Qnv7�7Ŧ{������O���C�~e�۫\���w�]��PV��d�S�;��[��zhd������aC񵠛�l��=o��R�!���bԃ�-YL��
=�g�Dj+
&0%-@ᾥ�f���{��9�d�T[,�q3�<9F�\���}�ͯ`y�r�7�}�=�+)��ϛ�Y�n y$eO��2/<�p�Pr!�C(4�'!�;��U{t���7��`�&L�["'�G�����+�u�3w��� d��X�s�.խ�!�RNkӍkؑ���ި��VG�(��r��t�[��:-�Ҿ�M�R\.�C��ٻ0�����jwj+��Q�*u'�S�r鉶P�e&��|`�|ҝ�$2)��H��@=��G�{q�wє�P��;5��Q�#DB1�~��g�%��{����(ŀ�����d�]RW3h]���/T΍�W�TP��N���mGy�Qkj�b�z�[��XL�n����&���q��mG��J�Vy��Y�
��	j��5����y�o6� ڼ���'�G(:s��|CϜ�ɧ���pDb\���L�0A���[����?vg�t.3W�Ԙ��zOѤ��s�j�����8�U��K��:��8OOȿ���t�m�����81�NZ�äi�̈́����UNu/�@V�J!Q䋔:�Kpf�
�.bי�U�I�P���>H��2�mdH�E<hhsU�Z�)$�u4Ѩ�_ҹ0��|��A�O֩8���*��� ����]I$hrm��%)֐�q��{	b���f=	���?������3>:SV*��DY�PNg�?�՜ ,�ؽ�����ޡu�3��X�����.7J�"�%�cmޚ��Ţ�U�D��'D��w�3E_�Ȕq���I+2�:��|�ٱ`�e�.�Z�����(<T���<GX侦*���ޜKވ?���c�c_r�H,p����L���b�8z��H�~u��������Q!�kBԁ�*JS[t�Nx��S5�p�?��>�b�9�T`��$s���'=��LEY���,9��=!s�#�o�O?c�������va�V�
ȁgd^���������c�sW�n���R�������O�)&N��}��3��g�n��f@Ap�@�e�P�T~#$�F�W���O v��C�d�:&~f�l�i����߸���D���s�=o�Ɣ��:�0�S��^>�ʮ@G�	�܄��H����)�Ժ*��6������^|.nR॥����$_4[9������M��l��YK��X�k�C�R����M�g�b������yzu%�4t�sg���cf&���'�wgܿy9L�%0��ȩ`����ue\��C�˭��C�!+ٳ�?�2��a^Fg�mJ�\�I��ΈhH���f��J�bY�tߋ.��.D�׵��`|
;C��}?�$ʇ�*E�}��k��1���Pl�=y�]�
ڽ�!���_p$�a+��U��ۉ�3s�oK#S����g ^e�}�7��R�?�o���9���q7��������|�H����<�;�|(��W�( �����;�pj�?��c�)H�$�#q��M�m�cO\�97'L;�SFFp���烎�"�CF�[1b�ﹳ��ڣ��Y���C��䎭�P�t\$>���$��q� ��*�ݔ���d>�)2,�1%gk��!�p,�K���Շ��z(6�#��
�+��"V�:���d%�����6G	'�-8!�&�r�"��� ��J��j��8�y�j䤽��<��^o�4�]>�6C����7 ��GT���M����n5�ẹ2�����D�1��@.8>���U�<V�x����u�� T%���yiE���z�Eg���X��?7��,��_">�F��߯U����0�<���Kֈ��G�YQ![<e2M ��I��L� x�	}�㒓e�sa�OKoƒ�JcG�m�l`J��K�	�at��c�[��%h7,��~�X�M�x���k�1�fV@�8��@D�<����UG�f(ҍ��!�~{i��U��yI��2'�tL����A����Q��j�^����5�r
ֆ��0_�U��E��*/�C�]'��~�M��u�+��;L �S��1���`���:)N�<:υ/��Z~�D��@st���u{l#	+Bxt2��J��Q l'YN0��e4�kA�+l@���`����-z�����"�Z=}\���bz�_�ϧ@9�%�b�r
E�`��5�2���!!�¡ce��&�.×��%!o��%�ʥM=��o{y+�n%�X��՜a�?$G���o��U�p���W���{^�ҫ�(��%qcm�Z�/ۈ�O�'Hr�Zx�۠o
3���1��&j}� Gl	sմ����Y�ݣ�_��SC*�oMn�-�LipjѝH�:�� �p���Wk�����n��v��"1��/���;ҖSOsd��ȧd�H(�+�Ҡ�GE(�"Ɛ�W�W$Vh����R�K�x��XXڈjsO���Q��o���3�����`�GP5(��J�r/E8�]�~�;�C;Cf��I�7ᅡ�0�eYϋО��Y��q����_J�0D>Fa�@�K��'���g>��˥%~��D
��H�v:2n*�.X�A�T[�z�<1	��B�GV�Qu�̥o��D�o�UY8�[�;�,�Z:�Bڹ�_ְ4��iB2k�l�����x-�h��M��-=�lQA��g�!
}�M*��[���˃Gm�!�H��ZR+�wTOc#aP�m$�����}�?浵��J��p-O�SB�7=�StJ��[�^��)�8i�#��6=Sj�v��B���H؄�;�ֺ�?�'�G���j=��7�Y5l0C��㾻0�����4�g���MHe�wC1����ĕȌf踉����z��2�x��e����r'uS~���(g"e�!Z'b���6��|�1�,J:j�_����_zF���j���w�=XS�J&X_y�5B=?O��};�1o7�8�������4�NZ��b/�`�a�����$�T��H~2�0�]���s��-q,�Ԯ-I�*i?d��MJ�,�dt8nJ��v������'�M�CM�^zk��;m��aS���_�=�p��,��O�`�$�|��)�6�v~>� �L"3���rJG!�!�lxu�G�?V޷���@\Ǯ�2��ky��`�N�7_E{.��􏌎z����k?�0V�%��C��U3鬊�<G*��m��}��◈��\q�c�l���n���+��	d�R\��ɺq���cJΙ�L�_�����ʝ�u��D?���&b����v��wJ����laV��1��o&�����_�(���T� 31g����<�k�����za<�O�pgb��(�E�}��T��EاX��a����&��j���(�����#��я�����'ۦ6v߆�^�ި�b5,�DO�Z��tV����e�0��Bv�����>�&r����+ΰ �M3-$o��k�vQ�H���4�$���+�wL�3�2���T��<6^�c�^���`)s�d�����\�����t��O���p �<�
�ʷ�l!2�Ktp� l�C�;�6�V�s�N�ӳ3����� �U�H\*]͇-�gy����N�/��a���wo#եG�6P;�Yr�M�%�N��u�d��XԚ��²��1pۦ�
�U�uo�k�����:�����MN���8��>9P#̻���{$�;b)�0����N.�8e�+��^BM�QP�(�</~�as�~1hon��y߷!�4^׌R��bȴْh6��7����1'6&����@'-lH���D�)��D9�%<u�ķ�1��,ͅ�u����V���G�2w����v���#�Ӂ����5����y����M�����0�O=���|ӽ_�A�.��\/P0ު߃� TW�/�P��u�[�NaH��H�b�[��D�9�i=��!���h�Mfe�G��8um�ĝN���T�F��'�%���ݩ�]������TC3>���F�+罩@�ME�{�|��>
��nH�H��6����C�����<j,�
c3�iH��� �'g�x�X��E��Y��$�
6��2"�u⑓{�H��۔"�.=6(>9��([�6A�
�E}�tŘ/��(�k�U���Nq�Fq���J�H!�*�Np���r��]�Mi�c�c��c�{9������M����#>���J@�������)+�T��_����+Ȩ#i)�0dO�,�SR3e��M���n��F����Cc���q�o�f�����|�pA�lzQ}n�CI$e�>�XX�Su#(0�LM����Jk�h �i�� ؞w�G����������e�B��ڕ�oMcN�;;_;�2��I`T}k$6��`m"�,����vV4�N�\��Ka;��{)\���m9/��|��a�!�(�x�H��Z~����3qd3��[���.���]yFJ@���-�T�֭�8�0�3�c]b��������|�o�U����J�J_s�5Z7�x������>�UD�@�|E#Y�Y����^M�� `+��Q�;�d��<��He'��	�����;ݵ]�sl�1�39A���z���3K�a�tJ�@�pL��M�qR�*��C�Q�/�a`��x�N��6Qde�(�fc&�W����c<�D+�v������xO���7�:��2��?�W�ٗ��M�1���qFU�tO��&�M�\�)��p9=c�'��1�!$t���q�I��,T�.����#n}�5�,�K+Re����FD�J�%C&����L@�E:k%~����Z����R�_�j��/"���l���9��� �b
����7?4%��8�#�_C<8�j6os��S�'����p�Bos�*��b�����	l笠;�>�i�}9j��~��0�`e�*��[���b�ۍ���>��+��Wb%=�f��3����h�*�23WYB;~����U��ȑ�iPȓI�1�lr���ޛR"�o{<D��2���o����6ۈ�؛\>f{�i#1[򜹥��qX����Lȵ�G�y�[٪}�X��v.����T��4�ڀ)�܏r�n��1�ck��܏Z>��x�HV!���V[��X�4!��j�mV.�/�FVa��5@G�d�\NqE��f�����|YRM�M��릾h�@S܇�R-@O��W_X��vT�[x�~c���fJ 8 7�>"�]loY���P`����#��s�U����y~U��:7�QQ		����W�ٲ��<����>��%䭥a�3`y(լ����FS¬D�V�$ͥ�`��O�����M>_{��͖d$�q��(����0��Z�HK,�.s<qϻ:��^GI��62�vK��p�ȧ�|�˫^����9_�z�k
�13�0���1*^6^(��h�Kç�߼�B�|5ҍ�Cd�Wz@��@�Le�*yC//�e\��@��Qx$�h�Wî�lL��5*:9���G��[�A���^p
�*1Io�,T˿��~E�y��t��k��GD��7�v������J�i��Qq0��5����S��u|�ή~�����aE�@�v�ļ~�c�Ô�X���s$Cu;Vh���M����׽j{r��>_�d�s���Sl�s��ک|��F�s�(֘�>��ag�7N����O{Z�u�=�#��|�I��f���r�j���r!@��,/G%�#@nT���9���9���e�:���B#�ؿ|\mU�xY��%�����f��s]۷4sILx��N���0�f��ߖ�����]d���� U�^��n�1Ȍ���R�B����V��x�E(O�/ł�HTw��.�rHP[�o�
�V�A���ķk�`�Ӷdh��k�gưs�ʁ���ƽE$��z-���Py��\A�{<0��뱇�/�����s��� 4�_ArZ\Γ��@m}������P�KT(�KI���4~�k5�y��r4sz���R%h.��"P��ђ$�����_���ğ���iOs[.��J�đ�D��4}���x�&�;���]\L΂�v��yZ?��2R��LL��T5���{�?f����p�=�~1��淳��#��L3�.Mv�n�>�r.���w1S��3��� G����~훞Z�n��|�E��;^o�j���3��}{�W#X����J9�H���pqN2ߨ�a ٖ�Hx�m����y��p����j}O��m��G�tU4�*��	��v]��1(�ڌo���	�]9�>�8��|��b�aL>o��ɢ�%4�Θk_Ӯ��`V]IV��d�)��B�)��EFM�h���<k���vhQ��v��[߾��i)�[|Si�r��]t���I�͢F��0��5�x�k�T_����o3#���wH�8�.��L�ld��y�U�=Dsf�lYY��\X;w���H�!z�7�or�?�c���x8����AԖ�vj��+g<*v���+����_#]�`���-��/��v�1%œ�C��Uc������5F��@� �kw/��l1��$��:J�\�@bxƸD�q<�S�{kA�(.oU�E�u ����X,������	��@���}�+�>��3�o ĕ͓~��I�Z�kcH��I�A�
pU��>A��d�z�����	��# ���6f ��]�đ�弈�6��>��#P�D�bΌ�(܁P8�ts�>J�HJa�H��co^>jkYа���հMu��&�K�F6^��9��	�N�L.u�1"e�8<�}o%}��IR������_����w��o����!$CY'R�ėv���h5�4T��F�`'�ChHӀ���vpd}y�wiӻ.��{�*���p����=z����u��šX�ң��縎��h3���u	]g>��H�"���1�uXo��4<�2j��[n�����ο����Y]�㽸��=c��̴�\����t�O�@��u5M�*��iƓa\�q�\�H�{��?��)�0P=�z�1l�ZEq���c��V)��#�>��<�7&���fQ6�E��*��W�V�q[ی��A�,
�Wʕ-�t�ݕm$K��ڌ���(��>��~���(������m�E���U7���0v���[�]��'@o��s.+,-!XP���F�]�9���f�8��E#����m�BE~l��@��I1Ml��"�[�lk�N��/�0���<�Bp�z!1?�އYo'���-�, ��>]��?6O�/+1�B�Jaά�$(á����8�x��]:�{���V�K�<g�w�&y����j���8�#s�ܽK��$��e��`
c��F|���Ye{;$������ ����ˬB��aY!�Ĩ�� ��\FǢ	�3���0u1�]\�az.֐�#�{K���ܯ�c��ט���Ĩ�w]h��^֖�ĨM���y���L��-#�8��y�*�`]/�/��Ցc/]�	--GZȎ��P;[�����f��i �lː�Ư7j8����?���`?\ ��O����x�z�1� Y"�J1A�yL�ZXaZQ+e�l��8bNg���<�#�v_B5�� �p�10����lW)K$W�
��| "�� ����]�j��۾��t�p%x��|������p�m0ﱳ<4�$�X�Ʌ$�5p�%������N�[lܽh%!��RnO���;���n_<p ��C[�H��sE!zJL�
G�/)����|�i�@/�,��Y
V�e��lG֟���(�������ݝ��l��P�|}謺�ұ��{��d'�+�,����9������ΓnF�t��
�ܑZ�f�ݷ��0�QCU�'�o�����˙ �j�R��E��9�j��s�u!e�BFْD���c`�w�3�%��miz�aM��M��6dǹ�;/�9*�J&��B�m�4�#��H��?J�a��"��8��=j�9���J�Mr�}'��81.�إ���G�� ''����C�n$C z<���u�#?ŭ���@~'������q��|M�Q~�9q��j�΃����X�� �&�r����}���'�ꉇL�*�v����(#Mա��
ޔ��Ibjy{5`��K���I\�8i_�U
��k���C�O�L�Y`,� im�=K&���y�93��ٳ�'��ݦ@�?S ���fd?�����,#�A�u����p�q^T�)r���r��a[�s.7H�ݸ��TJ��C���u�eX�/�l��'ז��2��;�K�o�xt��;�O\P�≳�/ߠ�TO�E����4�R>�u�Lvh����," ��G��}�l3*�a�K`\(ض+= ��+�'��;V��,H�AK��D"l���O�����˫V���]t������	"���๊�ZJulb�Y����O�:m�7����]�oD6��;��wP�Y+������>JB�cκ��z���fl������[�xI�x&|\�������?���D�_�r�s0�ai���a�Ì#ү.U>T�p���JT�@��ZU�-p�����Y+;(��r6�FZa�4��X�q�(l���K���`�YȻ�f��{�t��֑�4��U���f�������S9��hA�;�ݸ���j���]�|�D�Z�22F��J�k�G����l�����ż<Z����̀�ЕK*���K�:/I���(�i���?&�hو0����9Rc���Չ�|*I*v��i	X2b�-��(:i��m3�4�}�<Uc�4t0��U�PH��E���C���V��@a��-�ac6ݚwµ�dQrz�F*�6����M$r{#̡w�c.*~m�%���(����-��۫4���e�&�g�ǚ�����_3Ao�xI�b�7�S�(L�r��1�|�VU4,~�{	W�N�ê鼻(��"y&r�,�{��,@thVZ-��R�q�V�\��+ݎL��4q��s��ٌ��,9A�5���'4+{}_k�S��v.���,(	����LAv�j50!�>6�5m���$��b���ە�/�Euʡ9���rG�D���i��Qé"�j���A.��3�v.��߆���
��Ȍ�7��)�8c�Z�
��Z��������{��%C֎���w��	 5�&�#��B����AU��l��6�kB�wx��ZO;�q��Zk� �??�OU�w�+�˺`����M�����mӾ��m,��ۅ�Xɳ�F'ѓ@�8O��`]���sկ1��γL��҂��@��c,�k���^
O�����E!P�<(x�)8G7����z;:�Nj�����H0�a ��]?�M��KmY��{F�%�7b�~T�\�=6�BJ�K(k�E>������|�����,4
�WqI��Z�	��E���S��6c�
˾�7X���������E�t-��Z�!z�ʄ��%Dё�����OԼy���R[���ŕ�9�O�">�o���V���6�ֈ��?Sk�ɉ��l��\�4���2f�\P��O�Ϝ@��0�
�3)/�*+�f�bgJ�7Jy��Í�	�ɿ?N��R�I��P�[h��1���-�ˬv1��BJ�c'��.�.?��w�So�/��D��=G�;��D��	���*D��I;��]�r�Y��&��TV��M�Qd�Z��������y���1 u0�u�7[#eP�a�4�6�(@�O��Z�ș<��EVu���~����Rŷ�Y،����x�����5/@ʹ���'�����y�c*�e���"����3	O�H���-�w]��Y�x�3pPS]�q�""bH�R��s�^�;���y�N��� �BI�@�Npf��7�N����E�9�8]����u�o*�%!�@_���ր�AE���[�x���)O�J���1�q�؇�� B���be��6�hb7t��z/�D�u���1�C��Խx!���� ˌ��T]����U�9 䢔㎠�;o��ܷ�=�ٴ"�O��E��.�5�}5�f��SG�&佹{�(7�!���Č����!_�@żr�Y�>�ٳ��_I3Ȁ�U����X�cp�Y�,� ���U�p	���~����li�CqĢ�Țg)�Z�. <G�̿����F��,�'�9D���*����5�?g�ޱ7��8ś�I���3s�Nb~|��#b�w'?�f�_���M�}@�J�l��b�����[^����`�.��.Ր�2���������r���G�Z��K��ƕԕ�&��Bv�mCIra�oR��3��z��U�ICR�L&������/[k�J��	��>0X̕ѽ�v�=� i@z�fϝe��zm��,����#�0�s�۴Lz�:e�YK1�῍a�9w_�NA1C�������X�/9�.o5a����#���P����#��I���"B	�r�˯Z�1�����{&ޢ_�Z۹�Y/�
�6R�t��.
+̊��-1z�۫�u�c�4Ħn�ʾ��:��J�92��߻�C�qݣ&�f	ჴ�N�jS���|�(㖰����@6��3K��kF�+ډ�I)u�MO" k�AHq�4_c�]��}翯��N��� I����A�n�q���j��Ѷ���ds ��
�����>�+L4/������5��S���X>��<���B��w�9+J|6���Et�ᙡ}�#�t�}ʎ�]?����avq�G�j͢X�A���+� ���r�>+nJ�5�c®�$�.d���Zgn����G?μ}��=R�[\�ҩ�L:?L���] �xk���1�8��9�φ�����n&�pv���0Ȁ���ˇk|>f��籖gLy����sZ1�� �44����Qµ��²�7�))Oi6U�.��
�'�a^2+ ���uWP_�UzZz�8��v��gLbJ��{$-�a�+w0x���*R�9Xꉡ+툩��Ņt��jO"H��f@R���h�]FbMOtk/�����x�7<Q�D��z��A�G2�k��ż]���J��Ӣ�z8,�歹tA���!�LZ�m=� ]m�'�L�]Ƃ�E�·�"o��w���p�Ղ���Ma��˞W���i^Su�M�J��d�d�ɣs:txQN�v�l~:(L%^���b�QQ����ϖ
8��v[`ǂǑ�|&��'�i�%�� ZM���n0���yp1�����$di3f.�M�U[�em�+�sM�3o��&��������f̒2D�X�ԃ�[8�U.��o
�M꿀8,,л��i����3z�t�������"#�t{0��Q-�B���������ge�E���X}-���֡���;��)!{`dgm��6�j�� R�c��J�����7P	ś���=e�D��E�x��O���w��!m�:�\un5�x���9�wN�f����Dh��,����*�?H����\�G�s(#�'�*m�ڢz��6���u>����C��ǻT��F��`D2��9��v�y��n���P�n�fcf"ich��(�0вu{D���ҝCN��T�w2�Y��s����[�6�so�sGU+��
�!/���&S�2�r��^�e�&���Aq?�|&�RM�sj�p?Վ�����{���K�u���1TEX�A9��cd��ԅP��j#��UD���s�$큌��
;Z���0Wu&�ϣ���gdO]������g��7�vMm��v��Z�t�Po����ȟr�,�i_�������O��
t���T��"���t&�G�E�����M�ǖ�c��,<p7�o���8�q
g~��|7X��J�ՕƁś�^Wtg���(]W-��
�����0�.+|��2��9��o��!�Y���~2F�7��!��՘D���_�ûq«���ΰ@by����A��l�k��i� ��,�{#x�e�̪�K����,�b�Zr�vA�b⡽�>J]��U����Ie��8�~YHBVi�DT{��0���)�>�c��1:�?���m���`pzXݻ�A�C�)���8'�R���9���m�/R��_Si	�����l�H�����[�Gvɔ5��y�o5"����|��|���f/71��2���!�S�	�N×��c���P�$����������)����f��F$^]﹨�ߓ~�����F�)j�r��G�A�'(Z@j��:f����Y	��A���.�Hɹ�g���J�ݐb��t���	m�����d�]�(iUW��w�H�""�P�ҹ70��~/���K��8 ��f9Y�`y�䜁vO[A�j�zIk5����Ao��ɶ�*�X^��h�C S�9[$T�xy�{r��mbs���;��Jk����&�&�lw��.�� g-E��r�(�_WՒ�.<)M[m������%�A�kf-ٖ�����Ҙ�b�)ˊ�G��R�:h��9$}xS2X��t�{F�z�H�vMն�P��w39�L&�YY��_�J����4�j=ˆ5��v�������
��[��j�4EJ��8Ƹ�����yV^��3�I�2�5[V����4*-;�(����|׺E��&��,����}���SG4�m�ޑ��2�R��L�H�F���!��
�Ya���Y�������o��;��ӧ\2Ʃ�����4,��A�%�]e���%.��>��n�Q��.����S��B7T�Deԅ��kz�h��͸y�6�
���f!!���G�+�;��&���(��"=�.��	�m����տ.�R�X12V��m�4�\�	WsC�wd����9�-z������i�7|�0vi�
lҶ�8�=�kzN �}X9�w���~��D-�L�>�U��`g���?�8v�b�8�Zz��W���+�ư��2M]�5���@����<�_��cz�_��ެ�O�ߢә�7c�"�F"�j�@�Ȗ�f.�T~������H�D_h���`Sh�rU ,J�Y	�����$U�Ǧ�̈s���o���HBe����/72�0t��L���!�����[�-�y��qD[R[8s{�?	���)^���u�Ɂ2:����%?���d�d7Q?��ȺF��JkU��SѤ2�C��4&I"���_s����j	a������*��Y}�V~{��#���D	�)����s;�Ԩ���KV���`q��#Syi�_F������ݫ|��$�7|[���%��K�W����h�Ef��嗂k,&�;�[%��ާ`�ϺX� �����cJg��NX����0B��q������
���H���c�����Ծ?0.�s�35g��.l���ce�����JŞ�4�K|y��j��2�c~���`-bX)�	
\�>�(	v�����24}uueH�I��Pc��,?��p���.W����߷$�kKف��\���ߪ�@r������c=}ޝ�4�JF'D Ke��#�|)��~��y�~�d�U��~�J��|i�=~Ɇ�2�����A�j�p1�/>i��P�Q!3,M�n�)�ě�evұ�7���8Cc�}ۡ�$��t����_�F��ρ�t����!�M�?
g��X'��i5~8X��,�U�CҲqL�&���7�F���4����4H�x���������Ȟ���Y�K�l]�w�/���Q�s�>W��0��'�����W3�P�Y��w��t����ċ��N��ѷ|ϱ88��o�,~��i���}���L��C
�D�^g�Y����6c3+���.���N!�w	�&��M�	}��?@���t��pr�KE+�����W�QO(�FR+;�Qq:�<��f�޵�ʽ�g��V���}�CK����~��n��a8��{�m�pՆ2&oZќ��]���ʉ�:�|�:-�hop��|���m �iW���%Y�	�����ڟ�ƜQ�˺�z!s�VG(bܤ��V��������Q1k�����q!�;��\��Y2'Q�`>�m�a�W��,���8�����ԍ�N)���m�8x'P��� !���c�
bNN�=ʥ��.���~�g��!�L8Ӱl�ah�q�����i�T2w���喙8��&���[�\��T��"���w}������aL��u3Q^Y�f|L9fMsr�OL��M:5M����z؄�@���mÄ"#꫄S3M�?�-���-�����[�����>�	�Q��<2�T���^%�a)�����O�^"������`�,
"����gz�b_z��f+U\__?�(1T��rD�郣�H�ѕm��᛿C����o@~���:d�X&��J$�*���l���+������ߢ�&���u7�YF����a;肋�!XI��4{�fg��	�~�����D0�GA��ߕ�]*t����ç��>E.T�Z��ô2�p&����Z@}=�`���>I�lZ@�S���6=��Q��)�/j���0��D�	.�i��8]��J
�(��ih8x�=�`�}"�tv��0!����4b��%z)�d
�m�$�޳x�����uR1�V(Qmv�b�+���4+�.APn6'>�pAU+�<�Ŝڗ���4i���(_��EݾGX��<��?I�I����-B��Q�6FV��n��պ:�p%�n�te�(`���0���n��]�E'�<z:w��D��a��DO��)��	�.�륤�7q܅��~��D�o ��k�-�%Z���-� �)�,h�>�0�V(ܷ}��鯑�}�G�Yx��$U�[�e�(~?�r�`�P��Bb�0li8�'�L2��t<XJ|;ݖ��E���\ �l
���8��,iȨ��g��ŵB5�_�.�y~ irS^�D�B��L���@o\f��apŰL���9�>qN���Z�@\,iD~wC-����3SW�b��&Jr��M�B�>cὡd��#e�����q(?�^(q�_Sb#�o��&VK�ſ�b a�rу�o��ךkuA:X���LŠ�ֺkG��9a�$�2�&�!���pK������|�w���MG�����̿��)/��I�9qM`Sz�UhN�yC���^��S�te$ʒ7C��ܣN3U<c?'�Dh���pEU����z _�등�0'Z�V_��A�Mm5�_�[�.��<���l�i�zQF�b�Q}a���׺����=�Za�	ҩ0|'�GOs]q���@�B\����^3���d�D$�!�h!���H���OP���\�u�bq�x[��В}E��R��_҃�~���_�.O�gcf���,E[�]�
��d�TO�Z��uY��e�vɗ�J.��!�J \	ԋ-�����m�U��}E7� ��M�*��q)�n�*�����J�`^j[9��}�2�8�5=�(��:�JV�^�(��㈂�N@���>]
s���u�F�7��g�����M
�{GԆ�>jя0��.�h.��<J����y����o&�^�2G<"Q�!�����nH�&EO��ۥ�1c������c�(��<���\9+�q��F$�cD*qܰP�T��� n��x��T-�3+��������ɕ ��v���Οu�Ix��l���>*Y��UbY�f?���[w��������u!�~v�����ѣp�Zoo�֓�b���	�ȱ?�C��5!�yD�2g��q�7�!�{�4x�3:����D*��Gm�T�N�:KCGu�sal+N�Pg��m���	�Sk �����᠖��a�q=�����f�v7e������<�Ic��=R��+����OH`Ë҃r"��˵{�ڝ�	8�m��H=D��UΎ�8b����QD^����ڮ���{>(�=6��-��l ��j��*z�a`��qSW��>,��*����f���rɆ�S_�5�T�Bf�PV3(b߂ �Q�
�M�zp7&�-�(���H�~��\�6�)T�e�\�.)^�J���l�#0E8���`�y�ӏ`���S�֘�̸��$y��"(:�2�����jK���"��A����y��%��k �D�~.��T�v�����~RnxQ~��aqH��1���e��_��<4��O���ň���������x�A�g��
j����%=��&�7��+V����D,J1'���%�sB7�
Q���B��o�1e��Fİ/���@V��	_�F�N�h�FF�̓��^|�B+Ghf�aH����3�HJ�R����X���Q��T�*I�ѹ���� ����i53�"H`�K8�g�-ZnB>5(���,�9��.!cz�4���w|4�`Y�`w�m�/
|�)H���O%z�8���¦��ꇒ�=ip��yT
��!l>u}�
�ݢ��^/�y��|��������7�������{e���>��C�-�f��T�X�%��X>�*�C�F��A�� ��5��%mH����+bo/-Y:V�����h�I�(�y�}�F/߁��]6C�����nn��������v�%�4��ss ��	ٴ�q���C�ꃻ��,��d��J��ԉ��" �)���2 �z����m�s��w$L�l�U	�!w1q�-&�A'�q�Tl��}���#��?���9 N�7�lϽ�(���S{J�Z�ٿ��Da�@nl?%�/u���ķ���m1gf~�fh��\=\�_l�}�F���;W�>*��J�ڠ�o`�3�]�a�5f��iFW�5����|���$��D��Y�}���|�`FR���<A���
R�l7(*��c)�0}��3�d�P���c;N��Os������$c8��T_��-.��$�gb�)�d��#2<ƍ����ʧ��qU��>H4n|�qZ������?R���hY��N��1X̓`�-��^꿳_�<]����T�� �Ԃ����������P�� � !P�;p�f �-Md��b'p�E������Lb>d�����hat�̴��v�Fh��m~�X?2Q"��g���&�-�9'�k��xoM;��Y�sH��̂ت�eM�gk{��	�����n"�0�W	.�q?#���U��,�[�>mt��&�ᜟ����3�A�s^���)�.N�-���}����>���$,����f$���J��(c��2�ɐ=�����	Y�Af�W�鑮���V���y�e�Uď
'����c�K ��M�}4RM6i)BR%z���B���r��>����.���Z�,'�~�=7�uz�q��t1_�0�I�iY�ï��Z�9	��+�l��Dm$I[��Z��άp�q�N�ZWX��)��R_# &DDj,�'B�wU��!����-t8�D��p���#��v5H��*����� �$�<ij�@�F�x��j�.5n����_7���F���]�.�
P5Z,��������uBϤ>A�nX������y�����:?UP[q���9��O����Nl�&)��6��玈�	����2���.�o���6�ʨpV�i)�fl>:T��R*v�m��0/дZ�Q���8�J/�F&"5�i.c1�`A����}���@�#jX�xڃ)Q6�A�_��Ȣ���|�u�<navɥZ��T*����5�;BT6��~�*mׁT�a�n�I�|x��`��L8>Іܟ�O�ɫ��B���
�l
;d�d�n��H���+�:2ԶJ8�E��V*wz�`.XL�6<3�U�'RL�$Ep�����Qꧼ�_��	A�&/0[�n��
a	na�3��>�;��*�T"�vA1��68;���A�0��NS*v4}`����M�m�=.�>J��wv7	~?������KS�[����WR䗔�7�7�1��C�X�WE��݅�R�m��Yj��.��O}�=�.y�F*�3��p^b/7��hR'jlJ9�
�5@��˭/*�G@$�(<:�q�&4B[	�`�l����'���R�#p0<��
Mqt�e^`伅ihx׮E�t̷HQ� P��G���~��O���>@�p����<�j&|�KW�Aϗ����#�/e�B7j�_W4n�MH��O��}æ&n��Ԛ�B���l��5�4�$��H�I|����H�vODrc�9��n��DaWς�!,�J�W`�s{�nrf��4�&VY_9n��?kz�'u�N������=�J�i�������E?H���<p�y�{�Ԝ}�1X␎���F�Dld�����^�2�d]kP��kë�Z�t�jTG��0�H�������!ef]����Z5�ؾ���=�r��b_�F�M�����{����������Վ����9�������֓/d���݌�Y0�x���~qJ��s��y�5�Ha���	J}�8�|����!���D&~Wk�l�z��]ة����-L9$-���f����(�3��w�ոi�]4'�'x��Ű�������k.咂�h��:�_[�z���;�h
sA���҇}5��K�ZH���$p��sL]����U��'�8��ciV�A�٧x����3�^�9h��p�10�\Oq�p�,+�L�E.9 �2�/����T��t��׮(�3� �<�w�b���o�����p�����P�S H<��jV��LTW�q4��v�cm�M�y���ͅ�~��X6���x���%�<���.z&)[[is�>C���->:����`��j��F�Pf�d�fJҮ� ��6X����=M����p�t�Ţm�}���ە�-U���n�dƘ�?�MN�4�Uݡ~�*B�[Q�ݰ��'�ǡ1���;�J�&ݼ� � (1�{��:�ߝߟ��շ	)Fb�]��_����Y=u�10���|��c)��97�ؙu�7�!�S����d�!�y"�����jD+h:peu��"k���$1/�-'t�*B}� �P���go���ŕs�p[�{s�A9d�`��\�a]Lf�����6����:!tlv����MW�D ��A�su�"��^SZ3Eڭo÷���qӚ%k���(�z�U��	Ek��TWh�}�?½��%��X��֘0�@�_����6}��	#U����JA'�.t�dck��_��I�� MW�`/k谁�[��4��Q>��,�x�b�V^\��4���3�a?T0��xE:ǽ���R+�ٔ�g��֙^�e�ء�I�Ľ֧����#���n-�v+���Y#hl8f�4�H�R�����<#�=\Y:����9�lk��6Q@��dLob��s�Zp1��B:*�v�8���?���,�6�J!`|��KZ��
c�������@�L�NR��E�׎K���m��)���W暈�R�b�#��iu�'M؞�</�d�{�����\ktx8��snLE����ו`6�~���^q�Vk2�[F��� j���6�>��;)`to<���.��NR|�Y,i�;����3'"�*2x$��RQ�.�&�ԙcaZOU�|��?�V@m�q*�crpE����*�cS��E5���B|u�b$_�g���Br(X�FI�t�"x1E`T4!"y��V����L����#���[���)�	�T�G���gX���ꍆZ�d��=��/r�a���Y'@�gx�o1Qԧ�vZ𪄎��0�s����"4�W:O�#2$��~�q�ˤh̼����(�
|2�X�8��W}fK��� !�1�e.ab6p臔�j�Z|��
��N�_�9�h�~F�=��c΀-�	���.Q�� ��y��L��Oo�:5Z}�M��q���W��{��m��e.iӑ��w���8U%s��L�#!X�8��b�����t�
I�&���v�J�ƭ)=O������������~�y��t7���^ZdEr=��ϑ����}�[Iz�{e/=����"b��:��ef+A�2è����F־��������S��G@Tʒ�+%�k���+ĢIі�*ن.#���P��E[GZ��u%�q����c �~	I6j���k�q�3@>D<��(�\�@���c���"a�'%��ٛ�we��L{���d�
>�A�(�f���k��<o	��)ωz�I�P+�:����t��w�}��B��w:�?̓�٪3��V�\:7.��(�p�����Yf��\[D yhL�TZVi��ll6�2)��|�x}X֐��r��9DR�ƜV�����Δ�������Rd^Jk�<>N4�"&��VH���q�����Ν�@h���Ved&��O�/K�^L>S+2%��ಞHb�[�	�
p.�d�-�����G��X"���hD�?�QaҚ�B�zq��7�T\��]�s (0pe���M�<��2/��=� ��Pe�(���������p+�̤&,�-,2�Z���ˍ��>�8�
�`]6f"9�阎�e]��b�Q�HF$a�D̟.�\3�9H�����OŚ��5����d���m�����4ƪ���;U�cs�]p�f9�Ȥ
�F |Η�Z7� /�kQZ�"Z��߿�}��R|����Х(/`v=��2kB<����$�!�3��kR������!�ܒ� f�-K�F�:�}�3���Ds�V�H���*A��g���Ӯ7�*�'y�(|Q�ۖ��^&k��Dl���ĠN��.(H��^��]�Fn)D�@��O��l��ᣝ�8+��S����C��NY����ʐ"r��V�S'���s��aJ@ƏWa9�#뼇rSlE�a`J)hmq������|��A-bH����3���ٴH��I���Y-=L�⌤ig�?DHTԮ�	������_�%�@g���	�`��Iےg�z˜��5������P�K��Qu��ݜ�XN<m�Y^'Y[]�+}��J��#��$�5+�΀��[G�8��U���i�ka �iX�i�iKq�2��0��_�B|[9����k�����/�1��_�i!V��~ �
1��\?S� /���Y��JZ�!�=�ǽf��@����ȓ܈r�:{��4��*�ǁ�{���0��hFGr�>�x�7[x����N��&	o�U�Rd�F��m�A����{�2��լ�;���ZD;��GF0 :lǢkT�ε'EɊ���.XI��!��P�$�����K�ͪ�?=l�|�����)���q�wo2�����_�@��\7^�Q&6Ƅ����EK�t��wٓ�(`6���#��sY����.��vS��[Q��m� �vJ���k�<&�}	�,܋�����<�'n�f��]�g���_>�g���Lߧ��T��R�V��Zt� �I�� AAn�o�ڒq��g����o���0B������aBl�^?��*R#)�U�k_Q��0�}p�^��@V��
Kν( Y�D��hi��J�/�X�n5pg;ǥxR�������MtZ
��ok��&���+~=�����w$VJ����Z�-U�ޖ#UA�^v����B�_F^�a�(��@X;����h�˯ΛT�/rf���-���ќ��~L�k�:�<S���#8/��nî���K����[np�3bh�SC��`��V�t�~j��A�g�%�,�L���k���1T�:7q�ꩤE�W���#���6`�-�X���m!��1{K��B�D�� +�&�M1�9
Ѷ�\C�ٟF�y9���H7�h��I�L���T�ؔC&;�1�]`��J=� *o�b���xL��A'z���hֲ�j�r쵳�.�80a�y�� �������n-]�C�e��K�s��g���X1��3��gz�bn�`���$2�J���.��C�E�}U�pr���!L�G,�� ��b��)W���B0g8�(��i*5�K91��2������Y���u>4�#�&���*;�%h�=M�2��!@ϭ�ү��gD��Bo	�`݆	P��,�a{��&��t���'�/w��l�(-g#7�x+	��������q���V�Q¾{kwG}�^(�ܠT�՝�x�rjg�N�|7;~D]cR����?(�<��Cde��PZ��k�$ �Uz���6h�1���Q`�$��wȷ�(&�ɳȷ�~�U��i��o��$}oC���޹��a�Y�Kyz����>���)�s�&���c]a�^�A*ɲq#�5_j������Os`{�oeӮ5��v<��� �8��/�t�<����{XW9������ �g��S��X��SR�>j����b:���7u8,Q��Vz{_Ģ�0+�cR?[c׼��xw���ЊV��V�K)w|KVJve���G��u��CL*n�6U(���4����,��
�J2�	�"o$&�fdR�Qk#>c:�ހ]��?�F���F8����`�x�yy�0��Z�>fT�e�����:�YN���r�_�ߡS�h��ʒ�dzա���G�ʹJf�c@֌%�>a��8)nł�(v�/�/��ғڏN����N�?J8�Q��Ŀ��ƿ��h/�s-<a���7��p۽-�%���OP�/��5����@-��95�;�r�L��ajӚ�S������N<;�����`�=�43�G�E����!MZ�T8���H��Ԇ۸*��������u ��8�Z2p'I�>J���^��JE΢�d�����	V`��w����C�����(�&�o������Ë;�g&Ë����2�i������~@��i��?��[�T�t(_+z@���کP��ݹ�o����>�M脠���3��v���g�d���(`xA;BP�h�H��j9V�e���v����>c~��*|b���z�%��Խ�fP� ��hb���:����H����w�b�DE���C�sHz�3E\V#k�� NY�UZX�,��>��	�zZM�����2(�;��4M9�?�Ęlk~�Vm^$A������?�8�q2�����T�\��4R�4v"��Sb~d�,a)i�}�	�ʵ�߲ަ?�Os�+]�!�[:��G���Y�R��m��At���j-�7���~�X��}'��)t�Hν���skodE���HP�T�
���d�y{���d�P[:R��+�9�J���&L&�|{��e <�	��޻�@,ÅU���
A79g4���㏽j�c���()�q����S�c�{jt*�j�	i*����4͉��f�K�(z1�;)�&������
��
Ap�n	��ٵE�ܳ�jSz+�O�������#��e?���{EE�tܩh�$R�?z�j���S]u��g�l���������Л:P��L̟,�'�� cY6��?��q�@N���~o`��|�L`�b�)&�X�J���@;�.���Ҕ/����m1��̩賁��:�2���Q@����w�:�@�	j��de�$��H���Z��\l�e)�߅��P��!�>���U:&�d���9 Y
s�����zd?�*�S)��)���A���Y��,�g +�|Q�=�-�[>��AF�鏴�dl���xJ%�9��&����[�]�/5tt�[^���#e�*q��'�FMn��ĭ���"
'G���8�7 L�2]tp�-��EӰJ�ܯ:u+J�Z\m�k'�|@6fq1�e�Ά�Ã�Ra:v��zj��������&G.9\͍����t��y#�:F=�G�U�=߽�IJ�F.�e��9׎m���ṇ���/��Pr����/��r-�DzB{J��s�2��pU[��"afJ������Տ���,�;�_W��Ǒ�,H�3��W8-c��2G�����d �N	�M�0Տ�� �Q��O�����A���^I1��Pf�隬��E=���x�#N�d7?���O��5l�p�ҤQ�,h��=��wo��D��Y�R�4�5���E�3kV�5V��_fە+BH$�.0~�oe����$٭XM������_c��������Cϵ��������az`_��)��~N�I���z��}���+y�.���o�)+!V���l�K�bi&�w�f劙�tO$A��Ps{�t7��F(7��D�c.�i^��\��*�d^�A�'_z�R�]8t���mG�h�)p�&V�Z��4Ȉ���Sc��y�:�g��*N���{u`*������]W�Í��B��oȢ� ּ�6�c)�1�/��ez>�y���N�%6H�+�Ƿ6�����_8{P�h�J0��[����kU�j�b��K��l ��4��˂������rD��Rq}���O�򕹇�.�ؐ�RB�r���
߳�@���Y�L��V�c�$�N`Vqy1Y�O��q�]U�u{��E1���w���s ��S����C��淲���Q6�<�_�8�Zp�=����ǡe�O}���`X���h���>�+Fq�V�6e�ŉ"�K��ד>V�9j:�O�8�.���r�M�ݥ�PI��d;����6w��͂[�##o�}+�2�~O�jT�h�%'S�����V?�b�B���Ғ�������Pͻ���{z�2�t��B����	�B2��p��аsAz�y�B�7�;GN���m�3b,�������p�]�����U��m����#���ȭ�;�<����l�o��P W�L��e�D�b���`}n�2M%~BUnڬ�� ��kjP\{\�8,���V��+/�{��ghCzO��g�6�u&<t�v�}�x�[*'��9�>��� ��$�y��T=�h[�,��[�^O	�~��^cN��\bF
7^�Q �5Vz��Ƙ�paRZ��7i5��(8� ���[,طr��jM���Y\�4�i 8%g�[�1Qa�[��Nr]]¤h�d+���y���.׬���#��6��[�W�2<p�r��Y�ӸpM���F�E���OA|�� j$�]Ü9���J����G��k3y���V���em��`;��}��~ x�
�w�DOY`�3�W5b�B�ѸI���"�8��M�q�`�:+.P�����~������ݘ��R"��84	-z	�~l���>�4����#*s�����Vp1���EY��IX�A �1XW�|�W�Lu�׾�Lk�;?��\S�Hˤb�,��Zl5OԍbK�"��zym�84e��"%��}E�ބ�+��nx̍�^�J}92;5��ԅ߅5�x��o����T�A��^�/��$_��䘲���{=�%8�Q|�7�����`9A5��y+��9�yA�R�@��\㲮�v	�r�lOj�-趷r��d�\v6��T/�Pe�����^o�K��z�#��2���Zo�r?\/���T�ߛ�gP���>i��'HG�m���R2�e%�t�(�O�kp�o`5$|�ఽ��ű��wQ���\���>A�/o�kjq��K��vҨIDc�iM�H�㵡�3
|ER�Э�տ��1/�/���0��3}��b�H]�K� ��/�-:%�\H�cA��_������$�|�4������/K���x���OW��H^mv'3�'LI_E�Ü=C�W�5#���s�4ϴ���b�h��G��J�-���槍rY+�QO�`�O�o��%��\)�v>Nx��7/�$&J���z���o�L��)oW\�]h��̒�a���)��sF탪 z��rFT��FP���n��DDbzi�w�&���߲�¬7��JҸ0��� e66��J�)o�S?�޹���-QI�	�|$/�,e�:7`
v����RQax��AL<�i`D�>�,�=��;��rx�Ç���D������,��ܘ�f:
���<��5/,L��kw ��d��+X�`��蠂�L'��\��2��U���?�Ry^!�#���~���ms������WjIv
�C����4N��& �>��I<6�H��:����~92L�;l�a|��	*ě�N��{�w��<��苡�JӠ��m1y׻��O�+���lu$7nc-uG�8by�
fNW��'1�"���A��]� �p=�Qo	����?r��H�%#w��� �Ǭ���+ϲ.����-�7\b�ؗ��J"[2�!T�%���h�t�N�[�)o�ŀ��К?s���,S�<b��+����@�ݖ3��`��N�2JOzO.�WoJ��e�d�*�v	�h��ßxD�p^�ǫ�cY��������N�?���J}�hOj���,?�W@���mr	#��N�Z�U��=և9%��,v�զ��d����y��Mr���p���U�W��3 6�m�x˙�F�ӐtD��l��E2\A6&:��l���Au��{<�a��LbHCldĐ�'��Q �V�lCs�'.T/�4VpH2�|��h��Sy�"�P[����ߟ�����Ͱ��[r������n�����r|����"��,�$�%�5��K��s9�Ģ �{��������I�BC�o4$oW�{���y�3���-9�,jo&��Ae�+�I#؞�R�m%�ry�>��l�������l��HV�y4\v����}�ݠg\jA��1M$s�s��@�t�?e�fwA�C��,�{�a���I����<��1�7�������YV���`^�|_/��Q{�G�݁���|��	����|��&��ӧ�FAm��Y�>Ke�cM�ţ�������]�����vNw�0(0?Jü�*�Kz!��O&�+�G�����8��w�"<'E�:'�M�W:]`���� �D_�ܒ1
���e׀�i�r�'6�,ta$���������B��W֑�@��j{+�A����@�vJ�P��j��|��AlVH�{���!N[��"F�_�D�V��n�3RG &j��_<��d6+kʻ���e���f]$pX_5[��+U�Ѓ��X��v����K���x��W���t�n�����f܉��M1>��銳o�̀~��g"�9��ʆ��	v�,v@t`��,;\��Mx����)�'	 �I��4�06��G���Y� ����r��;�UP��[�sݸ:s�1. 4>������n��N3
w.n����F>��*fY� E?A��<�P���ɾ&3ߛ�Q���y��%�Ka�l�ҴL$Z�O(#u2]�<�֣���"⅛������Ff��"w��D��k�k��~&���r��N���������2���.0��"��Y�&�ٮb�(m�{L�%�M0R���>ʑ���oS8���h�7&�+���HK ����N!g��q8��^�v�D�;8�I�Dd�4�0�l�KhR�6�v�3� gd>p�&^fژ��gm��g��v�Ռ���sJ��iO��6�(���3�
]p�tO�R�z���ɼ�5�W�8N�zr��7ź�?੺��5�o�>���$�.��������Ep賙����#�F��/���,A� s�%g[���2Nc�e��_u#�)�F����x�P	1	�u�Ɣ;�g���0���6ܥ#3DZ��D!�t��Zr`O���Y#
P�`1�	��V�,���{E��Q���1\/2mz,�[WrlE���+ I4$�w5,��¸��4 Q��GɎ���gj��ֻ�Lh c˽e"�O��:b�[��"�Q�Z�<��3j�KXl�S�t�h��K�BR����t���V��,ҥH�%�?�t�u��:���Jp��1�V���=� �bu���.|�j��x��2 ~�L?x��m!0��ؼ���&	U�_�৽�z�h�� ���;3����Ua��㝦���jJ8��C*pȟ��ݚ������W5Kr�3�E�=��3���b�3���3N���csl��>c�R�G�ֹ#��=H��;T������)i"�+�U��d�1��=�<�c�Y�1��2w�����u*�������՗���W��Q��u�0���beI�t��@59��,��bbIԾ��H z)f(�-�����z��6�T���s��?������ 1�I��~jF��	o��j��8N�M��I��c����~�ng�T	�*{rPצ\p�&B���������⠒:��'Ӽt�X��#�z�l�ˈ�i"Ol��"���=F05Z5?�σ'�R�}��NZ�Kr�E����ø[},NOt:��/4��h�3EѺ��U~��c���q:��\�XZ�(���S��D��j�`��:""�DjpR�bX�l\U�z0o|ɜ�@�+�d���	��M���Pw~���+�5us�E�P�[�����S�e�]�8����g�XP��s�*U�v*���,�6��a�	ɽ��H�sdY*UR�䂨_;�g4�q��D�c9N'K����H>�#��'�	�^��i���Q��ש�#c�)�u��6q)?:�:2z{��&��#~!�6�� ˨D aA;�ds&���;Z����8��X�F���|o|���g�j�R����`V�#��I~`����W�s��'x�sɥ��^{�*��V��r��P�A�$�p��Z��{���t��3ؖDI՜��!C6>IE�i��J�o6� �X��V���F!������g/���z(]&b2m�FA0Խ%�6O����i�w�}8Ň��;��]���kl�is�N;~cL�R��ϔx5C=�l�:�<�"���W a@j��ӗ��e���t*�F�V�&�8�ٝa��Q
О���,�}�K���m�n��|�UD�֊x�с��(���T���5\�pZ&��.+y�rW���Pp>-.C�>�Æ�5��Bǩ�ܒI�I�w0�h���0�c,���ʊ_	ˢ�Kv�J=�-w�Ez`H�I��;q�|�J�!�g��C���|�T�5���"�ʣr���
��wkmaX�����悔&���b/ }9ֻ��$�_R�vЊ���Ō��~��'��	oɫ��9�ќ�37�37��u�c��O����ǌ���geKNw�kH�E4Kiz/�:�^q����5N�ڛHF c�����1v��jt�AA����⼎�Z7��"j��KƤ��͌Q��P⩰��)����W�~Z�@W+=��H-(w!9r����V�-ʼ���p���y���Ʌ(�ݾ��g�2���0�a �F5v
�O1/�O����0�"�:�8�3�$q-ߛhA���m�
i�0%]�F.��oC�n����
��z�G9��h a�Z�L��/���]b�>^��w)��3���4�}���#��/� R0�X��T�/$��z��9y����,�G~�9�(<�3�{+��/-���|c�r �a'L�>�M~�;�y8���7��
�>?�G�V���Iu ��Y>�Ɨ���J&�U��,��>��������T�b�݇BH��>qw@uI��ߴ{�D��BQJՋܟv@�����}g��1C��n��2�-pMJўhI%?m��'���D`�~L��mz��D�f�.D �j��Y$�'�T4J���}+�iM�����H���i�i�����-�u���RuVqB��/��h��=^�x�E��(d�lcc��]�Ϯ&9� �[�a�
eCb�}��0v�ѻ]���!��snM>#B�(�1�/����ҋ�&-�є�A6f�F��i^��c9���+�L��O�LLk�JM�o��#��EZw�6��W!��Xy�$}]�
�1����"����-�,=D���d^B=�c
ŵ0.��,ܸ�8k�0���s�D]?�_J:���lBc�6��d]ED����v�!�����Y�^{��c��LA��D�E�|�ny�� ���m�`��A<�����R�H�[[�9�������;��'yo�7=�<>B�2�n��O���ڐ��9L��w�o��t`���[���@��o���k���`WȘ�Zx&O�b2�j�٨�1m�\4q�
f�0rdz�D��3xaY�Ο�)u��m㗧���I�}��d�F�8$d��ۈ�n�_hm�(�p�c#�9y����LN��r������X']���V�����XtM�1�M�m�i����P)�{�@�3��:0�h��2��)��I�����@J<�!���p���^~m�S/�V��z\�)���j�Q�r�J�2W��*�3�ZC�06��X�lO�1�yg�X�m
O5My8n7~Z��Q&IY�����qk��٫
弤娡�����~�L�⻹�Y^���ࣻH�w欍���2���@��>�g��I���I�{���0:�Y���܀З)$p� �І薏�q��R*�L�������&�R#��4�UXNR�j��h7����p��/�#�u�AߍC*y4�G'����Ak%�T���$f0�R�N^N.�b�(g������jd�,3��A�-�rү&,$b�0`�(�����9�1��\��Y$��]�fz/�@�hdV&8t�J@��`�z�#s�-��M���3?w#PôDp"{WV�y��6��`��.D�o��`D�~��N豏3�w�r��I4��f\W1�n��o��vP$�Z�<�@�u��Ng5����p�刾�s}|
�NHI��k�z��ޭ�ֶ�c�K}��6X��laR&[$mj�5��D+k��

�ί���ݺX	�������>��\���r�'AV�����j�
���u�odG�Fb{ua�YlhC�����U�F�f��ٻ��E��M��������P��3��������\WslG8!l6��Goc�ko��S��s�
GV���w��/ThP٣]EA�r'��9�W��eYl8$8��h>�A(@i8ڿ�zL{�.��p�����Sx�y�d���i�Z��(�6*��D2=��HQ��L��i��;�f���z��CIP-%@'Q���b(�a��E��]�٥=�$��X0S�IȬ������a��Ӳqp7��'٧&���B}�z���n*��q��/��F�=2p�(Щ4�,������S$�}�!��S<.�{w��Mo��ST.�a���He�Cm�?A��2r��v��+��k���|9��6덟��9���V�8Η"%�్{A�j��]�{W��y ���S������ht@��X�����G^^Mn���	2�_�`�t�	�d�}u�Z9�?�g5w���Cw<����Yn��悡����O	;�!��Ɂç!��xگ��d��Z�,g�A�N*jo��0|2=�J�"�S�2�&�37�$`'�h�6q�+ٷo���|����_��dr,��l��	]�_�lԌ]I�ݡ�Y�*JR2�x �0�k��~N��<�+	v����J�&�Zvk��7rV�f��| �'���F"�Sk���CS(���ҏ����-�Ε,2]Mb��2�w�9[�H*-�Tq#ιИ6s���ɟcz�v���E���[��cZ�(T�n�1G�b�D��(���@�b�uy����+e.J+Z���:���h�e�������Zى��wS�t������EZ�0!�245RRf�5kr��Wm$Ȕ`X�_΁Zsa��Rݣ�ڕ�>m�ef��V=:�{=��tar��Kw+%GŜ��%o[�F��U��H %� 
�XM�l�Y̕�y�KIß ��5W�������0�s��W�^E��*\��nD)!����rF�=CX���l eז.���ۺ١�O�y�f�cGYG(� #1��?�I�-�Q'��i�2�0x�։���O`�Ɵ�[>�[^Aڹ�.�ף���ӂ�J3��c=Z�l(�ϱ6�h"����F�ܫn�9n����_om��>�#������c7�b+F�82�=h9��?-w�;�D��J�#�{�4ǻy#a`,%�� �Ξ�!�f
<tQ�N@���ȫDƧ���洕��ʔ��-�|�x�2��-�˨̝b5h��xu2�8�j�V�D�[�&�}�,��Q�(Y(�쌓7h���@���f&M�`ZYC��6%���W17}p��3���!.�ӣu+��q1�T�b;ŧa��\ W�������A�rO66��00Y��g�5�V*����R���h.Yu�so�1',����1�4��%#p�2� ��B��?qX����'hU�>�FD��%1�x����-��7����,��~��E���򝪖o=6��q�^�	FΜ8J�G�����;"Uo\�u6 z�rs�$�b8m����]�b+��rr�i&����|ژ��F��0�Q$o�'t�38pi��a.�~���x� ��Hz���,m��Ea2��}��i��{u7jL[���V̸w_�t�0 ϳ�(��Jo�i��sC�aV6]�_~p�g�g�Zp����嚖�,m��ya�X=(�?WN(\�;�3FH@��@ty]�) �MP����Σ�qu.�/�O�X�QJ2�*�[�qRM����b���ߒM����v��� [�r�O��Op���{FW����D'|r��'�rŽ�����+}o��w,�*�Έ{U�=8��+���}n����\��'��*��
�Tx����C+M�P��@>�^����ە7o�u�z4�Ѻ�7��b�4c:+Z�O����&4�J�#���5P�]4��(��ܛ�K���b��=���tS����T��w�e�,�>��<����j<��N�H�+��	.�!/�;`�z+41SrQl0
�N� ��B-���3�~�P�C���	���A�V*�9�d&�yC�^T��l�!�B����O����4�Aa�(r>13�RKh���Q`��oT
��]���f��Їf�d��*��k<>��-��Ng����Y����0�U�uY3ŵ���X���ec�2}Ю����SWA|�t<�|�����\� � �~U�a㪚�S�ъ>�U[��V�����f޻4'n�e)xM���qg��E�{z�b�u�X�X��B����H0<�2�V���#0�r�a�3t��s�^n� }7i�`I��n�1H���ƹ���'p�&U�v��l�w���p|�JS��^Wjz 
kp����J��_����~�'(r25���WT�/�������pr����-%�p���x�a� z�햭������ Ē$�Eo5�Ft��x��(��GJ��9�͑OZ�Z� .a�-P���]�� il�G֊��|~�w�B(��+� }m������J��xQ\W�q9|[���"�"<�b.�  !�&׃�n�C�i*��;j�ʌ�RYYeVv����3m��X�	(��������g��qv��,Oj� �#P��i�P�p���"�(���)^�Gh�B6�5�v޴ao}:��'���峒V[�oω�cs�=k�.k&��n� +��7W��r
��,�m�eD��XXcI�i����nE�����o���@�*vY��/C5�n'M�%�Ǔ�I�M(��Ƣ Pb7 ^��$���np%m?� ���↠U*IG��t @n��^���&{�ư2| ��WM�����D+~�ޙd!��5���[4��܍0�oֿ���%�����\���)�"� )�{xp�ңKqs��{{(�Ҥ���d�����)��A=��;~���(��B�&�b��[����<.��VY����8S�K6j�����>�PE��O�%�B�.^�K�YĚ\��l�N��nO]^vL_�%$>�ʩ�u5�cP0����j]����e@a�Pz[8P�aS�M�J#ȜA�y-�y�YꥰBDmRz��]C��ɉQ��ڪN?C1����W���	���I L�`<�y���h��,:r~۽�����J|ݐ��P�=��g��$Ⱥ���JIS��)�"���%ƴ�][	�P����e��dd#���p��G:?���P�]4�n��ᗃ���|�RI�>+��Pi�BHk���elUU��5?4V��-��vX8��A&�,����Ը��h�Y:p��\W�.)*L5ɉ��
F��NAc��ge0u|���wd�RN��S鉵�մ*,���e�4���ڵ��roo�4�5ַT���iW��ե��e�t�ƹr���"���@#�ͥ�|��.4 ��%�E�Fz�>�fNĊ	���w�	�T�k������2-J��(�A�4H@'��H�vk��]E�M�Ψ�Or?7u#�� ����r�u�:֟�߈���N�5���Og�ч4VXb[�U��u�_�fpuZ�Ps�M�d��o�-}N�@&�3{���+@[�=E��4��3-���x[�������Y~w���r����$�bįj�4x��K.f�t9_�Jt�i|��輥��?-�bΫҭX� V�1إ�|Q�ܷPʖu�$��o�B�
�H�x{�g��i]�h�ì̐~X�J�^�^ 4���/����fl_�%6
�`d;�J6^��qF�B~����� ��<[� w���+b���S���Է-@�@(�W�bŷER���ڃW�W
O�� �����X�m�7�Pd�Ͻ���~�{���7��&�����_����ݖ=i�-��q:�&�8~H���b��1�c�IO�)<]!�Au�W�-,��W-���hW��";u�:z�C !�c�T�$���d�O�s��{�)��O����P&_��� ؂ܒ<b��Z.��б�ίg���E�_����L�������g}�I�BҘ��=�$vg<h��%T ˰��d[@��/{"mJԮ�-���=H�%�- BM��;�:XNI�74�le0kN�tIt��g��Xr?�pb�dL}d׬��xhWn�;H0��wh"�>a�j��7_M?�29Ӷ���a��l��|C�g���z枹Z��&)�����{D��)ԺvS���̘���2f1�4F~�?���P�Y3TB��QȂ�ګ)t.B�Թ�J�R#-ld���H����h������wF� �?��j����S�i���0(ldnV�ϭ�*�0��;}�MU*,���f���*�>Ăt��X�F�~�NU�j�N^)� e����Wpi��9<Wl�u��N�0F����P�c�c�&�J��=R�ꅳ5�1|9���$�q8�����)M8"o�~`0h�MW�.�x�,��H��n��+W6�
�L���a��up{��`[�T���T�W��
�V=��]6��(5Ny����z_:T�oYr�����/�.�
O(����<��k�{/ !�C9Kw����L�
%/�L:�Cf��'�c��^5��.1,���Z��#?��`��zέ��}D���nL.ș�5�v��(�����4E8�3;��CJ�#�[!
!$���m]��w��}0�����&�Y�3�m;�pෳo�j��3�_
ԓ�7~[�O��"��Es��/���P�%���x45j����v�T[^��$���E�,B
0b�@!Vf�uUw�V}2P�뒱�8��*� G��[w.̞� 7�8_��ۣ:XWVAX����mȁ�Ӏ���KT���3\�q�ߣ<�bnln�������`��l��k\z5>�u"������͔�󲅼x�u��u	����S1y{`*��-4U�sB2"�0l#��ICwֻ.���	?���ɱ�̈?�Yy'}{;��J��86eܴ\D��VM%ˁ饯�� �B�7u/4
/fc6���2!�P���;��)z����&ȇh�t@����V��]pv�7��:ah�_\�D��Tb
{
���61��Tz�4 u�:җ}8?��X|�����1T�LD]M�r��	������	�����o�������5�~�J$�v-F�bgM�^M�e�+ύ��N��o�;ů���կ�l�I&��Mt���H�z���J��_�̞ i�\��]b�;C��NNi���y�Y�����r�"��#_��!���::Iͭ9�N{K0d�>8{�pJ��",�mŕ����G`�Q��\#t�����#rc��Q�Ȳu���`R��9	��.*��H�ZM{��4|�ƅ���ȕf�����S�-Ozp�GO�"c����,��ÔH.��)Ć�_3<'��w�p�`�:b�</�uS>J�&g���8g}�?�*J[q灈��0�Q�H�6�"�~�
;T�l8+}K�Ж�je���c�p�A: �sY�<~�����z�j$v��~�N&8�:�7r���m�M}/|��]�SsC��=�L"�����	$>,�Çe��h���St�Ȕl��4�%��XK@yw�'9�$E��V�bѤ��M��O}��7�X3�*�h�A;C���0��XC����-h,�v.��ؔU7rה1�H�7�M.��%78qp2��Q�"~SuЬ-����l���C��3�Li�3�_2U��>	��r��0.�6'h���AqhlBn������h��T�˖\)gq��z��<�X{�V��ʊl��@`Ԧ!/�6��l�?���4E����绍{QofR6���қu��Y�T�pa���@y)��]Z�1���㘿QKf�?�r�J`�"C'�OS�U�����3m�c�s�H�M��_�dG�b�b�83Y%�=lf�񝢩�GJM�VNE��zj���Z��q�UK��˭�wy��9^X0�4Ģ=v�g���u�GL�&p�;a���[J*/��*o��Ϣ�a���sQt���l���7(e����ܠ�S�^���Pu��&�yX���M�/���̽�I�oX��X��!��r�*�"F�m�Na�Ƌ�}��R��r�ܹ`2��+�V)^oLꋾ�7�h�c�l�Gz�6�1h&BJJMi6@����˻9��7��o�P���3J;b�U+2kk-}G��RFT���l(!�:䘝E�6�͗QbWB�&�FwaKJ��~�"�5#<�+×B�$�z-�-#�#�N��0�Bi��}�G&>�8�O�)?87̗G��֭/�!5�I-�'�pto�ǬbN�K[�\����~l��d�C��������oJv9�I4��TyV���9q��?��\쎧�TC�p�ɍ�&��D�T	t;�G�+H����6�F�f�X���2��������C{��@Qi�2t��Ք�~D�Sa���+C�!��� �F� g~���A�hڕ���|�U�#= @ ��]�$5I�i���ߺjE�;�/@�r���v�`w]��_������r$�4�f{�Z�;��P��\��B���
N�^Lװ�;p��8/U�����=�^Ђ����,�nв���\�l���(���UY2���@�pZ�c�<�܋�{E�G�قek�Đ���[#� ��	��� M���R�Z�9�&�����Ԣ�n�x�@h-}���Bj&��T���E�ƍ�u��.l�Bс��{:�nUz��|��+Pw���e�A{�.��+s��%N4�Τ��w\/QT��zR�xg~fI!ٓC�9��_h��[7��Z������E�׽��Q��6KV�1F+� �0�o�Gs�l	�9&�	�'[{Z׸��I�,H��Y`n����"}z�3VΉ.> ®�B4�w�P�4Y���]�֏�����v�^�3����*q�����0���$����z���Qb�E�b�d���vB�~I�֍<C��e���
�C�Y>��'�LM�� �_����d*!�.�g�&�3��p�Y]�φ.W���_�˨ѳN`J�bq3
C������+K.�6������]j���B2�
|�����[3��/;=Y��V���&V��t�,  J1�5�� +�91�G���/<�I'��Id��~��?���xD����T�Wz!y��U�(K��+[R�S�����Tgz14���BK"�|�"28���>�i�6��#MK��.A7`]ٶ}\�aS1+
2�a�b7-�5���m|�P@~�N�U��;Ľu\���{�j�)<����k�a��PA �ǔ����ʈ(Xh�3q�w�cG��-:v��`hv~#~�j�!K������n����1}��*pyH&2FM^O���s��I̫B~�͕�7��ӵR}#<�3]��7m�����7w�Ps�|���ӥ Eh�S|Gj�n� �?MU��7���Ƥ���9���m�LD_�	�{�	f@�}����aE^���9�^*��5��n1�BPO�ެ���Y���y���K?S1H��Hr�j\z�d�rw��ڒ�20�r��P.GN�j3��eM5��B7c���r���Y�wO}�r��P�&?�џR)����1[&Ki��d�1����� �i
�����W����r�d7T�������x�odH*q
즫�,{��E�(��� �+��~����?�>��ŬAۖ�h��M÷�ݍ����'��S<f$��;��
���?%j���-�k��&�#ȧ�8�f�f��� �b�!�+���^�Q��b�c�,�I�w��vg��9��v���6�UR:�:ү��݊�����t,��~�.
o�j���M�o�"�:�Ь��@�q�	YR:�Q��Q5]����I��K%�6D�S��,���v�H0EAj�?Do8BguN8� ��͟UI)@���G&�"9�>��?�b�X�)p��nX���J����}5(AnE]pg��)�Z����ә~ҝ �ŹΣϷL�8�	PWg��� �{a��'?������|�
ך.g���CfG`�bs"���9�'��f��;�􍞛�:���4��ׅ�T�yЂ�b�#gE3�[F`�XM�?����
�7���"�:��;D�
�N�� ��3Y�#A	Y=|�!����Q[P�L�c�VTA#m`D���,�<n������H+��N�����\�_���u<~ϓJ dP첬+6#����	]�L4L�����m�����vU�u��ZqZ���Wi�}:��k~�]�h�)k��!"^��Ze�Al��q��2�NG�qp�{�7�)���&l�Q2��;�����
8�ꖒW���u<d�R-E��X�����"�6-1~��O:���ѩ�e�\�<E�?x=�{��<�XÅ�3���jeQ}����HCŕ;X����k����uӁ,ώ=����k�]/�;K��<�H��D��d=�8]:��2VY���[˲��<�6��Ro1�������f��������J�1���:����o1�7���Ov?�䋿���*ǎ�yQ�TC0N�٣��'���2��n`eU��4�[f�q��G�g��#���J �WW��G�Xd݇���
����Q�
�S�%����J��I��	�I=�֏��SG�h����H���<?�^������O�����I?�8�&:�Ӂ�,ú>�u�Z�/�	�9N�a�\LL	�}-�S�nղo��&'���^�M�0�%l�I��d��1ޝ�H~._o�m�kUb��FƢ��A���Rӷ�,��� ��@��P�<r2��4��f�QF ËO���������/�yT���<H �c�o�/[`a�}Dz��{����������V~j\�ru��"���QT���&`6��&1���l�;Y�br
�{R�Q�k�Ę����=�+��A;�o���
JQ����u9����v��O�B��Y���B���e�q���q��p����I��	/#u�}�����P��{���e~��\ [�Bհ��\C��O㰸�K�ϝBk*��Nr��>�mHq%Ϊ�ɬ��N�~V����0m���ʙTEe��i�&��5�[��g#�aB@V5*aL3L�Y>;��G���B5�mC~Z~up�\+��W8s0���B�����N�aN��"�˻b�s"V�b\鍤�������M��V������������F�a��,G�3� ��	�jK�{ CR�UeZ�?;�֓r�l�Մ}�?7Ɨ=jFF(����:�Δ���0#���q�����"�x-���L��(�c�58�R4M[טh�:Ķ����G�����i��̈�/U�>j�CVg�����6��׏�:�"k�g��䐬BQ)����A��((�gHK����G2� �o���o~���T΢�-�������׃��S���@�8$"`,�H<z����n�S�����}"z�>�Q1�ȲW��I�pE�m��yD��9��P%����lpJ��d��&
7��֫ʻ��x�~����W8�{S��.jT�
x�p�ьi��MF��$I0_�0=�E�����/&t�{��8���{�e%i�*?�,����:/�����?�ҡ吿��O�&&������s�׳ʀ�v2"t/��+.����k9�����|˘����sLH+l�Q�����8Ǧy�u���-�Ky�,�q�+CV��Ej�/����p>��b_��M��tK�ho�Ɓ[w�<�k*�P��)�7Sv��YF>��Cp��"h,�}��Oe�)a�dr�&��"ݶ$�Q�+\���(5��GY�yz�R������%z�����ǀf���ƚ$��������#��jm��3���#"J��L�Ϩ;�v+�"�ag�{W͕
�ޖ'�mn�׾�������D�#x�ځ����b����BU���z���Z �o��˱�ڈn�>0�_/��rՄ�Z�&0k�pF�Lޢ�Ft�1]�{�SHe	���u?���2>���ET��e?:��n�����.�@:)�t*^& J��;ru(���R%$#m�^��`mP�k�F�vv0y�ܐ��=�y6h�w�$�����Rՙ#<�U�BƑ�e^;�g�� ��\��HTq۩�d���{R�S#z���vP=��$��]��=�������M�6�aB~zs���lD>�1K"�z���� �b�6�P��,c�1���#}�M3b���7l�
���D"�
�Q�AO�;��̓@�xQ��Li���C�D�L���%볈���tԊ�"��ئ�c���P^`52�E� �@[��\v�[f"̟���<1���VP��e 3~�8�_�qн��PPeC����C%¦B�vQ���)�la��y�a����5�}#EZEEN�%��W���F�ޥ�nO`H�.�W��p���jNpC�bhU�*�{��1���:Ha'/����1��e=j=Z	N����}���Hn��h'W�ӏ�ZǑƖ�X�E�wki�?�k�0�Z��.�������, �n[x������I�_c�o�v�f{ϯ���H�K��>��i�z�LmF���B���I�Lo�G�1��G�#�q�	Ҳ�a��P�7�<�o$[��f�Y�����xi\8C{=�M���t~Te��di-g��b��[��/�P!��b�k=T4��:�}y��!эW:�wo��C�:3�8߫��<`��͓ /<\�)��a���O���	�$b�gP?�-�1Ll��b�l�t��_�g'�9�Q48o���gD���)n��s��N$��
�h�٤7����x2�椅�B�,�������Ka��2Ɣk�{4,�%��`�C���/Г!O��k<��48��.wX�{�/�*�����4 g��;l񜼚R(>Z̓z����걼�X7�R�"e�2���Wffs���ñ�CbV����;36�M���/�h�n������a�mhm t��Fd1k&yF��P� �=�t�#�";u����㱒�ƀ����)Ak0m@�B��	��!��̇�/ K�N�+Į~`��Q��u��D�{|��^���Ɠ:�&yq�oZ�w��Y�2E��%���U^�ؙ�v<}2�u��m��w�č������/硬�ئ�I��˨(�[e�����M+�\��L�͗��e��Q8�����u�������i���Pd o��3���.MoU=ԟ����Ή�:���ѝ�Thc�&���0�,
C��)VK+ײn�0��;G� �UnH=����TF��r@KG�K�DO�E�����;M 
�~A'��
+c_�f!T|oc��o:I2>��X��gC�;���$	-z_�@	C��(4qŘO�'�����k�d���zo~����5�"xT��1�5.�#��=��j~BEk��t��١�
2�>=�Z3e����"�S�DRzV���\�6.QWy�`�'G\*�د�kQf��BQ��2�B(ϓ�V�$Gַ�ȖM�s,F�)޸�K+�i�ϛ�Ȝ����2�1ׯ���Au-d��5�0��MX^��! �׿lb��<P�_�?�R�ɜu�PY��&���~� �qQ�s:h�V~����tI��SL+�yD�5�7�Я����a�4�brFli�U�9*�w�W;'?~/f%m��=%��p�S���n���k��V�̕�#ҤLh����^�QL������L�������A�ͧ� �29�Q�`цh���$8(GuN����X��[��u.�8-=e�W�r[�A�}Y:<n7Xm=�1�*��|;P�B��K�c���!��lY5�M��j^��� ��+Y�t2���>�Xļ�������(�(q�s���؅�ܙ��<��O|Qv�Q��_9	/N��9D$���b����a�|�\'6���5�ϛ�Yj���E�.ʖ�\y�̃:����e�q�A옝01��ث�3đe�[<�-]\��f!Ǩ�vR�E�gh��.#�xY$,*�Jj�c�CS�s�@A�!L�̞�?ݖb���a�V?��!ԝ{v��qu����5"ݭ��f*�Au�����;��8]��}� �Q�a��"!�-��ؒ���3��+���`��O��*��1�1h:�>Yk�Y���\�r'6��> f(�>�F��:��RX)��#'_��0&��gUG�*�!�呒���ԑA�vS:5����w�*x�s�\���<��6�ff���ƖZ�L��c9
i\�7)��}�ya�u8Ӏ�_y ȍ�^�����'`��z�eӕ��"��l��i��-���o#�>WKg����Ԁ��,�>��g�'ɫ2�u^�ڒp*�`� 鉚��_������
���T��^�~(uEo�&Oz�շ��1��d|͗~��7`F^�/�x��2:�h�5<j K|f��h�U����*�& ���R�| �C!��Ev�ןo	�|�,��nt�՗i}�LY�<��@��	���"=� Ag��cW0H�x�zA���3��a��MʡD��]4Z�d��<ڠ��y���{ӓ<�� 	��2�O��FA�Ԯ���7���Q	�6�v�p+�tNO|����Ѵ�䚽�Ah�1, �)f1#��F�jUv��u����"� �)&�%%X������WYR�C��ssw���"^�ϸ�v�� ��x%K���P`�}.qAW�'ᝍ���`Á� ߰i�S'��VJs0Tj*�)�����|�d�����J hNc���v~�h(��a�4!�r֑ͩ[I�U��8�e�y����x�UM�)�t��6�;s����?��tF������S|4�ɱ���a���