��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\�J�"�r!�_	�Z��Ѵ��n���e�"���?k����ƽ���Mb���J���$��-X@ʫm�b����^��������m$e~�� ���a��j�h/� �������R9V>D�0��s5Њ�����Bko��6v4��s�q��p��U�|��^�ӏ��!Q�`�v�id5N���L��Q�q�B��OkNjtf0}�"�h/+�&�1ko���B���bB�G��z�^�>�O�;L`� 5�U��#����O��i�[���.M�s(�x-7.8w�[�K�z����m��~&A̹�
�
X���nȻ����~�	"O>+�|p���zG�`$fי+�\,�uK������M��d�d�m���s�"<�-�RW\������0�c���Y���sڽ|�ޒ��q�>�~��ws��6SH�����|��8���e�ӵ\�^w��w�m7֗їr(�#��h�%D�K��)}�x�7r���/�0�y$��U��O��Xe��Rz����_\�M�<Wy�r_�k_Fpn� J���'�R��u�E��t<��ip����zKQ����)��a����7�Q��}*�;U�_��3�xO�8V��	�%�v�����|��v�e?'��Q�����*M���U�Ԃ"~����Zi]��մ� 2�f�Ys�*^>�>s�9�8��	������O͕���O�4��ނ�^�Bb���#�!9�H(�Y}��^���)���K���\w��2����/We�/��-���	�E�^o���O�ӡ���:�}Uz�~����c�3�R�u���L�kJ�����|Dk�R-\ˮ��#(�*6���$5�z�a���/�GiaS�Ļ�F%m�'e3�����VA���|�D�\r�bLa���z�c�T���Q"�����Z����=k��5�&'�VG����(�zso�v�A�����L-�i��+( ��+>����5H�j;�AĲ6��Ř��[Z���!�(ݔ�'),0�(n �^�L	� \�����E�?�aJ�6ѭ+G��G��Lj��[�m�u��5��Vz��(��[4a�3Ԃd��<�ꎤj{�kV�����vmD�ME�>5��t�`7�4��v�kzB�}l��7BYI}��"c�^��+52�?{�� �
J�����͘�����7�� �o�X<�A���d���<��8d��_���T)[}u�,@0���+y��Q���X&|d>*ӹ��nV�$��,+�
VnEg���`����ZUB��T��ɒփmE�y�3� �Y��� S��r�1�M��7�3�B(�:��"R���ȉq_��>xm����N�n>?�>w>��EF1���/��\d��C��O~tí�]�/��E
��[�Ty@�8.�����{��k!��:��nk��7\��y���5 i_v�R$���
��w��=(׏����eR�3,E9��L�A�G_Pia��z<��.@\��\�'�-s�X\$W*�;SK�����^<�0��-�ʰ��KI�&�Y8���Ł-�wvtԻ��LM���'�:�U0�� ���
�S�	:�ܯ
�1 ˅jY����F�U�aK�����7���~��{��o���0��^S��,S���5���}�W�XT	�°����m8�l�
���j����:Z5�8�o2�����\ם�6��N�g��u�Dg�(/b�2��)iod_�����h�?�΃��ʹ��u7�t*�O�*�Űt������I"k�W՚(�V�Ta���x�.##v�;h,�A�\2�ĳ�/���v���q�����&�4�u���*�D�
��3m��Qy�&J"N�K]߆��e����ı^D2��J��s_� �W����SHG��[��ڊ������\����%�ﻀT��}�cXd��C�gy�(*Y�%�A�v.N;Cf>KY2H��)v�&.�m�&�t�L��Q����������1,j@M/��Q�رhB�=����6�9�`�]�Q��+�r2�
�Ch�yB[)�~���_�P��	�g��=��q��gJ��H}>��),�KJ�WƱ�&������K;�C��� �%��X�����i���7=c�<�^�;�^�+Ȁ��I��,�B�=*{Z�o�JE��=|�F�i1�9JM����#^n��j�[ǋ~t�ca�VE��m�Pd��y�*?���AȖ�--3ihZ�4u���%�[Z���gTK�&�=u�٤� �gZ���vH*1�t#�&'����,�n~w�a��J��y|��k�G+��j�AX�[az�l/Yi�v�`mDN��<�Pg\�b˰�c� 0����4�.�(E�O��9N|悠�z!)�(�a�	z��q#C�k�����Q룷����M9B�!A����y������n2BkؘB�WTW&�Y��-�ӹ&l�<�s�FY��[��jd�������%h�g�I��_�s<E
3���_N��7����#���F1v�P]揎� �ε��wB�e�*�w��_������B����}��8yA�;$4�򠁍�3�����=nR��L�j���[��X�6n|㞀Ԅ�,7�#I/83��k�������S�8CM��L�x�H۞����c��H�FV(�6S#�(�IO#_�$ff\I+$u��d�ok�(�����@��őC�s�LS& ����=�v!�p��/	1مr,���<=X�P��%����~$6�ZK�x�e�X����v�DcI�,����!F�W�� }�e�āe$P	mp��NYIJ����dfj��J~	U\qޡ�+oЫLm(b��>\:_��w�y�:�)��h�����P�(2�uk�'��/�ƞ��_,d���hG#�Z ��8C,�v�ؽoc��4#]KB�v'p^���|I'�y�KX��?h�LL
"�
���ǭ'lT���ZGJ��9�+L����#(E��.J��a焜��uP�D,i�-�~��%�����*�Xt���R��m姻j����JG�,�@~*Х����#	x$��.���d�f
?��%DD����c��$���h�t<�EM� �x,�4�+�3ba}Gʳ��"�k��Awr���j�"�I��Z#�.Y	oO� �e޾��rz�K��J����$j6$.�!�3b\�l���ݤ��}��e.Xݧ��x��S2��Ibh�����h.sg'�!�gC���J)���?)Z8���/ڒ��&z8_�A4���xl��w�+�׈&'�q��Z ����P�f��LPx^��X�$��w��f���Vm�w�N;+�qYvm�;�����az�F��	��)i�d��ށ��holQɸ�T��~��ԯccWA*zRC���/*S1Ϛ�q���"B�$ü0J�-�޾�H�.��2�������������^a��t�߼]=�1������̇���C;r�XL��>��r�S.h uN��M���[(U�5|�K�4�!2��3$X�'D2�����K��Jw�=�����;=����p�C�:������b��H���،�o5*x6�Ya+%!��p�l�LW>`��D���NL��c9�u�|�]�"��uZ�=*{�xT���"�O��%1x3�����9� �ܣ�݈�ɏ(p��O)}�D���A��*S���%
�Fv��	���}���������B^`�W
��E���4��6���75����7�,��L�g
���h/`	�o_�Ӹ�z&��ϩ�WG�k�f`����]�%vQ�}A	ݱ�r�Ǫ� _��+\�W/wz�l�W��\�ُ9��:���������C!��W��z����dGR��P
�@��Q��p�/Q+�Tޘ�n֑)���ea}���j1Fbś+�i�I"ĩ�Q ���*aH#��`I�Y,�L�INh���u���D��*�G����Jzob�4b�_3%�N����#U�Rf���z�����*�QH�c#p:LV�t�R9�J���Z�|�V��@����`/U��f�<!�:���� D�߰~u���s���1�|�Fa���6����r�ʌ���pg#.k��e�R�P��f�HB�/�HMx%�{{�7%9+�hUO_��g��<���UF�K�Ӑ}:���k�a�16�>��N�L��G��H�� M�|p���j�v���P�=c������|���܈�B�e����cVcd�!21�o�y�+�ux����O�vY�������0b:���=?TUEh�p��![
��;`i�����٭��~�P��t�ó@�s�"p-��Y�ʹ��ݼu���vh��|�|+��݀�%Q����V����������G��K4���N���s?��u�X'�����F��r����B�ޕK�y�BHW�Y��3�C$��첂g��V��!�]�^|x^mN��=R8o1�(�
C/��=��g�p]c2{��}jb������0-�eK"�	�潱��[QG0V�G�����m,xƛ�@&�|Ű�m!2��@'?��57� �btT�E���6�	ʪ����+vǨ؟�s�Y�ɩP��1?ܟDPA��T-�@�S�7X�Z(5�BL���s�ޚ6?�W.�-4���S+��C�p�Fڷ9+��
i��Ht���l<�����t�=m�O0���~ Yo1"C��Q�IM���t����pT��Z#���	�g�I�϶Vm������%B|�SEw#�HW�yG�_C`�*�2�E&L�5�^˩�0�(�� P�	of��hqo<�W�5��2Eކo	���k��9.Yk<!��c�:1uճ�;�9�伦���ZgOL�ࠏX�j��VA�b�a�K9y�rRr�"���hD�~�Mݭ��i�Oa� 1%��o�$���<�����Mp�㒈׮ػ�s��J��M�s��!��	K|��<:d���^2� "���T3�ٴOѝ7�*<-���������LP�e���:�B ^���=�	���(�׍��8������l�/f:S�i�Q��.�^�,�����&���tڍ{B����a��኉�,�l�{ m��zFG/��?�"o�0鮌�V��b6�7���^z$9xCǶ�L-4z��3�Vx�1=��K���]�mF� ��DW��}�q��H<��v}�D?k�h��V������e��uEнDj�]�˯�T�����O�
.���穣�:~�'����ޤxW#D�)-E�2��_h��&MA\�L
�-ⵎGCMzc9R�Ԋ���^��g+ܱn�oKnD�V����~ָ i�.x=������uC>��4#�s��m�꧜n'�|cR�$��6�1�$YsJ��
�zJ��W��z|�v��iӺ�Sɂ��!c3���_��!K����A��@�hQT�#��E�`O���H���σ� �_4�!�7zhh�����}f$�dP	��6�h�c��F0ڀ�C,�Ȕfګ�$!3��e;6�z\Vc@��#�����7�@Z�˃2{V���B�ȕ2��W � E( �Ғ���(���9d��}�������]���i�Qb�:]2����t��I&��y�����VU��՛�@g�T!���i�a �m�$<=�XXo�O7�\s$��!L!f��]w���"O��5�� �9�u3/���V���	���`�~�����3G_�J&�ޏ0�kf�6w�۪B�_0]&��e��k�XC�1������j����3��5j6�-�����t��/xZ햎�C8;���?�>��ڡ<�]�"X��R'���I8ԑ����u���7�AP��ڢ!`O� Rtc����Hmo��t���Xf2O��J��5r�3���Ÿ�(����)�S��2MA���.�G.8��J���n*����o���ZT��d�p�����:,��Ji�n���4]�M
顥8�u�'$�3T}D��yw������(�����i�2ޠ�%|���v�q����5���cwP��^�]Q#���s:R�m#�D>�)=�e�r�y�}R�t���	��i���MR�H^��ށ1N� ��&�;~�w�p}z�x��$MqI��8g��D/�6�9$�EO^�y]6�%Rؘ0��$�tI�r3_:9gV�pIH�/�GB���H,L�ѡ�o^WM�p�݀��rx��6�6̆=V��;1"�ߐ�u��y-b��浓��}��Ԣ�8�:���ꥡ	�a;���Ӌ&��ԓ%V=9B�h;�(jCn�77k'����h#�;��<�O�[��[���>�"�Y�ӄL=��h����n��2)d���ǣ����k�`��*��uKg?:�^����GK�A��I��`2p�H�qd�`1����}|gce�B�i4��K�{[k&E���Q�����%k6��Mk�<�5TG}�vr"�L�+�*
m/5Ґ�"F ėOr�w��bƏ�K����e̶�-U�EԸv*P]��"�
�6G&Gayϐ%�� ���^[T��}�wA�4	g����n��~��?��Uт���
Fx��J��7��׻�07s?�@�V���!N2nA"Α�'��l�HC��uvY+Ū�ǒ��Ŕ���4r��u�ww��ӠxӁ��X�{Y�C�U4_�DF���ēӧ.����f�	�yK>� sH���`8ej��܈�Q�����V���f����8H@i�S���I�X׆��Ɍ�%��3���T??�F��d`+H��M���3�<�j+8)����&�v̘�)9�x���HK��
b�e��/�g�@�K�����>;ү�����������@��E+�>��Q����]�E����"�6�7�$����� 3[㩗�"xY�[Z띂�~��:��R��!�j)^9L�D�5h�p�_�>��DJ-�˚$�,��F����pXu�~�g�����wK+0�a�2u}���;��W�f)XY���3�t�=6�Ī����U2t�a�v�\&�;VS�A�0@��v������YκSRz�������<��&�����
���o�e�2+�!���A��!��K����I���CQ�5��+�g!�%F������!���q�?7�*JoQ��j�# q��L�>A�q���ݷ>k!�������ӜE�/��(-�@F�Dh�6$��μ�͟J���Y�SʾbE�x��"_! ]�߱'�`f�sjwK(;IS�뀤�(4�w��|�z2�O.H���$�+.����*ɵ���}+���$Kb�]I�(�P��r�T�4�Л�ru�Q��C���Q�tSg�\~���!����$�NW>�H̹s���?6���H�k'�bX�ԘR�q�z5�"#1c@�ծٮ�0�fԤŇam�4�|���H�o�e2_�%�{-��iLK�c�p%.�r����g�(5����9U�����Ox����^�����Oo��C�zA�8Ya�,_��^���DP4��F�mvC�g���݉,���kᬋ'�7'\_[F#�ȻA��8_O;��O�9@)��1osB��Xñ��q�f�׈����B6`g�qQjg8'������>00>��\����0H��`��Ҷ�sL�3��B�>Ҟ���r$� �������um;��-5!l��D�V`��^I(	C���ӎs�~h�q���ɩ�Vg �H���2�ӛ��m����\B$T&�ȹ��b�+Ш ��.�m�vY���51��.
5!#r��D�[����!��+�h�m�Q�B!ɜE]]��~�� �]r	�?��'W9Jo�ww��ձ}�t��)X����{���M��@��zm^���_S6P��+!DB%�8&7*����G��IiL#l��,