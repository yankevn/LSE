��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��c~��#�|G�R�~��䣟�"���g��k7�����b8ƻ�a�2���S����%�ۋ��3����|�rV�g��F��[�%�d�N/W�'��##pv��n��y�8B��C�|A(��N�z��?� �JG_֕pkD�&nS./Ђ!Yl>�eȟ�ơ�ʦk'�S|`�'ޜ5�SQ�^C��ֹ��>�FV��)��_Q-i�Fo��H^=���%���O{�k⩳��{��%q?�]��Fl6')�gp�q�H�%^��9��iУwb���kj������G�@�n��`T�V]?NH��b�$tAl��;`��ق��emj�!�&��yk	����U����a������(�&�g�HҐb�=u�\�� ���A�dsxu�ɶE\��*F��!++6���Cc�8K��ۜ'��#�F���O"��w�i {߂�1�����L��D{g�{ϴ�39��؝/��ș�
��%��LT�P�����W�5��e~@�.YF$(ӫF�,^���c����,��>p]Z�~��h�'�c`M�#�TS����~��Ӵ,�+��e�e9@���U�4��RWr�gA&�����.�y.l83��"H�,��4��$1L���;�+B3�ލ~�q��t��Q��?��9k�4�16�E,�ǒ�Tcv�~�F���}Y֗G�#}20];�����.Q��feHR���.�!-[��a�{�xݭz�1�����?���2�Ď�����"`"4��`W��2�i�3J��a��9߉R:[�en�/�S<!�߁��g�.D���#��� S�0�Q��(�Q$d&{��(�p�9��`���!�	
DL\M}��97<���� vi���캹�>�l�4ɕ%&��$.(q�TZ�~j٦F����R�4� ��=(�Lxa!��ekGy��8���*�����7��Q�mUB������EM��D��+R$.z��7l㪓z�M���RMG��Q �G,v����c��N/k$�j��:��^�5��c�������)Y=��>�w��M&��B��
�˨�Mm��hԐ���^��9i�R4[ֻ]J��;�sv�O?@���z�m��/�Y�$hR�(g�wֲ��T�A;�q7�y��0��(0pa�H2�Kh�c����|��)
���/�m\���/�R�-�I�,��v{�M���*�ǺQ�Z�3��/��O|hr쁒�1-7�1���PT,�~VDӇ�s"���;_�_=Zr�_�P��_yT*J���|�����ji�-�I��a����,6����.���7[~*�� �b.���4�E�~�n�d�YY&~Z��C.���QN��E
�O�*:a�`�#���?S^�z�\פ�ȅ7�c�}�1�Z5�@�_"+���r�_N*�6��v�-�� ��������+*��Po|ܿ[������H7p�OYB!|��XK�� �J,;��NNT�'���EFc�~�@����-�FLw����3��1�4f�g��H���n�M[s�@�PC���gF_%夙�K��ȁ���Š���	k��5~��/�b�$S�����3�7�|����L��f�����b�ODpt��ËA��� ����<��8��r�;��TM�#x9�����&	�9��,��񙚙�a
k���L����kQ툴��ۍ��]|Ŕ����4n�~�-{����Y�~�+�����JqB��6�	�L6����Ь��q�.n��B!�8s��3-�����/��z��I��t�p�"������CXC̐���Oϴ	U� �%�2����	��N����~8�C��!�]�5̵b���d�͆���,@[�Q#B���<�����v��ʧJ�1oQX�l�;�p8ޤ�ť��e��F��$[���CW��Y;{ ���a�����B��� 2j�:��:{����Wq���yM<\�&
����+�)��ȸS
ŧb��i��S�oM���%�l|�Lc�ts���&�[�!�v�c*A�n��m��XFү�{A�;%t/'�Q;v�ڕ�S����ҹ鼼���WU�%��uQ5:=;J��?�N�}�N{|��c�?�)¼�
NJ[��;M�ipc����:[>��R��e��_vO���NT��ϵ��E���T]}�죐3ߒ7�mV��ࡇs(v�*6kt�Z�h}^Q�e2۟�� �ikg	A��� ��x۱*�)��ݻ���@!S�4^6�_CP��H�6xB}K�
}�,ɘLacN�.	e�_����y�3�+�t�w6!bdI�#^��+E;S��+7�@T�q���-���fV*�y� 3���@�6&*���$�v^��Q�B�8���~fL��R74(U�1�p��S��fxĚ�C�N.��L"�D� �~?G�b��h�t�i������@{��~�gC�u�f��L*�~�a�t��_�L'
"�܃�o?����Ǉ��Qz�$yOv�T��-e3���NK���i�����u�f�M<������&��2�7hޠ�6���
�*ܸ�CyNG\*�w��!!Q�0#9D��e��>X��e��L���� C�Ř�i�k��O��/\��{/}����r�SbA����{m�1�)�c�#&���դ�s�'ſY.��f\�9T�g��$*�Ô��	�)nV(�0�}a|�WFK���)��ׄ��؄�N�A�Y2<��4ɒK~|!�����jE`	��J)� �߷2�8/Tq���0 x��T��N�Cu����T�2�_��o��d�������)����pa[g��x^�c
 8��Kl(��dU6V��8Ze��_<!RP@b�z�0��K̭����cF�7!���Y�E�wX''���8� ����|3��*�⥎������m9~ �ǋ3��~~��s�Fr��^�Wl�>7y��L?�p��l���l�=��#'G�����2�Pb����ְ�iqF���:�k2/d�Z��3�ܦW*�T�X(��z�&�yI�;�!�
�]ށW�1�EPU�.u+t8S)�-x����\1�$mH�t|"���{P�6F	�"� q�Is3��g%�l{{\���y@nct҇P��9�%���U	������JmD�쳬��;Kk��,E]�ț}�"�`�>�"�ܪ۞]wwQO�ɣ>��5m�fq(�jJ>�:��vB?�G3{��}h�R �ք���C�����af�+�D��,��|4���4�0aߴ�� �Ž���ɷ?M�4�U�ZTXLI�L#�j]懿�I�[E�_β威���\�SD7{�F�4�q��ȑq�Y�z~5�!�H��o�_������r# ����
��� ���A��M'��a����6/N����:d2ǘ��ʖ~��߯�r9� GMmc�5ȳ/v�҄��4�S/���5�����`Q?�1��:�uҍ~8YѳY I�|	z�M��G�/��D!�N]b��N�w0MLJa3�����BMd+@��z��;fR@�m���}����,~�����@+��L�^�ѐr�|h�90sKd�df�����Դ��` }P�������o/s}7t}{��J�kn���UZ����o��E�z��O�ٕ�|`z��U�B�˕.��cK6�U]]���#SR���E��GBǤ]�+�8��3��dن]�'�d�WW�vu�5�'�w!f{_��P��^�$v �yX�#���Hqs�]�	���5L�ÿ�Akc�F]����}��П��K�X_�.�����-�V��'(���SW�m`�˩vA����C�얃	´�_Ә�~�X�P�l���>}S�#�HX���;�4���� 9�����V�F ��Fj㾯I5���1�i�>�EۃS�����=�8�����0�J� ��/g���阋bg��i��틋��:C�"���iZ�3J,�v7q��	RdZ6�k4����q��G-}�-!q�ꗓ��ǂ������.�LP���S����4���ę����rL���&T��u%�#~��&0s9"h�x����ٺ5��8��ux���ی��Ѝ8T��'�j5�V�E7�G_��݁�XfWXZ>t.���n��XaV�D��o�=`a̯�f�w(�H۵(�V�<�':�����E�go���,���v~d����d1j�d��V_�DFϒV��-&J������*�N�#�!�=?
f�i������ \������+䊹m]硨�}}зi.�ro3�!�2x�uM95l���ǀ%..�����+&����J��Eˡ��Kc2pM���u@��t��/ɘ>~��^�����	$T��V�ctg���	�2�.m���eEz���,_�5G�W��W������K�!w���iEWy�˚�>�'�=���p���%m�7G�E%���qw�/��/9�50+�zq�gg�4��X�~����D�����hW��i��<k|�����nv���0���,Hõ����x+��U����
$fE��/gm4^d%.Ч8����Xu0�$�h��;���b�,X�����œ7�E���F���V?�2�!U�
�x�iٵ3S�y!<�b���96Cd��v.=���3��t���x���	�I�.�E7gX��x/��:U�;)//���&�o6�aJ.Qb��<�~�<u�������1j��i�(����˧ɶ$g�<X��@<�a���� H�!�8�uSc��Ek�?���T͋x��Y	''#��AaȻ-��*��_��xezF�,0E�>$�2M��X�������O0�Uh�0�����m�Y�v�	�+�����X����������Tj��d	Ɍ�74����}K�>��W��ǉ�V�~+YK���Y��O����YBp5�8��q??ie���8����w:2e7��1rr�]Lٸd�+�e���:�5?�(����1�b�	��Edn9����6M[V_hJ���ZA;�� ��V�7�f��I���U(��y� ��p��]&%���0E�yxJ�����N#]_� ;��:y�n[w��J7
0Bj7jp		�r}�j�ڌF��y���{y�9����� �﫪��1�����]w i���¤��m�jaA��<[0ILΖ��g1�d^b̅;�ӊ�$H���X�-�+�*k��a.I�N��?�MĂM�'�m�'3�>���D2/��~�BN��W���s�����dn���D�b�ϒ^�������쥁7�O<�(�� /o�+�0o���}ðn�������i�x��@�_E�Ԫ�V���O�4I�������|�[Yؕ�'I�V�����h9�%%���~���m��R�B�ڗ�6tZ[���tb-�{�����Ҿ-}�^�$��a;�W���M�d9�0�L�F7���-E��z��M�uZ�R�D�������vR��Qg���e����O[s����!v��F1A޺����W����E��[	\w��q�G����+8J���(Q�T$h4O�Y��~r��t��)!8�vt!i��Q�t`����X��'\�}��(��d!�4��&��#`r�Q�	M�iRy2�.A�~r6v��U��D���h㬝��024�2D>�E�A �i�YA��q��g����7�-�1z��xA�LBR}a�x�S
,~��)����5��)h\�K��&h�y�-�r�R�����ޜ��w��q�)F��x�0u��q����cM�je��-�ޝi�+X�Φ��i�ZAO���I
T_.�%ype4����
�C�x���cl���e*@nm���Ԫq��� �n��Ř@�X($qO<
��E���؎�X�{&��L_"��e�_��n'w�;�h={a�6����ܔ�[�5.��?~��Xz5jf�Y�E(���-���3Y�]���������gPꂘ�=��V����/f�_ݥc{��@f�o���|3��n�L:�6b��ϫ1�4WD5���*�0�`�ߗ�1)�I�.�/~������|YP��!ʼy��g�~�����)��c�ntҝc	���PֿOSS�L6D����O���d/(�X����aY����2�S���j�t����AU����o�[��*ģ)�H�;Kn����=�¿��9��|�Usr�����Hم�L�}�(`�_���}�Q?m�Ecr�MV�K��4�ol������kIa�`�%���7y��p���ו�)�+s��a�y���G�x[LO+�^�)LU���9!q����5:UT�B�X�p��l�:�y���8;ո�%$��U-iB�n҈�3����]b�rK	���	�[+��K�TK�j���t��/bƎ+Q�+�-}l�ef�~�w�5`Q"�1�E_�SQ�(��[ V��P]�acq#ȏ���3Y���@��7�]���HÊXr/����廭b��I�p�_� ]�P�\x�)����ҭ��H�����0v�KҶ%��|�]���r^�F��*g��d�/�5�Z��Le��Ҕ��3����Ul���Mă���J�z+M�? u��EQ`�F�n��Y���(:8!�`�uX*��߄ �Q"���M�I��N3�H ���NK�����ɪ�V�f�֢lD�Ux��9�(3<�ED��;-^��[/E65��Ū���I\ݤe^U�~��Ym;���@4*����F���
_��,��D�#�̀�$�䭉I�]o�`ۈ�w�o:P�Ҋ )�d��

�ωV/��i�i��Y5g�� ( �ۊ���e�.m�X�m�ph�6�c��gd�ySz��[sΌ�@�t���#�+jG.��� U�;�G7���^���T��8C��@!\�[��R���,5)T5f9��J�a@kJ�G`���c��(W	?e��X2�>�?�-G�RU"��|`AE�p�!E�A�e�B�"ܷ���j)�ѕu����XL���9��1Ǆd�K�T���@�o#,'G�9a0��R�)��a"��mDHF���=�^�&�;�zX���V�%�q9H��S����-Y�����f�+p�}O�j`1f���n��G�W�E�q���J�1U����'t؏�΄�ee3
�=�n��U����������;d���, �&;��?Y�VP؄�ݶ?� m�E���X�E�����?<>�1}�P_��e}���{g7��+YBbYC�*az��=�sV/��<�zI\dt޽������$��[d�*zSj��W�k��|if��"Ђ%�`�~�`���E��_����I�K}��� ֖���gW��?F&[	Kߪ�ڝlM�:�	
��Gx8�ï:j�J8j*�@�E�g^�����5$�ӳ$�7�*"���n�V�?�L�sS�o�,�� ���b��q�)��d�s��'/2;��x�Q��f�n|����?A#��ڐGo�E~#PP�]c9l�,���q�N��!����3(Pz�W��:��&��5eR2�si�+�n�BL*O\��S���J��xY|��{ݏ|	*��MRIW��bq]i���m��.k�i{�� ��"�ש�����ɳ]�Q1*h���E0�=N�B9Tf1��d�0F�1iu2�,�����vQ5_�I���G���t3��N;��I�I"�W&�jRЙ<�*�r�n�X`%17e��"A�L�l��;򎂆&����h���K�W"�^��H�*�Ia�@�R\�CB�޵�l���gQ?�Iʜ:��3�Kx~9�-����/�i��V��h#
���P�l��J��K����ιm0?�����&��C�<��co�-��?�;(ힱ
eX�A���7R.*H׈-G���L�55N+����LE2E*;��EVK�/�E96����ِ��^cu
�r˧U�4]֐i�\*���o���D�uB���+l�������2}D�ԟ e��"	�*�{�i�H8@���� @u���J� ɫ��"Hs�͆�\�H��S�kč`�b)�lq������H��I����t�8��V!^)Icq,"K+Tx������� ���K�y�� �؃�#�X�;X�n2�{��CߍX�|��/�1f�.|�(`u]j��0k?.�\;���:4�o3F��wTK�{�\����t�}�Q�蒜,�(]����XWy8��C�Qڔ�}��n��+�<�ʊRF�!1��T�6�l��̏ޭ��'�<�M|��ȶ\�#�-ĉ���8�H��9�YwV�����@7>v�A��ӈ�+`䳞dڭ���~R>@�E� ����d�)�Z_ 0�}�c�P*p{�p�����jк��sل!�@��Kϯ�)!J%��3�tS���k�y�G�/�Da����ws��*��!������~�����O���-����3��8�@0qy,��;����G ����n�Q����5'7�w�Wr4�;��n���YY�+�m�Ty�9UT!�HoV'h��#��
�Q��ml<� ���9�g�|h1̃�,���%/��n�x`���4yРW%��'Q��e<H*ߕ�}�?�-�ۚ`E�*QŌ`S��Uc�8tf`'"/\6I��I=z���ձ
p�V6H
��`� �u:���g�!ƬDX�!�ZJ˥�|ᓔ``CS���H|�R_��8�w��.8��8���`aD��}��1l�0�ZED�$�l��b�"�~��˶�2^g�H�?�2���P{��*Oİ5X�(y���"+o����E�#T�(���>{"����e��sl�����=+�6N�2� �Ͻ��f�̶a�:�~���[.֝�����ףah��?��V����ANl���ɼ:R�n�i�yŦ��،z�s1�&��X3��6�v����vm���+Z��Y��T��$�P8	�pU���Ub�B�A��0�QK���n� �=���y�w<22g��-`Ɠ���?�òL�AK�����5>�ۺ��F"ܤ��r�qa^I>�������>cLɴ���H�ӖxB��H(�C�>�Sp�U�y�sa?�c����6}����ZX���FJ�l���������������I�e}� �&��K��~7BX��� ��L��ȵ�U0���@	AF��y�8C�ϔ�k���C�1<�԰��c��Rɵ����jL�M�G
�3��ޓ��Z���U`��je�BZ�RR�{M�[��{��E
���U��;��N�u���Ip��n#������ۏN0�B_���fz�ݦH�H�pȔ�sK_�� 徭��� [a^o$�zJ���3o�����q����$@�>��%!��&Tꂳ[�2����2&SNY��5��֓O�]uâX�"#�gVp��%��P�|zcl��2���%�H��7IG���vG�Ǜ�UN��_j��+��gM%6v�pw�/��A4���0�Xr�n&�RROh���4��]q�ݴ�(Tc�p�^�]���.o�Bd-�:EM`U�*M��T��]��͍��4d�x��Ke����c�G�6�N��̈́�>���\Ѿkv%1�A��[C~pҜ~�S���o=�����z���p�g�L�9�4�o��r�m�x	%=�
�/���:a�D�^����4��OZ4{�8��w�~�C�_���=���n~��V�=�%_RY�{m�I�6�]zp��FQ�����Tw?L����M}�=� j�ܨ�;�Q�n��r�{�s��~;072A	��;|DL	����΄A�ʵ1��	8&���=������6�S��>�S4�sojx���g<��G���8�E�0�`)	���7�/7���+�˱"�M5'J�զֳ��\'4�Q�� s5朦��8��r�m���6Ԓ��)^M�y�|�)-*%��(���W^�n)��A�|�j��h��K�	Ή��c�Iv��L����x�疻�,�,!�>�� �C��ΕP~W������OGO4�]���i:�3����=��ue���� �^8ۈ����C#}8���D�u��\b;SM-.&����668���RN1'��&�����v�	u��-�A�.� �e�0H^r{J��C����&lݤI��$U2���!��Ac;����L��u o��W?�)چ�}�#~�� p��H����'�����~;#�ф-��;��롾�A���y�!��ti�4���N����$>%t�4%AT��K�Y�9��(.��;��9���lF{94z�u�Y D��&����o���������_3�hdh墾Q9���3��nt�F
�.t������C��S�����v]��INPu���z���p���A�RSP�]�ƛ4����.E�� S�v��Q���QJ�+������A�*�E��P�X��HJ��ƾ��F.�vW=��rP���9,}���o�!`�;�#�7h��Ϯp����P;w����._��/`�n�?~~�x#�H)�����g_�;���PS��zػ�sK������U�f�%H�,�����t�\[��G���,�6=�H��>���'�/kD �s3�������yL��:4͏��j���9��ڶΛ�c«�Ɖ�W#���B缐̠\��?s��r�!��R���ٞ�E����Ny�]@�n+Q^�F2`E*�d���A�}R5$���&����F���M�~�<Y	?� _�*�s.?$e���N"B��%�����K��;�CdG!�9n��ιA�E[���A�43}�\$6�n ��@�e�4V�+�+h��E����F�ϼ Q|$�Z ,L�`e1SV�@�B����o�+jϢ�N�r3��!�\>!Vzόß��^X`YbZ!h��t�����{�f�:�._��oU�ٖ2��̴Ji�/���Q��W����?1A�ҏ#�����wqπQ����}�x��ȰR��*C�~�+J�J��V2y��|��
�T��gFw�F�.�r C�dsD�w�0�څ��G����[#��*��gX}��VFQ$'p���Tf_�.����מѳ�iM��^���q���C�-X�h�e$�#zzs�j� ���I���{��B��T̩!���L�u�x�WJ�%R�(�7�3�l�[1�e�x�%"�
� b���c��d��'���)�=�����Qi�R�Y�a
��Ies��&ClĮ���W"31<H�|�X����{��� ��)!�MU��,�t�݁�"���/��I����Ǡ���K��j�";�ב���X>jS`���s:n6��8'�Bs��Ø̉�U����:�xNc����[�|��.�6�����X/��F���Z�7Ʊ��k� |��t��<y��͊F��/�ű���~�n� K0����<���9Q?��E���s`�%�D_�/��K���h�ǿ�}�A<>����=2�ɶ|7f�qde����K��]0%),YU�I�ܟ�ޑcnC�\�\�᯾����:?n����=��Og����џ�����ڒ�~����u*��D��"`��ഖ)��?�I�͆��I��?��2Ft�����#���{�o����\$*����[�S�׀�I���ϖ�f��#�cL�LQ���m9��H�6�%���	�<��W���x�r3~��IJ�p;x��,��s���ի�(��)io8�vTR֘Q��I坔ؒs��ݦJ�%ކ�GS��p̺��}�k��Տ	��1F�S�5+l�k�#�b,E��{{\�G�L\T�&��P�H��t�e��v�0~��2F��-�~Hj"��"�@L��c�W�мA�䓞l���[�ZrX9������~�{h�J��'3$=�@��x5tp��@^���\ے4�J�7���$-9��{֋���T'�TDQ��U�F��^u����3��Ӈ��l���T�S!d�$Q�y!`p�Iz��!)��8���+���E	{������P̗ o�?�Op��H��'<�=;� �Km ;��E�
�o��s�6`K.7�MxZ{�®$N�x�Y�Rdxq���S���M�"��>�����'����c�Ҁ�U�2�d�I��=�6���x��Aw�e��*��A�,�]I� �Hw��q��F1���"��?�?G�hY�^�PCE9�?<�U�׶����W��Ɛm��?��_x=�`' �ט��G��*�r�ݟQw�G-�U�S�r�о3l��e�c��Ԣ�&�B�����Z�&ʥ�Wi���h�<dB�w/�n�O���,�K@��i�ͩ����w.��C�2�Xc��9�� \�;�+
lbQ���W���8�����6� �eg�9>��B�7����^�]�Z�uNs�rYs���{��r�#o!�Qo���⿲R����ǁ����=j��+�8�q���2�{�I I�ES��~C'�?X�ƿ��'5b�!�9��8�k���Ɍ�T���9 �( ���i<5�#�)%�q�N��QY��y^����i����0��.�^�
���-�D�Ց����
Nk7�+�$-��{�Yyx��^����]}�1�~���gr'�K��_�"�ݷ�P��bp[��r����EݪR�
�:�=�!�z� �ofZ	|R���U���A=�X8à��jy���)�y!�KlB}_	�m����"G��u�	/[��Z�v�s͇�U������zRI%�gG
���h��S�a"�laa���y~~A��Էx%%��%�H�)[,��>�ڼ�C��7l��Y�S��j蠠�P7''~��w�ѡܾ�F¤�T�Po�~����h��H�=���%�Q ���b��y��,%�%>��x�=�8Ƥl�׊a���E`\�ӭ�
r;���r�L��n)��fb~�|:�!�(Qb���	��x|u�>�`?����H�_��8�M�l���cn��J�v��t�tZ��6��'d�
]��ģ����ҾM�W�f5ڈ���"s�*UM~
��� ���E�$�q�{X�,�0����{˚�1�9���[u�O���iX���Y%%�vLV ��2��ɴk6x��W_��������S���������v�Q�m��d��K-B'ŜQB}��g�$�e1R�SH����5�,�r�g����i����BUrc����.�{%�%���6����(��Ȏ�n��(����-i�ES�����c�t�c�6�Ġ�*�'�}�"q=����E����^SUd�S,�C��_�Lu_5��?���;�ٌ���E������E�F��u�ε���k����V�i;!Y��c�ѡDC�ssS���A=�%6��V,��j���<:e}U�����NP�������a;���hz�r���%�0�M�HWܬ�Qvi���\��gҵ�1�2��h�$z��X2w��4V$R�|���S��s#8c�m�����z���eW�S杦: �����r~�H��Hޑ$��H��3�ލ*&[-|,J�:��,ԭ)襑�ŵ��V'��S<+K��\��j�B�69s�
��Z�q��<�F�J&�hFԢ�F����l���]�0�&₃%�Z%徔�7�2À����urt��������OJ��6����5�f�; j�~��t2O]usG��E&Ir>������+��	d��l�;��y�"[H����#"mhاC���L�_R�m�2&I>�f&�!�ƽA�|(��o�Cc{*�Sg��j샂J�n%	BD�"�(��d�L�2���A�b]��J���Jk������}��[@$�+��]�jq�4�y�y�vY������7'�j՘�b�B��j�GePńsL�}�x��>�&`�饧c�6����1OT�M�}C̩�F��q��_n���A�Pj�۴�+k��]Ou�[J U���tѝ���0��ٲ+�cw+_��XN��_wm��W��c@��y�4��d�CiIFs��*���$����,��3���?�"g w2K� ��}\z��E?��.���m�2x�F!�-�	[B�0D�/L����=K�*�$�_5��jJr>�l����b�?�X�dz��d��Mc��9(��k���4h����^A��m�%o�'����K�":��V�/S0uLYwG�����,8ߢPQ�
h`E>!���V��y&�ک�H�Qc#����ę�7@���=(�:����}%|��l�3���c���c_2�K�$3�ώ�H��G� �c *4&u��9Ki�u,�R� �$�F��?�U#0H��wK�h�������*6�]�|$g�hG)o�`;+����A�>����2;�3ՀOe��J�I(���lsކ��qB+����"��-�ψ瀆ny�AI�S����]�LA�mC��Z��z����K�Lkh�~/����Q?��=�m��ڭ}+�س%��C&�J�>Ά�(����ݑ=+Cŏ`��BY��c|k�<�=��g;<1��ERĀ��CMՄ��Ļh�a)"`����������kE��F�*qm1�>V�JC�}I�!���O��[���%9F�/�YJ<���� �[=JLZ9.�Kp�R��E=,k��?�l#��@,E�Q��ΫA��LTa�Άݒ	�ո�K��o�hUeIƁ��ݹ�4��9���L��j^��fe�����m/��bI���C]K��,�=y"���U��0�fZ�o9'x��-��"���a�D�/`=�1'&srt@<T 5&uƀJ���8oϴ��1\�ҹ��X�]�@~~.hL�t�)��9@}㧕'u�*�Ak�T��tG�8JذD�E����~�-���wJ�1sYx.0DA;O\�9}��iK��q�Vs��j����Pn�`���M��B�Y4P�R�����&��Z�5��o���r<����ŗ9WՕ�i���}t������錓ϝa�~̎�_S߉��.��b�`җw�n�¨��A����1r��1�&�B�9]�q���#h-������OE�Q��B����'��)y1z6+��l�H��>W��fޒv�P�����
63qZ	^���3��+�� ��ضE���ʣ�S2$��@�o�8'L���,cG�� O�/��H��&�z�NnSb�v_)��̧�\�L�l�柡ME�<���x ������"�6�?���6��/�i����5q�^R���d���z3�Q[w��wʦ��,䂶��X�R�	�	��J�+�v��3��U֮��,:�R�� �5�&��ZM�ܻHp����Q���n��8�ey>qVokN[NS�p~lhO�����񃡂s��������np�s���"���k����K�H��݉↩�A��gn�c*���̕���o�g:D�F'FŜE����b�s���e]���<�Y\а���x���3��Np=����N|�Lk���/9kJW	��N]3�
��\�e�>/Y�H��}�Q���d.���ܟӁ�E��R�ic#�O|�$҄��X�lս+ti$�Z�,a8:�p�Q�Q9��aD�*�kc��M���t��ŷ�����r���A�-J0�,}gfQ<ޗ!� ��H
�*q�~�J����)؉sU`$�\/ &f��}���N�넶?�ݧc$f�R�)z�\�{�|	R��y�X�K;	W/��N��y.�t��y�Q�9t.ձ3��9��%J����I�����Y`Nuh(NT�,q���!_晏9����|:A�Q����`F�֔,B�}3�yj�U�>l>�;�a}�����X{Q��v"���[�o�Rصhg�<��Xд$i��,��i0>��qt��kc��+`i���>�
��Rޫ���C��5��x�����$N�[5;��uQِICB$�0 Ƙ"�+f�+C(�OH�#} �48['���}jm��n�AZL��S+ƛ�������9�`��Dّ<����{D�8{ �����^dx������5�"������8H�wK�O��MS\�H�����ඔU�щ�([��9a.�I#JT��J�y�w�"	�H�$���T�I(���(���,��e�i���X��?������H�?�Tڥ�����}��j6E�Ӭbo| �\���7I_ǻ���j�L���9���Ք3�RA�帣ty�Ŭ�l��on�f|�;UNHgR�Ƹ���]�]��E��{ � >z�jY]C�2�W�}�!"
h$�1����C{Δ�|�o�����+n�A(�Nx��9<�����~���h��V�G�����Ű��!}��EY-f��(���	sݨLF���G��Ny���(}?����P��f��E\�S	�X��^���Yh�#p������Y�9�O6�0�	�ޑl;.��ؚ,0�N��Xm���&n֞eE����S~���b`\F�����aw�U���A��"�\���®x�M*���f�tժ.�y�5bߣٖ3˩0F�QWx}��Yʣ��J��h��i��I��BYҢ(�7X����r���4�h�|'٥��F�)�j3&h[6 4����������<�|AP�����g#�ǌ`��6�7/��0����gOl�嵟�R��~�?J�M���:Pl�
S ,cg"���q�8l�&8�N��t� ��4H�G��ǫ^�}@G�%�d���{��w���t��1���x��m2�ݷ2��*3���7��;�ԩy.�t%%��s�Gl_;Dh w�/�n���m�c��u������xJ�߈�,�V������k���Vy�J�*��i"6:�IJ�ֵ���ZcD�L^�����pڜx��c�1xRϩ��cg�a�]UaD
��D��[�L��ì㡶��̃����D��o��Ml�Y�o�Zc�����0�0H����W���  ��
����X�Y��y��ӣ��������$w��֗�x"�_S̩ꏮ�(�i�ɜM�h���YH�cLe�;))(��`,�*KC�j�a��v�6֍1�x��E�-�&;\�jV�W�;�����$��q�Lr�Zh"A�+<��llٓ�@�����(M%�����)��-FI�?L¿
����\~�=�U�F�ʬ��{^�v�)'�JU05��F��-��W�!�.�g�3�w����`����r��)|�EΗ���g��S.�B9�`�.�hh�1yVV/43�כ��-F\mm�D���!豽�z�$-��D�j��pɖ��c�>&�a�Ь4KTa�c@�T5��vB�4�m�̵���l&xī�$ߊc�w9���-�׌C�6��4���=9��7	I£+Syƍۘ�f'��K���bD듅)����e
L��S���K������������[�r&��,�d�W�v+�K�3�"d�:_p�%x+6BKі��]�;�?Q�l�Q�7}y!s��LE�}�;A������L�>�6�����p)ޚ��9�:��2�!ϙ�.q�c깧��ʗsM�"K�+X�ñ���W��F�R^��F@J܉oET��%h:L�����Wk�K؂'Ӽ�#+��X�v�Mf���)�K�i�oO�O9>rP�`>1��{�ܦ���aq��`DG��)�NÌ�v�}H"Ѭ�&KՃ%�Ax��0k��Y.�À-@��6<���7g�ݠ�g{,J��QY&ܯ�A��=���ǰ��tI�h��g~�ן�-3�[���gbrݪSw�T6K͏uӆ�%��qt;�����<=�6�H#��ތ����=\ϔ�����|�9���j�����w�ۤ������A���F��m���"8:��j�8�8�R�oK0���%t�)fB�ޡ'��J��Ru����g:�z@B�ژ����V�QJJ�Ns�sSx���b�=,�������jd�p�F�<�浗�����?����±�����*��و��w����H�9欧4A���"
��F�xu�9`ϐ+��\�󱑣t��x�s$�&O"в��uºA��.oD~!�Py�E�f��&\��(MQ䲋8E��ܿ�7��0	�6��c��g]k�2��J�H<��4��<���M���8��K9�!�$�"j�JQ�ܣǰ�߲݉�"�A+^�Fjn{|Iʛ��7�-����|�hm�n���辸<b�|"ŖA���X
�d�5�a����c����Gon%��eWh�kZ@M�E��4t��� �����~ùύ̬�ͮ.^<��#������q��I����cz�^����X�B�sŏ^�`7}	�V�N� ���ٕ�CH�m��k��n�`?��&C�g�傡����uH:Y��g�&�|8��@��8<F�HMJ �ޅ��1�4���1K��X���k^Ʋ̏�mdާ�F�	�]�!Ś�"�8��)w���!��mȇ*Pg$���(�J��GcG2n���i��(=a��:20�����%�f��Ώ��+��[��X 0�:��w�׌HR6g�m8���O��^?$�G9���,rct.Nx6��0y=�P=���:fU-MIu��f3��WC���6�`�]������C�ú*���R��nVFl�C�#X��x�˗�1{�L�Ė+4���L�/ �W���F���D82��'H�%Y�r��qu@��W�SV�n�g��`Ǜ���)y�}J����wT�Pщ�|R�y��i��R���� ��c��
?�-Nh��X���%���!�%�j�>H���\��`�K�����U��=6�P3F,��>C�.~�Y�%_��9���@R�K����J� A��s�"S�j���՘+^
��\L�&��i�S��X9!C
�7	�X5�_k���
�@�d7�JJLZ3e~����C�ƕdm}Ǝ���u��3n[ &{��>��[�2Ċ��nH��C�0/��N��S�J����ĩ6��-H���ϧ���"�������ec��&d�p*7�V��o�y�`'xP��@*��.&J$O�&�+��$�ryF�>�!ʛǔ�Ёi1:CU���і���*p�y��+aE���c�$E���&�5�:y���J�G�>�>�$��uvW�ɲu���T��F��Z���w��l.�vT�q$��uB����9-�_-��d��9�^q��@HP��P�V|C_�]u���@�'ĖbJ�2bvf�C�����m((��=@7�V�,���7��7����8�Ħ�8��s1+I��2�/����T����_���IM	U A�Og9��F�O�$K��8?��M���hq����N�|��Dy\=:}wl�o�U�#V�����5��8�G|�S����ҍ�&���l�o�ϼ~vS�Ë<�`����C����@D8�Mh�q	�V�'x�9���*Q�T������q`�R���\e��iYlW�Kk5�8}	��d�L��P�F�� F��$�H-u
�4vO�~@/�މ�i���0�j[�&c�Ý��Y�Yr�y��;D��eP��N���{<�3�ɿ����<'�ӣ���wq�*q/UX\b� q�>;���l���!{���'�t<Wz]��U�W�?>�`ɦ�kئ��h�"S�[�[Cn%;�����
Q'|;ޘ�i�Pq���$�5�ء<K1 L�J3�=)OM&İW��wPu�U�NEEj�i�+���p\G��b	5-q�rY�H�R�I���Sׯ�>~m��eLK�?pc����jze�������Oh����k�/��́�ym�����+���?ű�� +����Z�{f��Փ��ȗ��X�Sʯq��|S�oy�>T�<zhK!��V��������? ��4Nw���=��;w�)F�8����	edM�|�:���췸C�C[����.=��z�Ħ9c�Z�8���m�C�0B� ��^�w��O�a��H���zp��@��P�Eӏ^���qN�G�fI�H���l�{��#h���m3 ��&�a�'Q�M�{�I.�֐�!�9Ih
S�N���?�M�4�0�����+�v�p��D���x��/�P7�#"\��`��N��ꜭQ���efGC�*4�~�5652�QǽZ�ש\5"�&� /�|�E~【���� s���/���3I6ҏ�8�"����fE��Y���Ԛ���S���AUg�_�^Ci5��!�`�<L�#v8*��tс$Ȓ-a�oE�'B�� ��%���Q�N�3oC�e����ξ�x{��^Y	5�+6�af_Ʌ�%����������ӆ�-Gw	;eC��M�L〖���ҭ��_�</9�A=&Њ�x��=���u�?y���ίS�M��ʁcA�(�XU~GR�(A�:5畮*�V��fl�$�cJʂv�?��=�ξ�t)�^GBI�%�-�NLJ�����n�����v&�����.V��b�rE���:��f�5�lk��]���L?����	O<�1��/���m��0��ڵ)rr�[y��=>Q��i�cā�߹9[8l�O�"k�����_�]���d�h�Fᗧn����hY�~9���Pj��_��Ϗ9��3�U��p��ɛ(�t�1�4�'C_/p��k�Y�{P�A�2CU��zU���B��o����G�*x�O[�J����Ñ]Ϻ���l�XW�,ڜ��^\�&�f�Xu����2�m�A}������]V�2ZA�Ў ��N��4<��ue��Nc+I��E<0�T{��{T����5�m��+/�m ���+$B�y��;�rT��.@�m;�����_]/̘z���c�סǎ�_��豻���$��[�A���� '[۰,��$rg� K!�A@��PL����7��38{����TT���雚.r;�s�?Pw졤q:��8f��ua!�9����T]hpا�+��O¹�#��4��r}/����yX�>b�\z��g�h!�vB[d�f32#�4���1�K�B��ƈvLd�ǂ�Ʈ�]��3�3_H��:^9�S��|#?AV$p�{0�!�X'0�&,p��ni���i�0�H��d+� �J��̵d�� �Hb��sg��[?ScM���B���m��\�C����Qr����>��u��t�ck�9��]�
m�m��,��w=5��鄬%���n�=WZ%�Hi�ra�;*���@(��|��"pY4-��϶�f�[,��P�����Z|bs+����X�����6Q��`����F����O�u��btUH�����ý�����x-/І�{��Y�L'>q+�#^|�D�v3�?Zh�fH�wP�����̆Q�my��/�Ϛ�u��~�����3K����|*�RF�v"�i=`��;��<�ߑQ��-+s��&�����Ϩ�j��F����3L\��޷1D66�B<�:�S�~�{�4��P"�$�'j-STwɵ~�
f��lXBI]6�㬓.{ ��<��{�-C�>�P�9�/�����}�.���� &����>�"���H\*�o/q�+h�7�I��`�H����`�ǋ��i>����f�+���e�{r�e�{��ʫn��HY��v�֪'6�TE�м����t<�}����,���"���]£���{\�;��t���c�s΅�aggH���Ǚ�1���U�k7����b�-�c�&W� Q��auKѷƻb��8CI]�ߍڼ{FW0��r�nН���t4���9��C�K�![³���.���<����.�#ٶ�۝|�P2%��Ë�����NJ2�}�0���8Z?Uj�.#�`�(�������t�*�ƌ0ǩeW.�=%8p��Gu^�Ɯ2�30�{n��Wo�fX<ق����q��Q%4[�N51�HH�
!luw~��5r�����XU:�.��w�;��$��x��X�Q�K�e���2Z��}u�5�]���ښXK5����J�<��-b��l����4��$VeHe����=��g#i���=b��	C�-�B;e�HF�+,9z��M�o���-�0Q?zWO��F��00`*U\���b�˓ MF����n����J��Qw���m����JDjX+�J줾�V)�[�}��X|�9Z���@iQ���W�Lz7S�(�a�+I|d��#��V?2M��GV�����\z9�茍`p����3?��zy�g{��.	Թ�]@[�[��)j�-��1=:8���[��Ma���N����]�ALO0�ְ�%�k���.�����vY��*��`)�SW�B��O��ic% =R��x�ےU�3��e�o��������x��=^�=�uu�Е1����^x�syϦ@�*V��H���z=�T4���ĎnAv�X�6ңs�	�U5��`K�84����/)��lV����	v�C��q�)��R+j`FQk؍��	�;+���;9"�M�<���3��w�62�o���R�2��C,� ��7�Jb*�D��SZ�:��d~��!Gɡ'��nt���d��>�N�gߕx����:#��ܧt���Xe����%��Z���7�W�J#�����]#�t�r�z����;?��F�}ц;\�B��l55N���ڟ#iA�M P2��QM�;ό����X�e(-e�Mqa�Q�#4���p��&���<���l�CI�t�@`�t[CNHg#q��z�������z�M�,z���ȶ&!TyG~��w��6�ôq@��;�-k��5�E���<��;}}�\�C�ٚJ�('H�D�SE5d��$Gx�$R�sro`t�������O,���/���[�X����_eQ#^�]J��X��>�Y\8A�*iIZC+������ҐO�ou�jE�(u`�#��,�8����\�R<ߨ�L��f7�TtD&k��Ƈ�Q=�.�	(����./b@ô�o7�NE
����b]�?��f?@Α6 �ЧS���ЅWc�;��E�w	Ij.t*���,R�%ΐ���D�MdG�4QR�|�����{�w	dO{�A�פ$�e]������v���\��}�߭��s���R���!�Ї��R��hPp=.v�_r��J� (�Ⱦ+�M��#2���"�._���c_:�ޒOVʃ���Ep<Otm��{�~��"�ݹ3����ǝ}���w��8[Ĩ�]�+�Ju9K&�YS�W���7_%"��[���ʛ��p80V��M�X>0����cȏ~��ܷ��m�3	��ǀ68r��u^��wmMv'le�hfq�v��᭏�N �9Y�� _��"z��v�8`�>��\�E��o1�<���1/7c8c�O?�9���(��%�}\3</ �>���Ȫ���;�I�!�YD��h�y�rʞ��� $nN"�\�,��"�M�X�������?���9�;�(��q%�hnȂ�Ŗ��!V;���9ӻ*�;���i�ѵ7�ڗn7V��J���q6.��W��Y�>X��r܁��/�i�X�ceB�~;���l�(Q���Q
���`�طB|�<�(0f�����BΕ+夹�]�k��������C�*�s��[��0�T��h�sJW���8]�!��L�f��k/|�y� 6 9�:uw����8���1�w��#�����u��c0�)C���:v��EXʨ*.~�5�3�~�iZ?#\��G"�!���\C�G;���y*
���"l�|����-)��f;�,��r>etL,;'�Y�>���CDI���6��|U����5fm�:��o�,���yl����Æ�'Q�ӈ�R\�\C�TnYfd>�Y��ɚFX��>-���d���Un�]u�oQ�Y���0WzF�P���,���C4`����!\Y`G^��0>���� 6�	Q�Q�Ẃ�J��Fgj��ա���J �A�[����t��;��2�@�L�<q�g���0`u�^��Ix�?����Ӛ+�䝸Y&��|N�Q>gu��d}��c��e��?�]A(��f�zB�`�����
��I�_�C�_���&s�n���*�� ���q�XAc@b������P�T_h�]���y޵ʏ4!*�����l�,ru9'Ɖ~���:[���y�$��C�,ꐘ#h��-A/G"��J\����Ma�Z@@%Fh�(�,�$h̵����U}6�,[�ns2esJ�Tv���L��-�\��n�8���O�3s��ZO,��;*��Υ����pN��A=����M.1�1K��y{����|I�.	]�8���0xq�d�����;�=JwWr*փԣ~����J�H�N�H�X������L���;3dbQ䈊	�%Ʀ��:��z�5�Q��a�WC6t��p��i!�:!���h��@�
hz����L��%��B!�)�H�j���.ǅ
�?�/\�q��-%?S���o�vՙ�%�:���o�J�q2ߐ	8#A���n& R+M*I��~|	��_�9�����H]��]��s�O�Q�/DqJ (� �;��u(�j��Լ��oJ>Lֹ��Rl�zQr�פ��!�ʥ��b6�[�68������Y��I;+Θ���#��z����܉��֏Y���j@�w8��ّRx�ŷ�",�Q���f�W����n �K���,.�� �s}�o�}���`�|f��A�6 s����7���]�7fi�W���B��$��9�3!��x�+��Q<YgR��� u����q� �Y�cm t��SB��B���
˽Yvt�Df�UD�Q�߭�?��-��u���%in[��n[&p����|�[��_!�Em���	�q;�<��X�����܍H/��Ty<ђ~�g�#�dw9�\��L���K��pR<�J��N T?b*�_Im���-2 �oC�m��0p$>x/�{zw�t��#�X�E����|��YLH�U���M7�"�k`�� ��:�cAIa�GX�F������k�����J�o(�ޝ�Y1x@�:`,�Tb8ʻL�K�CI4~�a��h]I�w2���2=�"ձ��숏G�����%&?����镺l�!��3k�QS���ْZ��Dr���T'!^�?��+^߻���G�r�f{
����C&�S�Eט�Mb&Q^�J;�&�+4�ܿK���DAA�
�#(6!@�'N?~@S!�lF����+,�N���'��^V}DS2�$m�b�KiaUm�'d��qA���d� =O>n��SǛ����.��WH#��'$�������Oa&6�[a�Hn'p;�>����σj�5(��G��Pڔ�9/[���(�}�w�U��`XO�g x/��o�#�Щǒ���el�`[�-�ƺ.���Z���W?�8|J>+���I�E0���J�2�4�$���K��-���tU*ƞ��WS^�
���c>*�'3f5c�-V�j��x��5��B���z����e�4Ǎ*(;��3�Z+��C�x�����'�1:�%�	�ڠ�W�W����}�Ͳ*�$}8ZS�>�y����+O�U6-�K0R$/s4�'�د'��,�Ů7y}-�W
��<'�*<�����H�O��{��r'2�/* 1�}����9ƥ����ɛ�����z�}�nއ4��{!�����!�UP��0��m��M�jXksr&�� d�<�]���G�:��Uz9���Sb�1��Һ�<S����u�s�3�XiI���GZc��JC����m"V7�X�:�<��)$Ah+�kюRX�M�m�/g�d�����^N�,���h��.Un���1m��p�J =A��R��3��Xd��QV�2;Ȼ�+���KGv����+�q�<�@jkۄ!��Q~���q�X�_�	��M&qm*4��%��c�̊�h�L��&�ݲƦAy����.�v��$⸾���R�y�� ���Q^�㶚�i����T�/͉��6�c��ߤ�R�ƴhN�K�����3��́�S+�����ڇR2�Sf�m�liW,W����y��[sݪ�\�$�I�QA��vK�~�16��5:(���MaT2)���4��_���TO撚g�6�é$�﫴T�c�Q�X��Q�Y��<[f��0��N&���%��2���x�ס<d�<5��|�4À��5$��U���f�Ҷj��%/�w��_#�φ�u����!�H+9�B���X�Tj�W���C�z}���d1<���U*��E3���'��{�������%.�$m��v�	�k���TUSh��ST�!-�H2�!��t);Z�g�č��9ez�߯�X����ܸ�䆈e�󐥽"y	��Y�$�W �>�1&��
ojR��6� ���MGqtH92<g�+�t���yR�nKB�$@,�9BT\��R9@jVa� �3@���rnLz��KV"&��he���l���ْ�J"����1j%d�b4�	���"���D$ڌ�1���j8�s�a�qA�uWD�}���(���s�j�]�(O���Z�W����~��.������V	�驒��.�`�>GM�\X!�hq��zy��y�Đ��{7�	�6����s؍��A[�6(*E���I�>1h����:��9jw��CZ���X���_�H�	�/#D����O՝D ����kpzƒ�7#��B���pۡ��U1ijǝ���͟��o�u�����ow��� �Q�2��U_u��� ���eWx\"��$X�#<<�=�[:O��-�Ӕ���9��h�5����`>�)ZF���`PնQ�q����پ{o���K�Ec�:���h�.��*����x����Խ����.1t�q!a�ĺ�66R<#o=P�b?�_�9L:�}j���s_�AY"�݇(�Ń�f�ǥ�k��6�:�7�>��l0|02V�:/4�M���l�,