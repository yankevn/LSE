��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�tڐ�!��Q�����xZ�H��V�� �]d��� ��h�hQ�/���o�~�կ>?�5�z�+|��"D�[�!#��.J �SJ�Ҕ�5�Y7�0�f[秡3ڕ4�O�~�	����u�Q�Q�H��)*��V�o���}m�'_z�8�y�@� K$E�R�5^R�Ԇk2�vv�#�80����I��JI,3)e�[�i0��ifrJ{�#{���Z6�r^V���t�1�l������ĦV�M,�ğb.t����{���6�sLk6��·�#�XOߙ�I"3fm� �G<��a˶�~�T,=��fw�s�fk����?���PmTߠĭ|d��)0�C��F2��W-V����m�7���v�n��Tzu]
��l�2���o_J@ز�"h��#-

G9�|�0w﫨/^,�w�aR^`�O�?�����JP�rִ&�Krk����ی��n"E`G����J��&l5-'|�O'G~mq�M�NN_�������8�_������~�Ur>�h�3�Zm������}��Y��Ęr0n��ޝH矣�uV--�@�1g[��ޡH������r5��nĭ��^�S�n�{Û=Pml�A~3?����W��������!�>�|-����5�xs�����Ⱦ��j�fZ�>��ŏ�yy��z�S���#������F��3�Ƕk%ce��=�(�$�=	�dT�{��O������Qv9PL13^B81=�	qPbu׶�Xb��l��:;!X�0��;����[����b§�e�/A�%W��D1��q$���L��56��窔G9�)jg�L"����[�$�Ԝ���v�D0$4��0��^5k�Q�1���N���[j!�B�CAf�hH`l���q����:�i��#��~��h.��=K�
��6�yҥ`�N/�+3��}UMHc:�`|�W#e�G�@�WjX�Pf�[�Z�>z�������?��E9VdpK";�|�e�2. a���ߍ������rtX�Pi��m�v�_j��P�>$�z�̉H0&SԦjZZ�?(RڊR����-�y  �-���Jޔ�=�s$B&3������v�+5�; Ɋ�U�;]6�ʶuL�A�Ұ:z��.?�7k�	�8x�zT�ǬR�X�r&�ʆk��^GyW��������3�WW��>�;K�g��:�V��M$4Ȓ��_�f���P�S"�����h҄���ls�ޘ`�z��	��#npף��e�ٯ�w�FĴ����1��7'�9��8�.4��כ�
OW��7%��
��<���J(��U6�r

����a�?��M?��C��X�1׳���,�kר��ժ�:�nF?�FDW��K�^����2��Q6�ۋ�5_���i�m�NOpz��e���-ߍ���^� ��7s��)����>�ˊ��s�S�ce=��pZ�+,{�O��E�ESZ��a��Q��a�� F_ځr������ʽ@�����+">�;J�GK�1@e�y�jU4��p�Ν�d��JW/����363=�|5��$}�|#Ȼo���i{{'W� ��U�b��Aub�ʾ�~(xK���Q��*|�Y8�a��S��\�/T�*��T;�}e=��Z��e��C+1����!6������¼����{N�>gxE��c׫S<��-�!"
.4�j�aܲ����D��U�w�N3��d���v�`ԛ��ȳ�
�T���}��T@9����̖.SݢXc\ԫu���b)B���7Z��W"��&���ٞ��FU��[��_*�2*���Y�^��M�<[=�)M����>N�4�P �"���Q&Y�"M�a���9����s�C��
:W�>] �κ���;L��k�2IG�lDk�䄐{p�D{az�E|�h�z,�#H~B�MJÕ/�4Z%f���zտj��O_�_�G5*���>'����
E�lA�g���R��e-Wڔ��@��G�����q
tR{��ԿU+�	#Yj��'���w!��ʵL^��['�7��$A���B���2�Bt�!P�	 �+�N]��_�� m>p� �@C��z�Ήu�o��*�����$	��'f��S7j�4���=�!0��F�yttADȚ}�R�+]��lp�zw@�I�_�+O[CS�`��F� �A��P:⃊��/�{y���Z�7�����y��h՗o˵)1hv�px��*��	{��W�M�sK(�cʓt��JwA�ѧ\m$��T`��)�@�+|�S�[��L����Ҭ6��k�(ܠ&��^��1���g��'� ��Idż�kA���O�J{�SٵU��D�Q�  y�D<�[���3S�-ޠ
|��C{�ԍ�[˲���ϩ���0����O]"L���X����ğ_Q�FN˅�{z��m���6`?���km���<�D"}�%//����u�-.i๗�%�������G�JQ�u�l���͐��R>���I�Ws��j؉ <$�M^G��ܳ)=��-jSv���j����g'sLU������k	��s3
diR��t��Q���&�;�u ���Q)������{���q��j��L���� K�x*�)�\��>A,�� 
qtp��RЍ�����=�uyį�rvc�Hj��/��3�X��3>.a9r:�f������U��8����Z!��m ��=�n��ϱb���i�z{���'l���