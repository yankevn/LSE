��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���d���kYI3���;�����J.�Y7��� ��xh�B��e[�)�xo����~uр�I���,���r��v��1=��Z�Z#U����%I p��B`μB�Dv;"����Zs��%a���Iu�p�$>>ؙF�i�x�^QZs���zǒ��F�2͝*
��c-���JzL {������Â(pZ�mAX$ȧ�FG������;P`&�o=�+����};
(Y���1�:�e�I`�Wӟ����MѤ���(����6o%�������P�CM�m����,g�`o2!Ϡ��%������^6h���ag*N�B�����H$jh����ex��*D�G�t� �1|c���}Cy���ٹaW8(�t����'"+'}E2�el֮�r�n���Q�[�Z�!R����9��s���w�Re�y̙��!J.��j�nِ�bð������k���:�-�9���F~~��6�Ϊ�%�1J�˩�:�H�� ����܎��;���VS��6 �M��p� ��}��|h\ӹZl�������d!�F0˖H���[���$��+sP7gݩ�5�_M�C-dX4�,�f�Z�S�4$�����HY(I��>����^���ɨQ����]	2�>���[�:��5���t�q���3�י\�l֍�F�b��Z��=��tP�PX|Fu�u�{o����u�^F[�R(*	�Q�	���>A`doUuwZtb�r�0���乭�QS����Ƽ�2�_�i��Zǟ�F����k�O!}���7��{����g^�j�@a�Ƶ���>y�r�k<�c�8�1��>���1�������{��O^��M'G�kkO�J�������8�F��EN��5��e�d�V`qN6-P'��s���	�i�m�"|x{��h��d"��0(��i�x0��!ݰ�#�����J���t��k;/OV�?>�B�7�b�6_�I!�}S�2��S�¼���2jL�|;��wٸRR�T�m�cL��u�����-:u��= Z�H��(Pxb4�I�\���~ȡ�!��_$Կ�䭆�'r6´�gޅ8jm\���}�2B�EI-�E�z��������n�����Jl�=�]��6���7w��k�Љ&�{��1�^1����0���U��b?����OV����������m�j�C���d��^� E���8��.�Z=�&h����L����=K>ZR_��d���PE�,����6����X <�6"(>9S�Q�\����aV���;mt 騎�+w����]�S�@ӨS��,e��"uP	7�^S!E��di���gj�&�V>4�?�����-��eX��X�%#�6�Q�C��Ɇ�ƨ�(��$�2\�a�>Wh���V�2ZhI8��w�3ÿIz(xZ�"(:G�t�(����S���ݝ5ZѴ-�-5�@a���Y���k���=�]�|�f{�f�azt*�uӕB2�,t��9��!'`��\�<jq-�3�NChy9��X��o�t����ߛ����HD�.��f%"/�ؼx4��x�n�Q}����ٖ�{�L�}�}~v����+~�S'tr��v7#}��Ӥ3�,�Q���h�v$���M{ ���Y�y�y�1��� ��O�Y4�����N���v!������Ʌ"W~��Sm ��j�����M��-�������P�(~�ڎQ #�&V+]"ƧC.FT}�ʆG�Mk�A�6i���B u?8� ߽��Nڅ�������W���{0=3׊�r�� �~Ɲc�s���#.�m�T��G�2on����<}�k�WO�|x:Y��K؋�9Ϛ=���>���'��L�w뇱'b�әc$�2W�(o�)���a�-zZ/1հ?����4c=���b{dU�ߤ�)�6��*�^�@,����(�/k�?��^<��6�+?A����+�_��'�h�6��ڷ�+�3�o��qT��bQ���N�� #,ST?f(O���裘�t�^��euw9���]�;W��xd\���1���^�l%0d�_ ���/}�ȊZ+����݉�󟻞4!vA6���	���,�һ �S�f+� �E��:Ӝ��eͯ�I�z&���S"�5g��s��n������֞SQ�:�p���tpN�-�g&H7��I�a,��g�㞞�u�X����B��W��QܩLf!K�[�9#4��q.C:޿��.�l=��]l;S�/��:�`ǝ����A�(f�UEk��$�[�be�*��l/���/��pr�+���_$fS��v��`�������Q�1w�P����0A�(��ʌ���)��z�2�39FSh}�����y����Ή�m3����<��e��5����~U�T�������C�:��y�!�CU�J�E���[��-�I��O 4xM��"�~��Y�=aF!�<ڋO9��Z���C���.Y�]�B�'u���{���*۰%���#-���c��K��.U&.+}�nM-��)
�{`��9O~���Hq��
	��^5��N�y˔��T��ml�mjī��%7���#�l �υ��h�1��E���\H=�ߩ\�=
�T�Avp��8|4)�����G-xK��͒Q�4���1�C����*f5����
�V}�$����Ք*�%�LwUoz\#Tp��7=b�<�_���4�v�Q)�Aa_,��E�{�㣷��]Hv����T��r}�3�0�F�ɷ���	�`�sP��2.iw]�%�n���b�̎%�U��>�K���2IYߊ)��9l��<�z���� �,Uc���08�v�4\�`���y�s1���*��@��N3��8�D:����'l��s��j���I�5�*LK��E��k���l�o�=��&�Ǻ�U�sT��d`�'��y��+������Eȍ�����k��A9�U���}�9�����N�n�'���!�7K�_�r�VZRo�=c����q4i�k]=�,�0�T=�R����!����o�IF�G�#\*��eN��V$Sm�p\����m�a5,m��>POw{8�d�6R�����  �	�[�Xn��nc9LQB<�]�F��#�����Wd�0k�Ea����F�����薲;G��D�h���t�ri���y�E"�f�|�Z�)�����Q�Vrz#،Wٷ�knD�K�rQ�!���h/D&�`����`�w���y�[�`�5�鉓}x���(9a�ZV�Ri