��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�Oo�Ne�<��!G�u�uO]�nG����W��1L���a�KzܸƠC[#f�0�����-V_� 8T^(�|��Z0��+����[VT`�c��A�p�����	�S��60�W���)/��L��A�g87V�c�5�_Җ��sd�����PA��C%#!^��M[��[C�r��O�k�#H�w�c���T��7rC��i ��)�sI?�V�K7ۉ0���F4rg���W��:����J����Em��]������ \do<<(���1�'��*��{�"�%4P�D��V"R��G�xVxV����\��T:r/����q�B3�z��2z��un/D��QG%�=oTK�;�I%�ǿ���α��|��mی���o������?��H��t�x��M���ug"A��w� ��fS��������`���?��X���N�����^T(�u��p������l�YA?����L��bI���7lc�f�6FnEq��Fl��� ��g�Y�)RyX蚞�u����^�vTC��n���S���]���TWq�x�B��˽{��`��*����h*CN@�-�C>�_i���8_DyS�b�ʥ�^vo�0w�����a�?�1n� ��Ǭ� AR�ϓ\6��bu�_"[�P8p���	��1� �өVt� .m3�p���Qr�%���Z�^��'VHDb
v4�;/��u�_��e�T�ÙRj��]���u]/GR�r�ۣ|w{拈�?��x�N-�,����=����B�H
�b^"�׉��i���+$}\T~YַD�K�1B��q����u�(Rc{3=����ng�8Z���5� ṘB��h��T<�;92��W���}������F�b�I�:y><��#�c���Vn4�{Ʀ1��Qx�b*�G	� ��5_�����քl��l4���e�Iݞ>�#6A���ؼ=�gi��6	���D�8�/Y�ėגZu'���^��YD 0�^��q�<�l�Ϻ��+z���L#�ʦ�LA���d���t�.�PT4"�̣�H!J�5G���zR��h�x���2�E:�X������Ѻth7�]\r��cqc�\����.o��g�󼅔b�-��m}*KU�s}B� �~S�M�q��z`G��u����X�����1{��Z�7Z��1 �^>-}�cg�u�����ЍC�7���~&Z��c������^E����.l�+�0���qڞ�F��6�<��<o�J���>7�)���/Χ��vWew�U�U�p��������Z��Q%+��F�� cSd{ t�Ғ��A�"�g�kզ��ᆉx�r�vQ�Y%�K2Z�S��*�UEc��$
[�硝5h�Yi�Lښ��R��D�O�.�xWμ�ջ~� ��q�9�L�<�=�C^6�Y'ט�ў'�W��zV&�US(�9{��2�ly$c�v[����c�n����>��CG}�J���>����*�K�>��L�RG]*�@�ѯP�yi�a8fVݠ�Lb�ѥ-ע{e}�v!J�
]�]ĈYB���L��3���<�+��n2�
$+���PYu
�f�ְ�p9U_�8B��Fr[��2�>��+3�7�bP��z�M_�?�'|�G�d��@E6��>���z�>?�%1��{,:)3�����m����C����~���x�I���������)�7;��/_�����^WUg�t,�)C*�Q�0f�:��v��Ɓ��sh�o�k,;̐F(vW�[rx�9e�ez�q�r<2�a<�1GŠ�C0��(I��Q��wUr����s?>�����ϰ�?�޲�dv�/�R �>�o�D�Mӝ2��� 1��ILq̲��F-�X�c�z�%����D���KӅʟ��mS�����-'sPZ��j���d�ȵn��\K��7B��B>R���)���9�z
��O�S��t�,Q����=d\��� ���Η��d�����QJ��9�@�콫�'{�z�!G'��p��F�%0�rc3��jV�O���x�a���u(��h�;*�(.8S�
p�n�U2��$�#9�p$�f��w�2ǥj�����/�s�4;;�u�i�%�z�1ijEAN�譛@7W��n�E�lD`�J�K=�uP�0n�U)��G�PM,��v����So-ZO�����|�r�R��k5I��xr��rxb��C�>=��J�u�y�<��&�6�ʑ�O42�f�}t���ӻ{E�ᣬѿx39#�;�m ��o�ļ��oڨ=���xc��� X�f)Q�en:�=T)�J�L�"���Ԟv���u�0�8�j0�쩀rG��䟎9����L,s�h�G�Ǜ�6�'P���m@!H��ud������\���'|:�N��)�K��\�7�����b�`�"u��SBi��6l� �*�r=۱�Sw��]1�,Rh#��D�o�\�'
*���AɌ��ל�{u
!Yz��ۘV3�IGC�m�)sdHC{a�!'l�̣�:f;J���	�2T ��#��DeS�����d������e��r>5샻s�\���`*�k����dS�q��鄔� ��)��[7/%��ި7+A�e�oe"*;c�l�YS�>!?�ef<�jѬL�09i��X�G�<<�~�kU� ��iϏ����h�.��hQ�ҍ��!������I��n��wby��Y1��(j?o᪅���ͫxx�^ղ��y�5��Pm0L�&=-�3w0g.Zg���ѝ���������@p�B?;������L7��lFM��r����$��Ա�^����v�,�k��I�"��gߒFi���<�B{!�FRQt?񬑣0��U��S��&���dJ��d��|$&�,��K�>��5V+�[�A�G���<�[���Jְ8Yd�I^uB��V5|�G����矕��E|�|�m��7�RK|�����S�Z�51��@��R^rT�w�dS������'I��ݿ���K�S6{��v��������땧'	C�6	�q{x<&���Q<R��	bJ+\� jc�d��$V;»2��N$Ý�҅$T�g��B�r��4�͚`u�G�w�^a�t��H����o�UdYY��~�I��w���;\��e�|�gW�����ô\��R	3kA���s�~�guZF@����)��{��؊Cֻ��L$6W���4Q����|��x#�+ς>���F���Ͽ$! �TBX�|s�Zڈ��%=:
�+��E���z?����I��%�u8�{�C�ӿ_YC��/�+�}��B�/G=�RaW�d��f�N�i'�D,T>g�GO6D�|���Wd�>CoJ~F�6��V��Fei��o��+��CN��~��*�4�~!�^��1��p�?��F/�f��2�`�mx�k��P�:�-�@η�]"��we���#�Ko��lq�i�Y"|�Vdjf�5ϋac�d�õn��<�&�֨�I?�_�~��O�?ҦGHM=ڭ�`V1�y�SL�Ŋ*"@�����3�m�|Iӹ65C�m2!�i�����^H�;(k%̶,�&3��4CV
i����ZY���S+��]9�m�����0Z+R��S5�9� �T�4�9�(1변�Qd#I{s�&Ҳ�KpKk o��H.��yF! I��lx�y����@����/?!r2��D����Kr6$�3���a���j�{BE\�)� ��T���L��E�uB�1���p�Z��л��/K
+�.�X�e�-���셚1�:x��a���l���>�Z$�ɔ��e��3z�ᨛ:��c -�h@N�ʰy�zT�ľ-�hA.�6z!���;Z�U3�tG#ADL�~��Um����J���G���kC����]��t/���߮ K�'��W&K5�6l����n9}-s��/Q���>��ꛑ�l��CF
͵T�*���i7�3��%M�������Q�k�Z��%��G`:15T7;B���d�\w��[_k��a�=����L�
+T�'�p�Kn *�b�\����-�-;�U��r���!� �	��4&�}���Y��DՈ���y]��1n X����L��#��'+a����ɨ�B�pCl��!�4(2`�"��m�S�w�M��{=�N%)���IS��;Dlk��Ԭ�Kw*U%��JB�Pk��QT�p�U�Kf�`o9�f�i�3�-�:�S�@�id���;W�����j�8ɭ#N�W��C�;���0%����ᘍ>U:aa�a��/�a`{��n��5q[�^Xr������i<��;��4ajD"d��}U ߳��ܰ-b��.���7]㑠x����Gj9	����;$����@W�mW��Pm�D��x�J̔�c��,4�-�����u}����pH�"Jk����e������V
����8�m���'HԂ��l�+��GK�+�̼� 3�����2w��<��oJ�&6墤��Jp}	�������Y�cu
p��w^y�9G-w"t���V*�u�Dl]��e>��;�=EN@�iM$[�d͑gRy�� L�N����fW�4(�����[ �Z�bl_����zk�*LpX ��;�o�3��*�T}���>��_���&`����0�
��Β�0��Ư�Y4��kaCۦ�Ǟ(�%9I_�v-BS>�t��bD'�����"��f�m��Mj���=���������m�%+��k��m��65�i��J^6��;�k{�x�Mi�*��iH�)�$Rԛa�co7J?
����&P+��B�U��֯nu���UUD?p��bc�_�e����C�n�ʨj��B)��82������Er�$�\���~����"-�i k���~.�� ە¨�d\V�il3�m^�Wwe&��/3�k-�)�R�e?Re���}N��4�њXA�O�u����G����	>R���J�9��M}	�I�?���< \�/�C�Ȼ^�����0�V�.��#��8�B֏�vȐ�h^���C�,��J�^�0�trd�/���k��nůU���ₑN�*��c�����>�.�gYg;B�8]��NX�Kޮ�D�D���G-��s�tϏ��4��R���4'�z��ݕ��!���P�9�)sKM=�Nқ��^�Bq�H+�+�	�6Od>&�����Cw��Fɴd�;-���z��H�B2��L�L����WZ�o��w{$������K;2�y4%�/3�5r`j#�1�E O����	�U<����o��.��ڊC�fB�$c�y}7��}z�6'h���o�x����J�GU �[s;�ɣ6��\5S�����+��v/�`���Ccw��\����L�E�C���IfPr1]0S���[}��6�|g�a=4G5d�u��+n@��-�)Ƿ2u�R���d��X�Ķ�|�Q>�_����&bm]a�)L)�l������S&���r��2d��z��m�k�|}�C��xQG� ������L�A 7�����;�Φ�����^�����������t����En������<bi����7X'����;|����D��3v��P�j�Rjo���_JI��Hu�\�+��~i���%A\��i�=��(�������K�&��&��@��aH����� ��8E��!�Y(�r^IY�_x�H�,�թz�ޘ��57�~��������ef��%d�;�͖��DEw��h����!/'W�W�.� Oݾ��S��Y�Oi;�.A�sSp*?������U��'}�F5�]b�^X\��e*y�aEw��Q�Y1����g�e�^P"M^ΙH�-���gp���B��W��&�\�sVQ$/��2-�'�ͅ�X��ߧ�CT��H�!o��R�2/0�7�4	W�����a�o�� �w�Dck��z.B���j��,�e��P��o�CKJ�A��~���W�o���͏ϳfr���%8�3��F4y ������L��(�֣H#ڼ�d���{W@�I�� ��z���j9z����5쑻�A ��c�>cb�b*�yy^H���#�0/q��Al|�d���pj�F�+�0��I�?KЖ30g��}���X~���Y\/��M��n]�]�������
L��q�e�l6��n.� <�e	�,0�ü7�D��R���3vg��e���}��Q��J�*T���Č�h�6��D��"�.Fi���\����5���PW��2�>Q�SN 0,QSCdl���ҳ
��W���Luҿ̿�x$)�9����(C�E��=2�(�y�O�ES.s����un=4�U��-31h����H��27 z���'Dm�`x����P��B��$�����
}����{�(�!�����m�p� ����L ����>U�fe,�U;ҿ��Ӭy��9��͆qމ�o7O� ��R��}6"��y_O`���Ȼ�K��>��S�G�iH��N�w���Zy�9������a43/+�lk�K�63�c������ID�H,?�+���S���(���0X�?�M����zXd@G������X4]�.(+x�	�5`���z�Q��&��T*7W��^6��}��)�7R����ĠEX�U_a�i�m��z�M^�UG�6M�N-V@�c��k0���i���ׂK�O�%�
�lQ��;H�0�{�[��(��;���D�d�U�n���7*f��S�TLP�ݾ��F�a��+�ҟ��E�]J7<Ĳֶwɒ����(w�����7�Ø�Q�[���:�oI�P� H-������Ⱥ�Xm�|��8c�=��HAo|��t=4�D̾Nl�W�7��v�s�o[�d�C�m�@V�a���L]�I��=�ǼaK�i�x���>�Ǫy��<K�c1h���3r.�Gïl�%�$������`k���gl�� �8(����Fq�S0=�r:�c��
�z�Y��I�⃴��Q�#���.sy"��/�@�cv������O�Ȝ�b�w�s�x�. ���}�ȫ�3��	en�)A�1FZ^����Am���r\�ݘ<�p��V_h��.[ћ���}�?Y͛
x' �OvP�!��.�+YɡUA��Z��,�ٙe�gj*��V�?��\�����+��֍�b��\�����{u��8Lww�,�V��-��A�c�w�֌<�ڷ��O�*�ޑ����������Jy���ů�u��$��bFTX4�s� �s4P)i��ZƎ[�%ky�+�, F�;#