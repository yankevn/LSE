��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~R#b�Mҧ��p���;��aC�w�!�,l<�(:%܌�.x�ro�K[J*���Y�h�c����n�w���S�9�2�w�5�m��7_��^�3"��<�C㖝Y������H�Z�B�ַ{H����=�b\�)��fG\^G[����Ҕ����u�/����č����Q���?ݩ��_Î��km7A��P�G�u��A�褒H^.���Gz"�:���!�k����jt�j�ά ��֓B�\���N�6(� �y�\2������6��0���RMA
���4����b�'%LMX���(1��`%r�=�x�mg�8�O��B���q��`����[�%�`:�P?ڐ��%�,��ª�����h�o�����jN2�9ZY�He�?���׬SRu���WCL+��o#tz�W%�t����7$r6�e��ؚ�?xW�)<��~��H��'x!�� I�>܎��Ո*���v�Ek�b��w��^z����~CK/�2,_�¿_��n�@���������a��-4JY�}_I̯�Oo��
@u~��tb���]�x��|*pg���bm3Sw�W-�"�8��1���6P���^5� �����F+�˸>��(�3�6C�S�/g��!E=o�,�������{��ݗx���!C����*���ˏ����e�>[�f7��P!��'|�,x��'B�?�1�'VN�$f�U����9�r!(���G��-@��C�3-��YE���@TBD�d���v}i�N���X�3-�w��s5�<�>6"g������~�����?AP?�'��2�ED�,!;�	�|���vk����o���E����,���\\�b��b��̘���}��E;0ʬ�nʊ�w�KƵ�����I!{�'4��I�ۮajձ:1,�������Z�|M�S,��@�S��4��y"b3�;��>�o��Z��:z�!�>�i|����Q%9���vg�m�X�5���B���詢۽��)��D�����>G
���>����mgkb��%�A����X*ܦ��d������7����<>������X�=�+c:%q�0�l �G��@�XI7��ݰn�X�xp?���������a���.�5猶�.?��@����i�46�����A�V}V��^����Z倜L��(;��ޘ�$[�L#$�/9!7d�!\�w~ƚ����/�{L��5qE������8d���#������oKZ(�w�;���
�,����`�0�4�n:^���#�o�����ݓ���Fm���2ʹ�Լ�M�kj�c�aV���0�m*��Y�G%d�&������l�&N넟n��j�������I�T ��R�VQ�=`���Sr6�[�:����d�@cr�Օv�=�Αw���,���'����-.���p2�\�7��i�c�|�F���V_H�9	t�q�s���f@��)��a"��N�����{*���i��N�����8�Ń���N�_���0s���?�u9��!�.��}��C�{f1�c"j�uC<q
�(�`�X�l���ě˂2�H�j��j�~����I5ʅ���*�րf�SV�D��_T=���� v����g�S��w����x٬XA���QN7��3�����UH�7.@�s�:�/؇T�C�qO��&FK^p���k��0���&����Tӷ��*�j�����&�<!~9�x/v7�k�fg�1�z�Hn�|�d��m.���DHxU�:���)C[L����p�
���ҧy����y�E�﹁�rƽ��u�����.��i�l��~��� �q�ep5��.�T��_�cI��+mm�L�1��6�gf]-�����<'�0�4���A�e��5����<�	f1�eV��J6�h�@��?k�o��pLGe���4��Eճ�*/x�4pek
���oB��a��*�܋`vCLw��g�IʶD�O�������no)q2�x�b^����yk�U�Ϲ��B�BGi�����m�I� �~��}�C�LP��T�*J�"��������e~��݂s�V�iZ��?&�.[qs�ƮN��f�;\t|��Oe�\l���d�@��t;����6�BM�P��^��.~���KuGTނ��M1U�����ȵ��/��УV'�+�qA�J���]'g:X�ᛂE73T�3Qj�
9�����ozy�͍���	�����B,�9�ZI��k��ը2$�_���/�s��Wh"u95}c��T���[��8��Y_�|�w�:!2��x�#��|�^�iZ�l3���Sj�Y��@G&�YNHq�3��ݛ�po�(%\1<�\B\Y>�:>&`e�*��#�leآ�$ؗڔv--8b��xxn-\Г��wy��V�(��������$���q趕��-Цm�kb �w_�{���מqΜ(���rbCf}P���qf�O�r�Ձ#��Vli3:�y��%jG�4�Ą���\�uӞ�.��Aa={A���Rt�A릖���0u �1i�_�v�9�tX�t���}���t-�evOBO�U1�&��$�џ Y:��r�o�j.B���`�.uw��Lɾ�su��ݺp�*��Yķ��<b�gޑ�1k�!$n�7�+*+���^�T����,׵�,)�+f���T'Sb"��u�K���-O�0xI¤�.�y�V��O��1�ʎS���Wׁ a\�[�]�fmH����?�����H�$O"����9.�!D�\�7Y�<�j�e6�6V��)�t�+*�R�;�K>�]r$�Y�l��8�!�։��+憲�����y>p�Lc%��Р	�����X�����NL�Zk��n�Tw�V?�c����B��	vJ���#w���Y��E%{r�[d쓑�P���o˺|�	w�v�x;Ce�����C�*�]8�B:~��z��צ0߾A�eX�6臖�J��u�!��4L��Urjh@�)���p,(Ϟ��1��.�&}��Lx��c�-8�Qz�#�4�� �ZD�I�M��a�65�6{��-lS���\��K����rP5)Us��:3�$�����f��w�\* �j{tx]�ꐭ�윻���w�/9�%�)����+�P�GY�W�����ad�Lh�U�����F�DM�$K�������3(�ߗQ�Q135`��V<_���C�Z�[��0�����t��r�S��2�nUZ���׿��c�L��Є�rF� �S���<� ���~�_�@	�4\�9����Ys�3��_c@^�d�ZC�k&	+8���&������N|�~� �~񨜹@+ƇYBJ����RfQ@*ۯiF��M2e�x�`^A��&3�PW~p���j21	�SR�j���:��H��m��xJ�h�<Q�q�#a6Um�e6VzZE���ѷFc��&����^��Ɗ�+_1Q.B*��x$�����|g����!�q:��[��@�..�`��N�`����\o�Y�#Lfz���Wu�D���Y���ˮ0�r;Mw�`͎|�L�M-zJ�8dL��3&c�l]1�[Xs���C$R�\��9(E�"����D���v^�R��9E� ��(.r���e��@WR�K�E!E(/R8@*_���*w�\L��۠�q%��+w�b~�}���j��ښaz�����'6���3�N[���z`����qU.T��'od}�5��`˶�ˉX�� �Y�5�����|�	N�+�|�x��jj�g̲�_��T��\���)MR<-ۧM���_Mv0�kN������4ܶu� Di�F�J��^��D�ѵ�<{n��Jnz�����q���T^(��-mz�@�$��x�x��k�8�}�k�Y������m`�8^MJ�-�t�_�	~��uU��.��~�kNo���#��3�o ���gJ%eEʆW2`���,��Q��1��Y�y?�nD�3�"���4S4� �7�R�1o��,� �VkQ���d�r�d��dIh�6V��_��em�M����t-HhX��c�E����V�P<��u�J�^�F,h6B������g	�-0 �&@:���Y�v(е�c��I~�J5]#vS�l5���[C����S�?j/k@���Ax������!�`�+C�b�nǂ���\���HiX�
���%= ��>w�a��4�>���7�ڜ8h����?��C�5��P���|��r�&��q��*s���t�i�v*o.�6y���s_?Po�r;p4&� �� }i����������h`:k�,�IK}�*�fd��G����D6���Q���m�'�����V��M��ī���C�J'��|_f"d]z{�"�m�Y��[����N����@�����p05*ۆ���`C[��x��0��!������Dvr��ɿ�B5�Y�.l�-�
J	m|����A;�+J�%N���[��\��<���f��o���B|��Jdv��U'.����-}8Y=SJN�Uj�;�.|�
�[�Jf���OF%�/��\پ'�����^����c��	ޒ�o���g�JRu�Kub�	��l
�y�iᑐ�4��
�S �A����	��Jo�N)��Y����G�1]��ϳ
�@�m���hd���(�Vt�DG�o��W�`���"B]�D�n�	ܡ���0i
I3Y�x���Td^rk4K������ޭ+��z�D�j���X?�DiXQ��7W���S�R�Z!@��;]\��"�;��/g�6��} u�F*�� ���z�j$���n���鶆�9X���$ŃL����3�P�p���i�\Ua:|��ΤP �,F��Y<�ʍ�E	YpĝB���ū�����k��x+5�חt��B��QCؖg�����68vo+F�enf.T<��`�M^oz���o=����cߔ�&*!Ϛ�s�L��-D�l�a�g��;N�*��&�p�C��<j���]��e c�q��;����PKϬׄ����7L&�G�ĩ �b	��T�A��C�R^�G�WO�5C����?k*����f�bx�t>�X^��5��	�X�����>���;?���y�U�J�p�xo�Kh:�i
�SK��$��Xt���]R�'�E�S�%Y��h?E�rD{6L�5�����'���^IW�\�W�֯*�#��Z�w���у���Z:��-B΁? -��#4@��; ���D��:��c�7����q���+�d�3ʀ7����p�M��o-�TՄ'Ӱzi����
���H���ۂ���Q�g�<���ޢI!��3�[1�����M� ���dށ�x0����sAl�S�B<�ԕc@�!�^w=�����w�f=�Ҷ%�n��V&&�=����5 �Sq�*G?����zbT���(L3v����C6�����&��%�F>X�}A��:�0ޓP����fp�0��ˎ��w' �2SF%q��7�v�,�H��/��M��m�T���:�����G������*�q#��s!.�z�dP�Q�
�e��+uM��%9�c�/;�_��O@PB�&�Q���kѾr�@ܕD���OW�=�<�|&Q��ϯk,8΄�+^:p�m�C���Zg�l��}7�����j��@Kn|7�k�)��v����)��lw[��J[ƶ'��"�w\��c��������"�m̈9NC�g���4��?w�I�?!���yl[� ��u.�`�RA���Zu#�!�$����IZ�}��F�>�n���Ll��9�f���OR#	`NV�_��Iw��|ח�d��h��'U����r6����!�+�7��JS��Xukű��0���s�w���̔��`]1�<9[9[\�R��-ZL��Lmd���O�n��'��DE-A���,��w6���?����e�o���QK"�'��V��'��<�ie�0TZt��}�K����?$J^��,�b\,%��lL�@�9���P^F��B�����a�̱�Ί@#�J��ւ�N��-���Y���o��X+_#V>�0�Ԭ��}�>=�6�+!Rَ8���r��/1���A��y�pǘz�d�ww�[Vư`P�<��t��!ƫn�CA�����GF��{8��c��&;p
�ĕ������e#E�.��g��akKK&�n�B�8�1�
\�<dr'�V>����M1����I�������v�����w�z�j� �������W�_��O�R��}�Cg\���g��2��K�W~�rvO�J�P?X��N�8�w��������� ��α����\u��r@=cs��H�SPR��SX#}ʚD�����$���P�D{��������߃Ǥt�1ͣx͌��.�hC-zCm��c���b۾�^ ��������R�޿�'#8����iqxq��}����]���$n�������]���	5:��yK�-[<q���	&�����҃�`��D�3N���1k��5�*Hc��)`J�ko��W��T���]��
0��Mu�HqM"� 5W[���x^b��,WzT#c�l��4�Ef���G!6}��_���}�k��ƾ,mדּ� 
�����QZ�֞f׬w�_$3=�7V:%���k}�Z��#���F���O�������_�I�̛#8EW/�o7]�zis�r�sc=���Wm-q�}�0� �Ym��q��r{,5}�DuX����Ue�$(�y���6���[ �j�)L��F�����3buzR��Q-Y6�µ?�`��)J�۶�M��E��s��<�b�8�πwZ����E5.�9/U�َۉ>�%�=��E�| �`��\�H�6
�"ƅ9�1_߳�/�J^e�� ���Z��/��
Dy��TI�g1��R�,�ӷ/����>Ϟf�Ҕ>8'������\SG�_~%�WVg,��Y;Q�ח�{ן76���L�4ڗWC [�=ԸBO��:8���(�B;By�_�0���5����0#�ɪ�^�+�~�c�OE:���4��&�H�� ☚9$�g̐Q���g`�T)��v�axj��ݨj	f�[�Y�ë��i[ +������O�����~��6�D3�<F�5�ę��e2��e��u���x%�Qp��l�R����5�"��YV�͚��*8-�_�U�X�>u�e��u����8�O�V�s\u^���6Ue�Y|L^� 
�ر�,a���V3C�;�j�L�M�I���4����Nhͦ����"��W����E���S��Z^Hd�A�6f�z�O���(�h���/o��Ź&u����_�(Ja6Q�	��^����X�1}�r��ɽޅ�����ǚ�����]�̒/��Ob'w��������h�l�܀嵶�}Ls;�ӆh�X�b�A\�@E��"�
�6�~a��G�3-p�RJ����������X��fՙ /�D�wU:��OBTb��F澪�4VE��l����7C[
�/(V�d�*bZFX��=DN��:����#�o/������Ղ]>���0��+�$��k�
-87X��x��*������Q(.e@��އ�i:o"�u�vTЬ���恴)�x�����>�g��i���s����)����P�����Uvt���<gBa��J����WDwោlN� ��P����)r��U�J��?@#a�&��)'}9[�����[`�fӫ�����/²z���;�����9zǳx$K̃[Q9�)��J�\���mFr�,�*h��x��6s�\p��v���8��Ya��d�"��_&�k7�������N��w��;���nT����TϮ֥��1!`Lc#XJ�A!CP3`�37#h����_Xw욨
��� C�A6#�;��LC�r�[�6+���:uI��-�[�g�mXR�Wo�ekTD���	�x�J���*����L�Ȩ�ݽ���*����}:�3��E�V>�a�~|T��e3�8"0k���l��n�#'�t�.46<�cY�+�}Jo�MIU�WP����� ܂t8�j�o���;���Z��d�ϻ]X����5����HX�W��$�WNC����|N%%Vz�N���7y+�&���gꚧ�7B/X�e���bf�x3�³@��.�;�e2��cZ��G�E5��D�C�tk�l~�V]}3�U
D~$WB�y"�$NC�ɖi@���M��UH�{� <l8�Y3F��}yKA��RO�kB=)$*�L`��?L"v��ĥ�@�"<t2��&S��.7�DW*zGt���{�����G�n�K��$|�s�'wc~�c3B���ު&�5F��>8�g��v�5Z��(��3"�_��o��·��:)MRŉk����Lp)�/ ��F�T����b	Dfӆ����`���#BI�ݯ�.)��b>�0�+O+)�w���<���D�Jm���]��9����Ť�O�F�4}6v?֡�d�N���C.o��8ÄM;����������?�|�Me��~{�����ƏߓC� ���+?M����Yu�2�L�p�$�Pv<���(j�?��Z���wy%= X�K�k���th���S՞�@*�z���u���~1�3�3�R�c��|M�`(kN�1b� �Ȋ�7S|�B���_8s&��)μr�@惧dl��4Jb|�gR�d�<�K���q\��w��/k%$+����$����y��np#���~nA	�Cl8�	r��^P0�U��#��#��Ip�X����Z�Q~��Q�a싹�l\8�s�X�Ug�y��Z���"��K"����^W`���]DL6k��C-�yg��y.V�νJ#dB|0�:��k�<gMCʴMJs1��dK�S������1�o:w@h9�y��	k��A_!�pŽ��fZ�dfHO:������bS�N��1	@�ո����V<�l;���/��JM���*܎S��"�z�Z����X^�ft����u�-$�XF#���z$�-�k���L�GM٦�uh2}WK5U���l�<�-�μ>�r[���E't�T�ݸ;k�G2��) 3�b�B�{o�=C'}���:_�+*��g����S�����+v`��~���@�d"'t��I�]6�u���@��F��`;�K\�
��Fk'���ĥ�&�,U��%s��:_#p�p��bay�Y���DÐ���^����D7�Հ��ܧT$`�����;�[�Am0*�/x��j
ç-Mu^u��}:��X��E�!��RNZO7��ݷv�g.�ĉ��FtUf:t���ŏ��ϟ���٥�2�aτP̡K�yFW�^`��a#v,�������;}��������������F��׊�X,�_��	\�hrXY��#�Qw���L�׹����ZD��������1D�R�2��d;x3PE�@b�S4�}���j:>��N�mO�a���ڜY#�\۲�e=o����o7jdBm�sF_�ʥ�4�������B{s[Vk�W<�O�NV���+ģ�Ғx���LSg\�TB�Ɲ���4�o'iv����@H,�5P~��1)%����Bv6����KH\'߬YC���(�)	y�2�%Q�%���o�4���n����p��h��̂�9�8R���J,���8\wB��жꚴ�5� ��6h���l9��N.Bn��`E?[� �J��s)[�_�����]U��C˪.a�
�B�4����B�[1	�"d�[���JEǝ��G��U2��f�:�-��}B����%
8YT��9钘���ܯ���~�l0�jp�P���g2����&��F��a�G���B���"��N�0PE%G`��?ҥ2��xEnjP9�k@����C���H�{PxNW+�[7臄��p�
�^�JF��d��4�S���j*Fs rx�0*�v�\�\�8B�-����x*��a�<��j]�m~����o��Za�5~ۡ��y�J�N��MM>N-�>W E	���5@T�ɒ�E[-#��en�d�@���+&���C��.8�t�щ�R80�ഁ��Ϟ@�h��I���}^�1��[1,� k"�$������t�����D	�'��ڼ�v�������B����(�H{s�4��O�
����NЉP�r�LR&�@D�r�Ǜ�'M����Y��֢-b���Z����Zz�`{�֋֕��]�ɯ��+���.̅�҅<����#�T2� G�v>ɡ�� �����H�����Q���b�{�͖�i+Ѻ��~%p��F����g!�^���P��EI�)��-b(�W���Zwg���|�I%Q���j��'d^��6�"�
��u�(So����Ƃ6��.�5�(�H�W�:�}��J����fk<{�dʹ�h�%������g%W��J~K����o���(:�'����޵�����̉���1���G�1�`�3�98������$�y�����oA�����@ɗJA ����tB��8�M�e�Þ�`�����A��}��sk���4���1�>����s�;_��ls=X��T���^h�r1t�+�b�A,d��jڼ��M�Q�*Mg���1	�"I�ز�Ho����2��� '��t�������h1-ɣm��9��cV)1��Y6.'���Z�(ڑB���B���21���[�������6��:Q�yv�Ll ۙǅ�m��G�L`A,ґ��TD��Z%ӡl���uyƭf뗂2"$G�'��4eLE�����,J�w�FFxo|e�7<�"�r�_�o�.��Xtqi�����+�ʃ߲eB��\1�,e�VS�(I����r�� ���&�5�s�#���d�8�+���L��sm��#RxfF�5,h!�ux
�{���dP��A��_k���Ebe$9���?�X;���|�5�$�8�!��w�v�9�P.(�0nwp��z����QQ���-����}Mܘt�v�3��(�����6
G�}�2�ΫG8ќr����,!�Yf=E
�
cjT����y�YN6(��wk��ngR�N��1ޡ$UA���F�A;dY�M���&ޑ�i�5���7��8@L�)�gF�m��x[Z��Be�Һ�V�s��E��^>$#��{� ы�j�7:�̫<GvQ4�2N�q����>Al��9K*��� p	�%�}A�2ʖ�%F�r�!�:]0�蘏����t�>޼����u5����-�����LrY��;��t�+����i��xh"u3�+I��\%�v�k��f\�a{�A�lH_�$m(frڑ�t���K�%d�/�;L�{��:d�/0R��^a�J��dK�X�#}��{}�t���������}p���Awk@��BZP�ZS�n�	Z"��a��f�i������p�~�K-��41��%��d�73ҙ�P�
;�@.�S�a�o�I j\�L�ʡ��/@=�kȁ���֥�(8�-2X��-�2a?I�WF�YM��z���W���E�+�%����NR��ZI@'`s�=�>����Q4�@T	[���b����j��X�M4By�^}�W)�B��.r��e5�]��R�Q'�"���Ǧ���og��2DDj�ha�X�d�Ur%el"U�	V�Y-�d��¸�}p�,֋�7�'�6P1�l��N
������'E�3��o;ӿaW(�H�� �A��FlD���o�K�K��/���k��t�n�8z��u}��&���KC�0'�6�,�|����辛Z��'~�0�4�(_�I���-�u�FV��:�w�qva!��&���������V�<�$>��甃�>T�p7�����_����C��j8�(�1��t67��pt$���z�] /�G�C峎�Å���z�E����B�11g�� ��^TX%���jf�~Wp�.�v׉��_��݇k_��9�3w���LkW�#S�s�m�X��m�q_�K�PhX<2���*s�P�������[Gw��BX��kUe��~���>�;���K��Q����=h��8	;Wv+U�<����_fۋۊHLNN���q��s�Ŷ�Tn�7� �=H"��ޣF�l�xr*Z��ۧ����;`=e�ŇԥZJ`nSNM,�e�%	�^PŉI�#C�f�h��4H��J�JI�2�·���D���(��m�"�#9�v�y�m4q�����.����6�Ά�\�y��ܜ�ʹ�K���&������=Jq!�du�B(�ɒ��Α��ڱ����������̱�������~�&O��b��T8ͱs3x-���3ϸ7���T��ē�n�:�E���F�s��iq4�F�n����ޣ��V#�׏1k���&|G�*���MSԵ$��	9��;u��Z1�o����pm�{0W9��Amw�Q8�c�)��@6?[�]�{av���ĪarTX�f�� u>�"'����� K�\Q���F�U�e,n���uS�n8�X�9�o�~7�
6d*^�?c�Sv��at�ۆ��bp���Q#$�.hE@gD�l̮S����y��_��x����E��>��3�c�-î1��M��^��$��G[��p�/�6��.e5F��Iq�q�Ow;�����o'.�)�N��������StE�����@�7.i͵�eA��eTtZ���*Ԙ��>������e(�vN��l�?R�A���H�hG�U�j���� :|n����+z��ڛ|Hex����.2׶�`����Ȭ�~��Z��`��}
lgk2��}^]ϢOe;��J)�MZ�SV���O?]���f�Ýɍ�K����ͮz�.�}�8��%��'�X<ޏ�|�(Vd�r������6f4�`�a�o�"zE�s���*
�C;AhVv�K�����f@l�Z�jG-2����^N���>��A�譢C��V�3rZ�	i���f�DW@|O�:@HRz�k��Us�<)�V;�����{1,�����#�"E_��f}^��~B��3� %ZÚ� ��m�M�{�ˍ�G�TF�f�]2���B��w�t�c-��n�h�H')�ޏy�Ŧܩ�v�f����{�`,VA�(�W��Hg#n*�c�]��U�G���.H�=m�Lێ�*猿r ,��m�K;����o��iA��2�;;a����E��JIЕ�g��<�N���m���Hn����߽������P��E�^	q![d�+}�+3�
@�`����^�&��M��=�=DqZ����Cmc��D�Ĝ����C���H����®�A$��V��{�c%\]�/g��;�Jg�h:�Q�(�扡�����]g��c��N��/�tK����?M7��<YUAF*��bBw��B/�}���$תv�y��\~����?&V��;>���X�f��lo�[���� Xl3s;רM��T��6�hmbY�z7��2�l�O��QZ9����&|�Uѧ����wX'�4^�fW=�z߲���Y �W�����#/�����J�����A�y QP�|�מ'E�c���R
�r���*͌-���̢'e	.�+UjOݯ���4>	���,�dWz�;5�G�Lb�P�C�hi���D�\M��Ƅ����?T�s�(���j+6	�K�P�*�-�KZ�q�F�Ҩ����l���ݨ�ޗ�D,rl+��Rq�ք��~��B1CAuX5��
Ö�a�A�[��5Y�;��Ɓ�����&��1�gm�:�#?���8Q�O��;p6�6��Z'W���غ?R�2��vHB�WւЧ��M�M\˿�br�ך;�e��F݃���iɞ�KF;3~�����8 P���Џ������k�Kj�#�ZuX%�DĞw�ҙx����5(U](Ӏց�ygq�)�Nr@�T��$\�Q��V�D&�u#0��MΏ:�SH�+��%b�rÃ]h�?��1CT�!���l�K����ڮ�K|�e=�\�͹KPhes�|�m`*�r��W�q4��!����r^��7Ҡ�L�[���(K�WKc�-�<<�ܒ��a�yb[M������I+���L|�+g�O�F;j�Sl���R���񢢚�8/ i$�lE����,�q�yҭ�&�y̭��ll���ƈ(/��dL�*H�ղ�6��B�c��լTu��H�-�Kw�<ڶ�p(����WS���;%�)�ᒷ�ž�z�ő���s���4u����v����n��X���H�X��u�'G;�\�I�^�,��p��q��m]m��#��Iz�a7yf�K����Z6�����G�(x;��J�E�����j�V���r� �y��-6�w�$�v5(��1�	8�cH)!��oag"c��gݝ�C���.
�aM�TzM����o��:�>����Y�����YY������e�9̍?x�����z��V��	���Q��N�QFsR�ܕ�X��ځ���9)"0�r��Y֯S��Z���'�V�����t��>c�'�t��/�ZȺ��ŮG���F�UV�]6�8� ����ܥ
�ӒS&��lS���'���Ս�%�t=yweƮ$R�;~��X�};�j���!�����G���B���y����^牗�����$3�|Q^f��!~��Z��Q�y�Wݒ�z�=�1��{=!���*-�@7]w�[��Py��LG2M�Ԓ[Ʈ��ņ48cTO�v���W㺹��3��#��b�������
�V�H,/RS[G���V�c�o8�	T�|�����T�Yk��q�td*�׷������5#F�P�r�Z.2����m�y.h�����A�-հ}j�Fd�#6o�����_���r�Tt�R��Cx$;<)�	wf4���;�l�z���s��U��������8��\ԉ4�A�j߃�~p���?��so[���ʎ�Ӟ�_u�c:G �2�O�w�ѪL��qT�T<^邷��2��jƊ�
p
��T�4y�w"�|��K s����d�Y�Y�X/�熕�G�BC��� �r��:�!�n�*z.&C���<��hn��Z�Isy-�6T�n�`��{����5N �F㔌�P�^l�Es�a�}3e���"^5������`��\u9&W�B\��X�g�y���h2fSay�s�'��o!N".���+U�"BYx�����P\�-�<JD�%ճ��F��R�0�o���� C�@�!\�@�����m�TS%��X����M���ij*�ͤ�6��l6x�r�����v8N�Cjo0�N$=F��������}����h���kD1%� r��)�$:����A��VҊڷ%�{��C��g�n7�N %t�@[��~�&b�
`�Ւ:)FM9j4q��hG��P�E���.A��1B�q��P`_��zbm���$�����p�-��"��B��T>����r�[�d�BQ�ǷDbl�#�i?j�
^Y�R�I+8ƣ���{
��XM����1!�,]q�������%���|0.�/ld�`{^ Q�!��Qf�J"��AL�58�"=E�*�zмu�Jԛ�D=�z��"c�����>�U�����t���}�� \�v�M���3KT��@�<�c[�n�i��K�K,i�W�Ѫ�D���T��ʾ�,hw6ɩ�\!tk��9�:=��ג\��J�{�w���]�� t���l�%���U`��`�WaF�	dP1U��?�'pȀGv&��ywM���4�*� �a_�;��7w-:���{�^�eѐ�l�vt�$c���
q-�8��~졔�S@��?�w���*�5f�\�f�H�9\��H��6�B�
�Vɳ5���d���mᛏ���9��uxJz���.}���iT���������p;Xm,��/�m���}�!���"8�Ի���>i<�/�����ߙ��PSךU����:ô߮tNx�Nu��=��"A��G *�~{{���PD��p�z`//W�HD(��?�k���7����V��7L�
O�����*�$��NL��՟W-O��$ȣ:��1nl4Ǯ��>3���ݸ{��BF�M�T!�f�B��g��E���Ru��g3yǳB̺�[>�"�?���d �(;�ذ(�uQȐ6�������Z����`�(��8�x�o7����(��J/Y���=��h#G�K��:����
i��P���d���e��lL���ԭ�7�Iվ�ü�U��
8�?�� ��J�Y�ȼ
o�E�
ݗ��f5�b�g�*'[=aj,�d_�1ڭ�Ĭ��ґ��1��� �⯒HT0�v�Lc܏ǩT�?�9|,�F�I�����p����׿$�/��{���=�7@Mz�a $�C�N:�yd�VE^e�R�4?3�CQ�ꗾ)A��)�'ƭ�-�{�t�x'`}�� =Q����G��f':u=��<&��x��1Α��T��wW���˶��/.A�4L�(Ƀ�6^�H5i���&=���q��ҮI5�od0���"dA�P��'��mTM9BV]]���q�j ��a)R��c�N��゠�D����� 波4�_�V�o�Iocf�f���֞���	�Y�_�P�Z�e����э��<H���'Y�1�뎝�giTt�ҩj�^�/ŒIb[���G�9�2L�}�HvY�$���Y�XD�c"|��0��{ ��������V�g�|����RV�'K��J��C��T�ܟ�F�d�Zď����>\{�i뙞NZ[.�l�~��ux�V^���<�<N@�nc��À+�v~+�Pk���:�PtBi8�����o����E^�B$�ŭ���L�h]���x(��TH��zex�pH�Y>��k���u��ɹv#x���T�\V5��@G�ԸX�v�h>�d3��r[�ؐ��y�9	�����ef�n(Q�_�ը]�[��ٻ`��茢��@L�Կ�\�����"F.%sk|���	��)��KITb�E����ѝEmɡq��ǻ�]��������5�P�v^D�2t�[<�+�O��'=(�_[�	����=��Țїa]����wf�2�.V�1�.�3��c��v_���ՃfP�)<��a��P��^�
�.ǒG
����X��q��"����*�e�t��>�!:�}�'�/���
����kt,����)����%�ę��߿�,F���Y�
Ϸ�qSo�'��u�_le��cu�n�yu~�g*7�I ��?܋@\��,0CͻOm$Y�'2�49��e�N򝀞�%K�1���oi�p�~�^R{1�+l���J��Z�>�%2�����bֵ�2津w,��/�����!GM���S�y20�m��N�.?E��w�M�K�-����H6�-um�U%���p`J�Z�m�C�<��Aϭ,�Lx���Rȫk���L%�=�盾�&�5�f#iQ��UɭGD_�=���{ޮ��?�e �܈_U$b���@}�b�n^n���'�io�T�e/��|N�=�g@�_z0�V)-as��I��_/����<�;h���ѳ3�)SO�w�e�B�PLw�J��r*���D���b�Lؚ���i_f�+�!ٸ� 1��	�1���M�i�R~w]m3/͆4<a�l���{��J��?��k�7|�򷍪y��H��]�[�w|(�Q��H6d/�{��+g}�9�0q�G]Lt����:�����tK�.U�����6��(���n�H���U�:*6cU"���ta�/��{��؏�"���/�`�+�@�O�jgn�$-o����7X�����@x��۟�R�#�E#�k�!C��E����9`�XoS@������D�,K�#^r�������'K=[��/��P�%���-fk��;]$�1�D��?uC?,���݃����P�%�?�(��r��G�#��bJ�����):��ql0�������2/�|ƃ�o09�����yo�I|O���j'�y{I},�FP���`�9�ZH��������}L7%���p$���O�����
(�^�J��K�ބ<�hN����ͣ�q�ұ�:+�`0�дh��?�*�%�s�kԉԸw��K�"���c�g���������@Wp�����S=c<��܁�yַW\��w�����0W$����gf��RSW�H��6?3�Ok�Ղ�db>�j_G�<w��W���d2
�@�7��ް�36����'x�eF>�
Q(o��#��q:�rH�PP��i��=�@q�rxn-��7�Y�U���&���^b��3ov��.�/��0����3��ů'�r����*/�OmO?n��V{}��ms6|�&�� 7o����|��I��=�u���["�^1�����ނ����{P�s7xo���M
�y�MG�v���T�����plN�.V��g*�Y*�I��@��0� ���`�b��sW!��m�c��d��S��T��>Å�IX@�±~u֐B�����1���%���zPϝ�^��\�V;[h쾿�f�%
���4X�]-d�g���G=��)�<�
	�B)K�)��f��JԠmA��I�Q�@e��h�-�N��ׂ����r�b�& �G�N��x�Y��V}-B��.3%xb�e��r�  zt�V����D�>�?H�J�Y�MW4y��d���U͡?͓lA�2���e��;�Z�]�ɶ#P�mP���]��*��a������_���~~��{c�FW�b4Ƌ�%�8T^�&�m�Z����;��}M�d�����Y��a��c�Vx�LB�[۳�UB��yw a�zΦM;+�<M���ó٪"�Q{� m ���Jg落X�VQT��ލ�<U>WC1��_ه���)�5��Lj}	�8��AGh�
C��q�\{��Sy_����{�d�5dF�B)��rЅ��H��Du���DX�&�d.~����BL<"t�.�
�nNI�@Sc4I�(�9�eRr�FsP�2d`Ol��C��lm����(��(�k�������q�ű�'*5箴Ɩ�%�N���3d4��PE�Vڬ� �~rw��L�q0)�84"ں`��"��ʓy>\\�3G��Z#xxE��OE�Y����kS��a���z�-?=VZ��l����۽Ӣ��N�U���܋.M>�W]r�RۑY�H>i�� �O� ���2��'����Y�fl���!({�մ���6ym �2d,҃D�o�kWM�Q�z%�>*�R60q���`����@����=w�]�����׈U���;���#�f�?���'�{�?�@ ��1���*.P�:�À�s,b�ǖ�]�-W���X�{�C��(w|"�W��|�`Y:P�gW֊�:^7K+���@��aq�w'�.�Ƒ�<ҕTO����Yp_�R����+��U�i!��U�C��
vs	�.������y�>�"���g�P��l#f�1����qV��N�ܿ��:�!`1���Ņz�(h���qs��W@þ��fB;tΪ��LÈ�B�0i�),�Sh5V1���Gؠ�7�KW.���*3��9q9 n-�SC�T�7�֕0���W���su�E�BSr�I�KOP�����δ#�y;�P���L��Sm���郤�࣏�$v;�i��+'�����Q�L �_V�,5�4�*����!� ���d��N�����)qr��잙&ƍ�7��I��'��c���L%����-����J�Qo@ך�V����IK��3��A2�6��5�h7d����O�nY�|��+}� �uMK)��╻�v��z�y4sX��M*֙F?6������g!�UT͵���Ba>��<gΫ��Jc1^��}�R�Bt�@�������6�H���ma�V�`�+��;������O��C�6�/��.� �nl��0�2~7�V�tIuy��g�:�H�Q����IP���<嶎�j=��g�j/O�~�ͤgB�r��������*��q�,k���{X�rjm~�E����3�c�X#�3�HQ���I:�Sɱ�*:�Q�;-G�ˁ�j�"
��;!��/��(�JT�xK������J�����Xd�][��Ͳ�xqQin�� ��VC��mx~���䌀�s��g�F�U�\�������ʰ@�!�A�ͯ]aGs.����*>�5��7�M ��g���׾���A��`rČ^b	�F�}���v���{V����>����Ԧy���	%3.'+cR�HH^U���`��h�By���ҏNi^YU�)���Ēm�����H�e�����VG=�Z�`�o/H�����M�r��XR7��tj_����֊�K�KI��NUڋ�q)�{oa���%H|x�܀P�o��{u����^�$C}�.��2<�������[��F��4,3������Q��r�x�aT���� �j㌥��{�$,�&�ê�����q��,P�*�Di�M��pYE��d��1o��*��yi|��QU��o\*g�/�\]��`��p���4?�8f#=}6I�qZ�[D��IK�C�h6QX������֨��#��K���x}G�N�²5��S��_��2�L�	>�h�~��.�@|pVxK���|N�6b��b9�ŗ�����4haڞ��<���߼7��P�����i��UKq7��uJ 5����y��9�l�*+-ҚHh�c 2��q�Pb�^{�u#�/cWl��?+���`O=q����<�YQ��y��,�Aڝ����5ʷ1,�4�I��}w����Ɵb����i�Xj���N5��/�T��t�,���\�8�e��:��,Nj�D���
�;(7���o��x�:�`�&�n�&��[[���"`�<�܀�>Ҍ"������1�=���D�e:���c�?�����]�n�\&�FF��oZ.�;����k�(y��,�k`�]�����{Z�/�@{��XU�|�G(��~!��@}Yքa�X.j|<�|[��vm��(��gM��v��wU�p�j"&��J���B����G�u�" _�9�=5��m3�j{�<�ir� �{���p;�E6�?���/����ȇ�d�b�].5�M0�5e�p�g�>��$����=��}s@� ���	��Jx��G���#t�;�>�����C��_쭷�Q�K�ߌ�މ��G�O � ��< ������m+�e � $�pس�xV)>;��-��a��ihhe�Y*�^�J"w����NK�"���^����ɣ�n¶��y���!����j=�C�f���~L�N�n��U�ۆ�3���Q�UF�$	��҃�`L���˹�D�FL���A�U���d�2���a�� s*܎%+�>{�0b�k�D��W��O����2ݟ�ϔQ�9);�D��A�Z��po{	�)߆��>�(��a�^We���7hض$�_b!
�w���"��M�|����\ij/8q��g�1ŐëJҍ��J	G,3��1��J��9�p���2�^U%BoP�J�iZ�ԩbL���b�b�@;��z�`���<g�OC�YmėDS��nVQ4ݝ�<���d,V	�H�C)�g�������O%)۸�{�!�5$�������:��Z��<���R���k�za�w�Ģo��E��nw����gx����l����ڽ�U��^ѡ��Aն$ �ͦ��^*C��x�tYe��#��&]o*B_u�VH��XᲣ��W��R�>1}�(3vS!�EDj(U��4�3m��'Y�-�8+�#�� ��3��l!m����iqa��0�=�Ǫa���1o�w�˗��)}����P'N���bя��n���<*�c ���R�w��ڱG�_#8�G���܎Ee�kI�?�Z�� Ņ��]�ۭ8T�I~��/������*r� ��K�{�K��F��."X�cw�/������t� �O����(L�w��z�*�g��oZ@�Q�s�T�KO�*[KU��	3�����õ�����O(�'��9k�.��ai��ɋ��N� {nl/8��£	p�[��TErC��<]�SF`��~����!�+`58�b�����'`����WzV`(�^KV��ݢ,at��m����<~�JY��/|��H9�YOC����w#�)��{)Ƹ���p���,H�W] ��Z�=�j^�_J�q,�rG��=�CI4뼃�U�#� ���{]��3&v�N�瑒�����q����%��>��7��uE�x����������N��N>ߴ� ��;�gTؠ�9�0��W��OZ��;-����; ������:;\-�Ε���zsNn�]��|Ӥ%%u>���F�͜k����m���=R!�J)ج�Le�A�8�,�m�XrS���C���"�� �,�+){х�u�����\�S��$[w�~���Ɇ��a��uyG����o�����7�2�`z.y��#>ՙ���C
H����+�/��]�,�#m6:KDӠ�'A�Ah-4�H�b����5��5�7Ej�`��l����`�"�NS#��Zɠ+�=f��_����AFS�٢�| �"�lj^�?���B���:���+ʐ�&P�t�����&M�X��!�=�9�F�����W&���*�����[/�'�Ȕ�}2d�/"�W�D�"qv�W���NI��o��;����xӵ�����pm! ���M�L\c�� n�`m����o�~��2��@��NW���)ª3�[|cR��ӓ��og��u+�t��%2�~��7�-4�.L�'r� X��n
�w$7!�8h��;�y	Uir�Ƨ]YW�ڶ��������Q��lY�6ޕUG����Ykx|�^���=�	�!IK�lD3�Q���/��k�QA�=sR��m(�$�j�|���o#�ۙCea���}������uhT�W�B�@ץ3�(Ս�׊�q�\�e&�49�&j�VA1~g����U���B�8��q�����5�q־��B�"����^�IȔ���q����/�U��
-���>�f����f��M��6:��w4Y��'��mH�`���b�a�ʡ�}Zqf�����-�-e]j�:'��*]x%�Ϟc��˸Q�)׿�aSm�cS&z�&����p�n��03U�-)wCm��}�'D�G���~��^2��p�����wE1�2����܁�(���T!@�|o��4�����+eݗ�@�	w>����a��a�'+K�"pd�Qh=Ȍ
���aC�	k����/7�v���:���͓O����5%��K�����(�x�TB��Z�:���g����G�3�C��Ŋ{�����z{>b!a�2V�=�6����֋�	/��+FL���"䃀�|s8��� 3u��I�y-94ȅ�)�:	tx�H�d��F�uV;N�K}�u���b�J;E;���[��<�89�\Y���9Wײs����&�U�W��XT�6\H�UZW��3pxLRg��d4��;���E%��R8�2D55��M�4����q?����ד��/���Y��M-����"	u�W�^��{!%�b�-�Þ8TMxM�C��q����O�k
2n%k�y�Ҡt�0+�>���G�ǋ����2��w�+�~2H��y)^с���(�dAeyI��B��U�w��ʑ��~ͷOZh:�2xf3c��ʱ��A�> �HYw��A���Q��r�����<7���Ŷ
�z >�0�ѭ2,)ѦP�Afc쳱ﱻ6�^�����.�q���;{�z��9Պ���C]
|p����.���3���@�⹜��M��A	�H�ϊ�Β�!�}�q#�������܄���&-s�?BX1�����G)"w���������;؀:{�1!��B�e��U��S>�`V�гţe��"�d(�y��7�o�B7��"K�}N�a�.dR���y0����|��([*e�.�SO���s�tWc�U����U�˵b������ز)DcߎE0�JJD�̼�\�A����r�����p���?%�H� ��U��w�S�W'��E��2��_X�k�Mp��Y=����^BÐ&�a�=����@s`m�Cq���w[����,n��=L�{���&P�"�*ύ�1�9�#��iT��ƽ���O��{T�������_Ȋ:(���'L]�}��r!�4N����
}�f>��k�~-�J��پz	g�$�' �H��TϮ��M}��2����WYe��VG8s�&�w�g��H�b,Rn��R���cm`��%_�6�WQ�`$|�
MB���Ƴ ��m�����]�	)���8�����E�=d���V-� ��m�4�ٍ�`+�|U������@]VR�U٩V㙣FOؗ|ۄ�5�BS�P���9��B}�L{ށ�0�dh��9��67�"Ne.�f5�0�_�55�M�)�(Õ1��� ���2�����&;���ų�.w�wx�0]�-���S��K:�y�����AO *��c�b�����H�@�xޯ@�x��_]���B�"����Ա��@b�hp̈��ZV�T;�μ%i��jT��r]͹�K�S>��A��|:���w��6�3���
�GM�6����֭�cV)���@Yo����q(n5�7��o�e����g��f����B�a�B��JE��5���!(�.(���d18Ϥ9,�߅zi�3*j�#�b���ͮP��:�Z��j+�1š����(����Š{�GI���y.������:�R�I�E.Hy�3�*&�l5��E�B�V
1{�n񲕭=kp�)�E��!Q����@��e1���/�3I���F�L�����yv��aa8��6��4��¦_��T�hZ�TOY�*��|n|��}̲c�&����D��Pt��P�u�͌/����w`]@񉮿Z^~hv���OU��&���(fR��1����6y������Vz�"^�P��P�I�څ.�KR��$���^�Q��oLnřB5�y!c!�)k�0�J�*����%�l����c5�0=�4���hу�Ц'������u��Wg���z$�8�xݑGo��p��(_�N�,1J��Tz1���{�E��K�Jv�NF`���i��ޅ�e�iK!.��x�F�o<�4�,.����&ڢ�+�:9� �	Of`cx��?�:l������s$�*N
�~vxo*��I��9�h�d��#ww�����t�v��Ot%��U<�"m���"78|]e���\��G�!&WX"�2S�F�A��#�c�H�v�5�_�{g#��?.zP�j+��� uE�?*4cEF�ZFA��Ut]��
;r����O|����,��teAQ�� �� �� �3��цx�<˷�Pa�%��A�<�i��^�0�'����$���>/>kj�mאI-��f������	�����' ���m̸,���fS[�P5�����|�7�K����8=���8�6	��Ir�g�wWƊ����.�,���Ӗb�MB�t}�4t^�Xu
i��MU}�x\�+X@�e�b��%q�d45W-���јB���N���o{(tIⲺT[��=�-Y͆H�?
6�y�^P;�g�'G�����*���+��]{��b�H
�<@�b�4�:)	����f�,�Ɯ�$g��%�/�װ�x�p#���E�vY�&FX�Sߓ�	�� ?63��˚m���a�����@�'6�i�Xn���(���\F�	]q�.��G����E��#�2���놎��9���S\MP>A�챐�~D�d��zA��5��dJ�
ru�@��\.�����U���Q_7���; �K@�	���C.>�%�*�|��v�m�RzՓ�o3��n�u�F:��]n!��uR��ϊ�r2sp��[2n�h�;�c�=��p��k[�ʈ&6���O��������j;�B�{!�~TrMF�]'u�>�/z�Lm<���H�kɽ�[�=�S�����b��=++DH�����a�����cw$AZ�?�cc���7GҊq�B�w�s��PA�i,�j��Gb�q��I��wT~O�ă7<U�b2ⴀ��c��V��䭨�s�#��u8�r�9A�D+��9H �in�:ƌ80ѷ~���1ƽ��556���`�V�`��|�9��K��e��+��%�<��^f����
������'�]�R��!�"/���1sd�%�U��`��.M���'��`�`��7���-�������I٪�x�g��t\"+v݂ ��/N�Iw����4���
��&\��|�@��~Q^F���7�7�S���r�8�"��{�f��
w��
�#�f͛E�d�<l�f%�������`7y�I+�
���-�τ6��ɽ�7�rA�i�k�~ڐ/�x�����qC,�w@��͏�D�-�rW�s����Z��}#���)#�N�t`��,� �o�eD[��Tz��Y<��
x`���z��/>�7�tNg�N<&YV�~�����P����L��`�K�74	�Ć[�Bu!ot_]?Gz�Sз�p?��.���-�=��u
k���m6�N���8�S� ?���Ie��X�p��Lj/4��5g�E�'⃅_R
�3DKf�D
)�,�,�sˉ�-2���*�űW�DrE���&���̪:*��)���頺"7�M�M��I���[��:��
ݚԉ�vbє����o\8y]3����5/���_L�C��]w�	~�$�_7Ob��;=B..?T'4���Y�d����}l���S����[ܖ,/@|��M���(��I��EA��������D��#��v�b2�кn�c���A�u�6��oK�X�F�q��^c�7`J�$�6�.ƛzJ�kz!U�;覚&��OG��4_���V�g�-� �G���$����o>�,S[ �Fe���yڕR֑&�;.���L48��0�}�m&�k�����'rLUB��b��KZ�}&��ZE����R���Q����퉩����%���π}/��fA�y\E�&��߮���!{�E����%� �"�(,R�_;����'&J�#H�el'/�/���/7og_F�>���H2aF��\��ʉ^w��P�xsm���W��ք� zk��fK�PV)�j��E�����8��ӊT�R'3����L$���3�h��Xz���Ļ�vu�@���Ӌ%U-����v�&	<���W���j��un�!�2L�K���9�L���]D35o�����q�6�P���1d�l�f����$b�v����/t5R��@�֔�D���߁V���t6�G|KG'���	�}4�vүu���˵��[�?�-I�����K�A�4�w�G�:��ϠH��F|�&#
�c^�-�p ��q@MS2�^���2���������:ku�G��;{B�����s�/�Q���x�b�D.��\C�CJ#昒�^��7֯�pϏ�C� �j
��&Y,S�����r{��.��	�@�fu�Ci��m�{�ҨO�	;����H0I͇>�^�)���s�nt��B��V�Tͫ�02��]#BഓY��+a��9p��X�hT<eL���p7�S��六ȴ�#>}�ı��t";��gGV�8�Q������k�XQH[G�m!��z.�d��Ř+*���xz��$#)� �����<	B ɜ��;������i�W�b�����C�����щ93��kNc�0@O7�,;-����)	+7�1��/u��DZؼ�S��k���J�I�s�����}ld$�>Щ���'��L��q$�!d�6x�A�<c�Υ,S�OĵvY���K��}K����������R�.F����g��BP|`u����-�I�U*e#�kMV[�,{�bd�>�;�S�OU�	9����&�7����s[���F�V�b�w%������P�f&/������gl�o�ZZ&��Բ��<t����ǜ��ҝu#����
��茣�����4E�3ņ�L��מ�Y�:��&o�a/K�el���5p��BQԡW[4�@��7��=���5	�.dԧ�Nz�S{;��yD��R#m��%6P����Q���u��� _e��3hlE�3/4(��p�&�h�|�:���Ԋ�Ĵ�+_��l�M�D��k�3x|��b������]��5���ߏ�&��l>�d]#Ԙ;�I�"�c��<a:�x��
�G�C6>����!���!���s��<�A���'7��p���ÔT��[`��M�-TJ_������'Y�������?F��-��YK�����Y�p��`��:d�"�S XZ+o�}�������1	� dΧ�"���ڟ��(w��5Τi�緒�&��I+��֗*Y�ȊȻ��7�� �n[�9踞���{a�$瘞��7-��&=HTa�71(��;�n�J�&���+Ѱ���M$�����|qEѐ6t�
V"a5^�R�l��7R���聪T�3b�����A�cI��s�:ų6�ڜ�be�X.@.�q1xˎF�+��c�eR1QT�/|���E��m�'�f持�y�'�f�:�������N�06��%J1SL�����#/LR����:���Xm� 6�,?���H5Z��$��<:�*@S l^6�{����3Tp���@���2�Z��Y�&��AkKrA�V���n&U%�n 	Xa�h�����n����wBM��wK-Ǉћ��oPc�6ݒ�C^A��D������W����f�h�HXǳ�@�=l0��7�b$3�F"qۚ�aǥ3�zb;����������#@���AoWtaN�L�`�权I�劬SKL��*�����X˜	�1�P0�9�|u����Z���__���W(�c�g|��j���W����8�`\H꽤~H��Y����e�?^�z������2>i+/� "de�2�-,	`0w�.)���������H�]B�~L!î�߼&*�X�E���rad$��E�*۪��[}�}@��!+#�E��s���:Q/�=�~�( �!es��c���76�4�x0�Ζ*�����C���!�#Ⱦ�t*�I�9ʦ����TkXg���=�w�N�?>PZ�q:݌.����^��ḁ��*�� &p���T�*��=�y �4����!�*�Լi��K������y���.�)�'=��^���pF�o���1*��	!9u�瑑�1�H~��z�k�+�n��7��wP�������#.��X�����R�ƛ��.�C �X�4U�B�ޱ|�Q�2]�~��Kp������r����m�W����t'�6i���=n�p*F
�p�)�6��\�YI��1�^�Fq�_�a	%��$�����n!��ij����A�����|���MJ�쵇�n�%G/5 Բz��1YN�]��,0H�R�Icg��l�F���@qԿ�Q�uD�l�^��[�Rԅ�!�)x��|��r���-����W{˂��9w�(b���zg�n���*�M�mrY/|;����+X�C�����_�b5��g��HGf7[�T���;�lYo̂L�q��������O��_�'I�\R���ց@�l��@2�A��P�G��K'�߁�82�@u�i9Y���Ī�#3�>�����J�7�R���/g�(<6Ha�!�l-�[������KdG@2ciE�y ����\���}x��N�h�C�i��x)�n�7Zm.�Jh���8��y�vV|�Q�=����(P�\K���W���a�a	@I���%�igU�0kr�Gb�[kE濫/�H�w�E�%���Ϛ�>���F�6A�Q�_��'�v�(�m7��'�m�$��Z���լ���b��ϳn���ɰ��S���(GQ���(`dn�C�\�5�^�	�&+y��A1h�h��O�S�����00����qЏA�C:��o�&F���{�����zW�s�Ꝃ�R�Xh�sU�~⦇�^����R`�w���,r6�k���-��=D^3�v�6x�nP�8r�1AP��}rKi���Vw�\��zK��վ�4?��ZsG�=�Ku�!�n0)�f�J緪�j�ɧ���k��s��/#7����&�vJ�(9���J��.O��P(�e���b���k|�d��	������4oGHubj({ �[������%F���xk��1���tV�/�dg�#�@h��_b�Ǆd){]v1E�:��@S��-�D˕h��\ w���<ȸ_+�	�]�����5ٖE �{��u�mCV��r[��A�#�l{�l�-�zy0f���<CF&��^�(,B���q��I�5��]l$�4���ܩ�&K�����LT!>���c�s����3����ò:����xw��_'�����8f�>��<	᫭J�1�WC���z�meUR�xl�j�vKܷ;e�����I8H;;??v<�r�=�6µL�u��cT�S������,��r6v�m�R\�~�&�=����^�%��/���O���A1+������{��D{�����G��p��)��5
7�K=���^,$��uvXh'P�;�P�0dp�H
�3b7�:��2V���v>�8�$a�{��@������f���?[w�MyXy������|�*<��Cic�Ņ�W���y�V�%��%��\��PG�bW}Ɓ���/�4*��<;�s^����q�xC��uϏ��i�������a��VO�!]�v�E�{1'�������w{�ņ�z�;0q�?U�bk]8�Č�ІQ���;�1�2g���L�q� +������#r�t����&��W�G� ��]_ipv;�V�g׌�ߵ�71�m,�,��ϖ�gA�7Bs�/��h8�I%Z��x+�Cm�����\����{�U��M���)j]m���C�Hp�:�� L˲�C��зj��-j'��+�Y���@��^�H�s�� n����'��Ixv��ǥ3�D��;d`��"�����������3�� ����sp>�M8�����?L�$�YF��j�|�Ld#�X����p.a�C9�r�� C���d�ٶ��U�A���!K��Te++#5�?M��B� �K�)P�:�d�L�znuV嚯���s�5N�qj�.�r۬;��(�f�*p�?�h��1b�TМ�D湐�,t�Ζ	���&��ޝ+I�ܹۍ�*�γ���V����Ê��辞=V,|Av�
2��~��e��#Y��������aYq�TM�.��K�A4��DmLCY�[��k.�[%s,=��,W[H�Xt�x`%w���":	�w���ೂ���s�,��*�y
t%�g͗l쟣�e(�T��w�}og �*t�������0d�NlH��ҝv ^<�J�e�Br󮆶{�Ҕ�9`�O	�e�T�S�&ڕ7�t�J�'k2�T�_&.���'���`&c_8>��`Lr���q��5�'�s:�*��/����μ��	�8�/������bLd<X'��\��D񟒥��]eIe��h�V�7	��u��\$l�-5ɦ���.;S1��^�nv��+]X����^wDy�����>�� ��3�d�_J*L��o���H��i2��F���>#{��a��8e����o�
IȦ�bq[t2���,Z��|19)�<�����FN�����&XW�s�'��.�g�G�]³�M6��$��.�õ{�%�-��,]tE肛�A���+�����m�vu���b�E�CT���o���\�VCy2t۳+�M��UA��Ѩ뚺jI���������`0���)"���ہ�(<�6EU8}-@?�I��"΅l*)�� ���(��z[^��X�sD���'[>G%O#��yOBR�����ޠ�lq`��!��|�QR4�x�<,�2O�ܰ�~g��eu����0��2r�?K�H3��.vz��9no`�r�nS��XO�qy�v=���y̩qß�;��|��yb����
�t�ա:o@�
*	��6�ZJ��1P�()*�����H��}�X�����$Ό!��GGA��1Y/� �nw9I�-����+'.<69��S5aC&-��;����sr��G����N�Wq<�2Ĺ ���ǆ��5p}�+𩛄t��b�g��o�9O0>��{��R<7ώޟ[�J.�Ϙ��$fƼ �7��{m/�*��GŘ�Y<�R�����[�
hl��B�����7�s�p���x;�v��W�-������-�j���hQՃ�cN�xj��o����轗����p3���&#��e�h��Dw#� ������w�zJ�^V�D�z��d^~�|�$�nnڈvH�R<����[-���Q|[�e�0�_�pߕ���M �<!,Է߇�BU��9���f������un��"F?�0�K�c�;/�L�4� �Xy5�xw��Oi���BB���9��Cn�UDN}:p;��.Fp��D�Cs���SL��I�'�I �w x9(r�%��7�v������1������N~�,�Gs.���hBE K�`�;mn�Q�^*k	9њ���Єh�g�#�|�-;#R�nG��V��3��Z����N��*��8Kss�I��F%��I�6{���+�Mn���s�`�	:�-D��1J��i���K,=@�E7�>�r��)��z�7����!gϻ�T�E�חc~���l�t�:�U�/2�S~IH��m #	j��dl�	Ґ�]�k�x���/ʢ���(=gtz�^������pX����0=��\�d(���rx�Wf�A:��=UV��F�B��1}ь'�D v���7#��/��{|�do<�~5�7��Cs�l�S9���`M'w��P.ǉ>.�`:����ՌI�-��f�PZ��H�y�Q4�F�=����2�#?5[o%�ƾSS�j�kT��C��4���/�;}~�{���O�@��Π<�%Wn�M�"��Q�y�����=g���zh�����q�-V�i��П0d��&Jh��� ��x��	B�ohN�ˠ�;��NOy���X�ʠV����)}8��G"	Lg�쳊H��VUrp�*kv�/-q~�:=]��������3��2\v�@5V	��|�:8B�P1�ma��A
RP�{�5"{Fx9�}�/��#kA/x�z_�s?&��3�̘#&�����,zsX��׽h�D4�MLd!���F��5~h销8�k�b�%�F*r�J����[�]v�#����T�ѳ���Ay�0j��0���2%:�^]�� l��i��m�Ј�w|�ᴆ�e�w`��2��s��WӠ̌.�'�AtY w{��[�|�p`�6�*�%����B��j�TRX�ށ��t��s=a��vt?P^AtD[J{6�s��RqX
�$�
����w�XRG\274r���y�-[��N{.Ap2�@���"�[�y��Bk�?��Ꝛ�)���ʮ�5o�3��8�"�H��N��O� 2��O�yb�d� wؤ��z?��NFr�^э|>.��pu4�F��D+..�3r+	2��| �F�����ϭ��c(/�2�'*��)��s�x?B{��ف3��?Ă��^?:�:*SL�^���?���#�v:�tA�'U7 z�b������ғ�%�$��i!լ���=^��T���_��o9��_�܂��-��\;O\�-<������Z��R-䆄]7�ܼ��V�f��mJQZ:�"3�Q�N�/z�*�M���$��Cݯ���l�h1��	�u0�g�����rGc�܊���<������C%4�?O@��i���H�N^X��YdS�0'v~�Q +�$�X�w�cqVt���!�`����5Y8e�Y]�G2ɱ�[��݊v��{�:2�24�V�xWI��ѳ�4�.����~�Yzn����I0��/�3^b��gC_e7B�N��hqW�����������N�*���ў���],.��E��D���q�X�./�d+�(�ͱ����?�ı�{�o�9~��	��x�)��W\~���t?�f���| !\3V�qc�������n�To�S����xҍH�tP��^��j�o�A����!�k7�u�!m��r���#�,�o��gt��0��`�K�'_{I�y�(�_���^ʿ��|jBk�v��Z�ڋ-ͮ��T�.�ak����m+R'F͍���B��,����{��b��Ã��T]ZX�}��d��[N�<јh%rNGi������>]���V���,�������~LF��(o*��z� F�����8�b�v�QT"L�/���D^���9]5gm79�I���z2-���S��+�7��;�ͷ�8����t��U�v�WK�Ǖgc�Vz�vX�Z�b&�j�Z��q �i 2�6m�r:�0t��!�|ܯ����1�&�ao����G"=w��ޘ�;Sh:TX���ޥ�Lt�*�ǟ^qY��=�hC��1鹣7��I4p��]e8�5,��$���$��)$^�i/��5��]�d�`����Fq�AY�܀ IG$�����E^�L�(r�01f�g�7jd ־&(
��Qs�����ޝمW4'YG�y޹a��&�7E��i��k��0o���<Q���g�ۘy�.�2I*i��?@@����^�$�̣}���P����FvMjA���Ņ�a��+s�$�/��6��r^�ΰ�zֹ/P���
�zq�^V<"p�8�;�}eDך��\�91?��]�߇����5s]��s]��P�zϺ��l�&���usR4�F{��Xcܵ5��i�J8��0��v�R5���W�=���z��r�R�hi�ML�Lu�h؛�;ö��؆�$7d�(6EO��� I�Z�<�D������܎�%��-�6/M��c ����i�wen=UA����nwә���h"g�j*��Ŧ�� dF\X8���bߎ�3�����Bm�ڎ����sX��'A��!���'�`/!��L(�х�Fӣ
L=h� ��>��p�t�Azq�Bn�#{C̼HY$�ھ�7QfJ��i��Z:5�g3: �ͯe �+��ZU��g�������a!���ɽ�6Wru��3m�����K.�G�R�\k��[ѡ�YP+ ��<6���ಙ�z,��.�W��wҾ�W^䡻h�,��g:�t���_�#K����<�`���|dUi���2F�}��!�/�Zj���<Wa���YI�EL�{���B��Bl�M5a5�e�<�y{�UG_���	�J�k��\bF�{G'rca������ݾ
�^�2�i�gq�k
4�i9IS�G��=8�Dn��I+xh�P��	�j>�ب�g\�������?�����Uo��|�M�գ]ԏ�ff6ֺ����1��ͥ��Ε ���Y���{n���k��P��Ǚ9?��B���n����&A��]���4�`at15�A���t�[�V�{����eI����i��7�?�6�M�����x,��m_+�����U��E�y����?���SO>c���dϐ��76T��]t�	5�����4��%�2Ey �N4f�F�))�'��M�C����A��������:p��p��O�z7 ���Lr�~�FeG9�w,%��}�eEr W�(��Ճڵ��:��%��K��`�oY�v��������0�FZ'�t�����<��>ӊn�ZS�;�����4$v�ӆ��a�c<�)��Օ���}B�J��jmjj^y�B�`��6{� 6��m�$!M���E���Љ��I����<Z�f8q�j!���e Й�-��,f�inݦ�����4]o	x��o�u��@��Q�եA�P�c��S����KER�,�j�-�SZk��q�=����,迺����챷M?vXq��e�&p��o�W�oQVy\�Y��sx�;(���㿫���<Mc�4�����E��'����1`|1�3Z
Wg��N�w��=х�8/2�J�6jGFֺ7�� "�%�3u
B@�AO�Âo����V;�6H'�4����(i��hx���ȷϴI�8���H=')�+tTgnW�<�|�L]͍-�3�|��3�\B�-�lA-^�zЋd��l�T�Fʘ��wR�z���x_`NH+Y?��P�6�t�է�,�	}F\{Y����G�>����̦����*��<��{$љWB��}k��h�:\�5�����s �_?���r��P����R-��%�eN<>��A���75Lef/��v!�U��,b�@헌�0�c�s�!E��G��,���:��P?0ł���$��a�*P`W��Ae�M��ס���$����<]��mqUi�leRܮ:�s�қ)���,��t�HT�����2�j =xƾ@�Ƀ7���V�2��,%/�qI�6�A��U�S�&Psh�k�W/`�,�o3�A�T3��y�S�A�.[x9fϞ4�;�Bە�Y[F�A_U��_{%�Fː�2꽆����e�U�l�G��������Cƶ�q��U\r���S�f��q������n�U����adQ��t�Qs]�\2,��ȚA��.��A�'H6��9�X����t`��˪��ا:������gH���H6�E$��t�G�Jʄ%���ޅ� �Oȍ �.�2t�/��[�l�_*U�]"�c���zz��>뤝�s����|����$=6հ㗺G���b�X��AS(^�0�,g�x���|~=�2Nr�7g���@��x,�C����*1��S����r��J�eB��C���s���=D�I�8���`�cr�GP����.�$ �hl��6�����E�2���`)A�������b-B��IѶ��7�\c��S������n�d�Dzd�c�)������Z\�������Nԧ���E-=��@�"A�Ep(UG���~�5�������6��2!=���h�<st��s8�9�����А|�#ު�w�	��)<�[��9\EY���}0��[VN8	Bs�G�����K�R�*�â����)*XBSN���*G�4y(�9@�f�;@9j�����%��[�����ּ6�0��]EV������5v;�ݹ!��{`�?�K�<�+�+pQw�ON\�oO�
��͹(?���֥�^�-3�0^�mfq�$�߽��Ȫ�D��\��6JԐ�v^����?�!�u����Ǝ	yjf�xXЂ8h�Jg�Y�ۑ��E��^�����.D�=Zv�O�V��K}j��9�/m�v�~)����o6���RdÈ2\��?w�>��ۡ���D��M_�P�/��ǣ��*�X�c�F0Ga�T��~ a
�����D��H3�뫭6X�4�N
08���R�Q��O�ULm=�� ��y�4�&B����ѩkcu���ʵ�$ߺ@<
�Vͤjˊ�5D$7����L���V�=;g%�ی0e�E�Ė�ͷ��0Q��KO( $ S	��fnKNp����"K�zB}��t������W�\{d���D#�g8D�ßp�tCY�]����vb�.S>��"Ԟ�%oЪ�Lmb)����Y�n��7�^^�7������9�p2�&-ҠҘI����EL�-�fk��@1Z���t5�;h�"��b:��#��=[Pb]pPd������� �$(��+�ļ��RWWo��/:��B��!�V*��%7����ޕ�;~Î�2������/�;J6��TK�������ۊ��`q4uB{��v(���]�6LE
32Sh_��y��{j��%�LP�"`�P�p��ЭY�j DN��s�Ha˷9p��L'��~p����z)b��0"u<.ֲ���6���qZt,Ϝ~�����5���}������hW�v�ф@?t�*���'�#G	0�&�qҜ�뷚�_}�1�.%��6�a
n�|�ϕ�.��v_dۭ�S�Hk�B�f�!{&�$��9}���b-��l!b�t����V��<X�hhx�t\�Xb����k1`v�c��G�	����򉈷�6����	��:��r](u'�w���`�3�#�0�^�X�>vtQhs����#�8�p�_�*�,el�Ԭ�ve͍�M��o!�rW_4*��U��\ �����t�����¬�pEeȷ�h`�:` k߅J���_z�qݣiE�,�������̷������tR!lM���K����6S��Q�>�~,���.kY�o�\ۺ}��x�l�O��o�]�hg
߈������EC����?[Z�d(C�F}t�Ėo� #/]����^����ʯ�DN�D����%\W�i����]<�����ʽ���{�'�n�,�<2(��j��%��B�wF�9���;~}����;���|�b�US�X:D�y� 
@��mIQ��p��KZ�lV�~;{�c����3,�����˸�����2��w�s�E(1m�<sR���E,˪?�F2�>H7ld��cI644]�Q��D4����`4�S�"��$A���~���Ȗs����Ok�ERf��a܍~�@q��)��ph�L�ސ��� ��]dZT�nD�bh��rJCB%3��\0�ʋys$�i����zک�=�)��ʼ+��`|�<@���D�"@��U]؀�����#<R��8X/sz�1ފ�Z�~a�|�l�9aZ�/�N���P ��7�Q�-Uष�)�3�H[�D���QK>313Q���6�\�Ͼ����������z'�G�^aW���%�(�}�ɨ
P9�Cz�d����B۳]���>�sAI��9�*�����g��P��"%K?ɾƫB�_E��_�)���Vu���t��@d3�ǟ�&C���	Ǿ)�@�lyS�s�2��.�I��.������;��gN� %c�2�ī�f�0��7SWK���:Υ$�0�{��I�f�����.WCɶ�2J�`֜���f���͂�Ҕ<`�������s�ǆaR�=3�����y9�9S������h���	�����Va	2��,�\Ez�O�>��r*p}`�y9��3���Ȭ��%��R�J̽��͆^W�>�c�D�#@)��z\�-j�3�T.9j,|��sQ��߰�����y�K�\|zim~�!z���F�/']���]�Vn֧�gnEjt��RH0�����w��]���i�v�~ћC���%U��a��'�y2�i���ѲM�iW��`�Ϯa����\�e��V��r��(�S�DY�X�5~(R���*����&]5S����#��	 �+���3��m
��88�����I%�0T����MB���
�?��D��u��c�}R���]�5f@��I��_���~t��q��\�rf�E�H�'�,)Ԯ��D�Vc�^ �=�ۥ���f���8�E9�Y�����E3�C�!l�[~N�X|�����5Kk:'5������c "-����������RS����F\��切C� J�/�l/��M�R�>�0Jt��cn��L�ӫ�D��X��/p	��{��h���p�vb����|�#��:� 7͸�5���c_ֲ=�7�X Ա����b2SL͈�F��v6�r��V�`�GNw��CKxG;�����-X��AE�K�׉�P!eLҒ�͗}+@�F	��f�ɡZ_��b=�8���@�Xf���2)�����[��fu+�ˋ��*kB�o����<��c�j������H;f��$bC�F�\3�c�;�����Ҩ��;���)��}��EԴx0=���xR�w#Ƅ��|1s
u�H⯘���hE�LDpR�^�@�(�Y"F�}�|V��1� /�KxT��ﱕ/ڗ��h�$X�!���Z�����$�Y������F�f�ٽI1#��С�7:��۱����N1A��Ĺ	�)&��<a�ҝEVJ���ؤE����1Yx�:�tVi ���L�3��ZxI�6�bI�<�6�ѫ�lu��4�~�[�����R��e[ON21�zg����C�}B�]��Qa>��մ���G���9�߹�NYy���B;�SǠ=Qc�,c���ݵ�9����s���l����ؿ�]�]�L�����U����Z*"�v�:�z�Wp�Z���yơ�]�%��p=e�ޗk�l�=�� 7����bM�|:�|@�n�ة.���5�*&"����Y�
��Ηdz�)q.|�Yp,���/
Ff�{e���[b�&s��;F{�i`�y�݌����!��䥱��$'���Ur��.$���UA��6B�R3i����$(p�4��~J�9��q��6�ϓ�<�ܸ��Zڤ��iц��i�7s�\����	_ �2�� TzO�Ak�X^��9����G��<ʣ#ar�)e��,Cq����.w0b�s�T�w@�Ut�E|��L搚{�|)r�'��l�Tu�J���M�8�eQ�-��`�7gI{���R�a3��г��Ñ3�1�O0U�80�6�����qb��^"�V�� >u���H�3m͏�c�����Q�;�d-a�~D���P��H'�^�ɃzQ>6eŹ&���*���iHRJ|�)0����gc8"|�
J�xIr��(l���*��� ��o<M�v�;ZP�dbE�ʺ!�\X���وoT'��g��R�* ��UI�PQ^�N3��)\��CB�����A�j�t�Z��Ȍ]�%�/�_��\a�� ܠ�s䭀N9E��ĮSKs;vpI����`ݔ8X�R*�#~�P;�a+�_F��Ȍ��d���:/�s7��[\��W�Tӫ?C��>�Wo�����t��L���n|[�d�-i'8�����
���W�$�\����nM�`�a���������D�U�p8��}�*<���&w�md!�l�����r�M<��m�a=����m�L ��?�jF�`��p�h����V�تu�x�"�q�k��:<cAc��K���_9�,���!����()�K��?�\ r��J��ru|R���$��IH ����*���߬O�~�p���Ҁ��if5�{�ls�U������X9��(�Gq?��^�\ŭ9Ǖ�X�u��`���iݜ��uu�/@ۿ�MV��{C��^����������^��A�k�萓�@�j��8mVm/Xs�[8�2=�w��3C�/�k���	3���}.���̴f�ێ%�gG�b�`�jz#���G�$K���[��]���8��c@��x��U��E�Ѩ�O@"�!��/���)Er^���͍���!4sH�a�d?Jy�E����m'ӽV�ޑP�]�
��)zu^�n������.{󑵲��Y	��1�
(�Fa.�'6���Låt�ۃܕz�<s潼J�$�k��f�q�P�����h�\ģw`&�ӱ@��H#���۶��fF��om%6*��8	�(���c��~z5u���Q����X�T�'ń�� �tD�Suo�/�����m����]pK�k��N������������dr�e8D�/(��6������Ю���� �%{��3��^]� N��>�9�+͎7����A��NQ7��S�s�`p�N�33�.���?�j���Mٻ����ź�فM���n����A��i���#�&"Ę�S\��)�/���r}�5�_�ᱳԯ�R�'��C���u<��铈(~�z"ԁP��Ŧ�6�����yCiN�c�e���&.EU�g����:�f\�����m�C�)׌�L�_I\'�l��eE�-Q/z���Z�A7�D:�����	�3�G��n"�+I������>D��8ճ��܇�k�.Z�S������'����)i�����eЈ~��.6��˄�5Em?�v��(���6��ʍ��d٠��A��M:�	C��	ad��X���p:��|�*���Ql���6OTU�P��f�J�zn�#�Dݯ@�J��k����g=ş���Q �����^����d����6ŨG��ZbWV��ۊ�É��ȧ����IMܫV�-�!x�5��r1�ȥvC���5�h4.�8���{�)m�#��q���7+L>����h��و����j�b�����㸀kT�*,jW�����9�WWσ��[<� �_�^���y"�b�P*�ox/a�ʆ�adk���f����qϰX��Fu� ��xH�;���Tz��z��@�L"��h�za��'�R�ّ<���� �?p"�kkl'�w�Nr�w,���j�����w�C�W�j���wH>�s���p6�:uT�ʯ�7��$z�ϥ�uE�W���	�G30�6������Y׭�JBH3�G�i![u";��?Pꌐd#)	1��&2�|�W��mfrz�g4�����/|�(�ě8�4��G��>�	��5�`�T���a��'8%hイ'��-)�FP��Q���{7խ�gy O�W�� �g�ױ*,foWCr��6�1����[hµ��h4sŎ2�1���R��}d���~�^ނD��ɏX��(`Ք/�:��t��,惯R@K�����T/��{u�j;�"��.�(�+�{@����~VUE�Txh_��~~A��C�*_S���&Y8),~rYNez���Ѳ�]���>`�I-��.��"g�
<�=k~��f��	 �����:�+F�@�FY�Z+� �f��Z��>a�S�����!AL���4V3�:&�@��Y<9�<�T R���oA� w��ՙL�r���&)S|�&���ʽX$��=�g�3Y?v!%�7dQ�"xu�ٻ+b�.���Qy74��;����+;��tW�և����c�,ٞ���>�K�-)�DP�6+V?!6��wWҥ�����|9�o֕���@ᘨ;n�F9r�)�&|�$*t7�E�v�^�ʅu]釩T��;S�t>fT��O��]� m�F i��,��UW��ԾE�eJC�!�8s��[�L�3��#��5U�G-�޽[�/��\E�&2~̱�"B_κ��Y�28�_q\��@z�n�b:)@�ٖ�e�r�!�5��Խ�$�g��R}d�3�2?=����0��Y�#�2n ��� [3�
|����kp���=������F�C�}a+kD�;9K�9� ����>}���kLy�9w��۪�1''�Ѕ��ͮ�����IG0E��[�s�h��_O���cUs�k��{;�Bn^Ǉ0�\9T~r|�'���v@�{$�muz�Z�I��^'�C��ZJ&�`y~��]�=��)�0o�g����j��X/�a>.$Ji��f-[qWu�ȕ�q�c�6n�-vB,�����)=��@1�,9b][ㅣ�R�rS��c�٣�XQ$��c�����ݿF\m>�K���S��!ғ�i`w�pf���\�����j�v�V�r�x`&�F,��pһk�g�+:�Ah��Sw��T��&�O���M�Ie�y�ߠ�#S���y��Z3�Rm<��C�5�k�g>����z]�m��*�I	E���"k�<�w���c5����L�$>����?�f����^��y�4l�bKv�3��]f�'�
�'��7l���_�����c�$��5
/�ڞ�����u{�v���,��Ǒ}��b��BO��)�!��!����(9a�=��Q��^ݪk{���]V �~Fl��d7��O�����[�6K��棶�S��\V{R�ZF{����eq�*Y:��2W��_�"�K��D�Iws��4RJl#r�R�����q�[��ϙ����u)� k�NwN|�1.3:�����|KP
Z���v���0F[�M�[9�Px�{���H��<���y^�O㞤���vМ����U:J�iKɂ�,���"ju��^�����4!͜�Y9ø��{{�!ڕ4�Gq�e�橖�,I�W���&��y�����^:	;F�|����*ǲ�IS�Ը�`�Q��wHN[��`3��/��1�{�k୪����N�N�ui� O��5����G��i�Ԑ�#�g핗P$Ǵ',��0�8�^��F1.��r�9K��jr���Oв�z�����}<t!�Y2
�.I�Ű^� �L-�-��[��\4k�sGc ��!�U=�m�9F�����HЛ�L<@�B=��W���x��[�h���."r��cJ<f��ǽ���ug"�R��̂��Y�ё��ڭK��t��_7�&�t��F
)kRU�n���J�R+W��s��&n%qDV�b���'��!Ђ�.�ެ�*:�AI��s��.����@��ė��d��N�XMP�*��p����t���̌90���Ԣ5 �K�0��N���$�K��,�KO`�5��
Z���# ��)�1�[��LL�T� a�9� �h�3_׍g-�%��`�"@��J����İ���K�k�؞R;����ÒQ2L#���*	7��'��˭#0*h�~����{(��Q�/!₵�+��zoF^	$��Đ��͕|�)�Ǒ��q3i��L�_6�Nu��=s�8S��  �7t�b�������d"�	g�Z֝���3���i˅��y�\g��B�x��y=^L�Ѩ�F#曈�l� 7>����6���~p��rJ�J�=�گ���	գq��$��w��do8���E&�4&D�$f��Muԁ�~�f.��Zw&��C�{cx�=�ʗM�1����� |�E�#X0�!�;Y��:'���C!�)��^��}dpk������ �HoFP���|[9�U�Z�����Ǻ����gu�����E�B�M��!�g�T���Z�٦c�%����(�W���1a0�
AQ�Đ!|�-���S�{�b�RA��X�U;���k��� 2�zVo�$�a�����z�[?f+!N=�+�l*M���J� &2�w#�5m�&��F1�qB⇔\�r��{���@ԩ/�p�Z�D�u�",�N���QxNx�+�������h}d�܍8D�E����t�!�{R��ȳ�"G�~����%���F�q�qmZ�Q[�I˅խ��k��nX��YS|H���c���[�F��|�"%+F���Āa��2�3a�*i�y>J��n���^��!��-�er���Kč�'��7�H���;�U(��+���m�叒xIk;F�ٻ�OQ��l������K	��!�y�Aḯr�b��O�6��+��z�Ԡp�+n��h��k��[��T�V_������rH'�(!qU:~nI>�x7�%n��+f5���Z3p0G@b��@QG�bJ�`��?��&�_��09X,nu�L;EY"6[��UHh2��~5^�;�L�Lz�u��n!>�Q�o��'##v�ҵ 3b-h�})����2�CH��u/�(��/ĠWE�?RaZOl�N�����FJc�ʘ���;��B�C�N���ZƸ��(F������@�|�0�ho�9N�z�-�vhw$$�Nઠ��%I��{�dx��t졸�U�,v�D:ս�����)O�3gD��)�r��n[�)Lo-߁�� ���>l)[O(oNx�L��;����s@�����̰�ݓO���� �5��l�p҇]݁v~Voܭ�-�@|b��k��#���捡M�v-wgˇ�E�Y����lJ�� X8\0��G����w�m�X���S~�ﺙ䴾��O�ɌO�6��3U~}_��^q��B���HZ����ҟՈ�f��b�J��/���1�zO��噔��Ih@*ߠ̫�:B�	�f��H�̙D��64��E����n���"�`+ƸL��ժH�h�&�~���\�8�*7#�7���FªF�3�L�9W�m���+� �76�&��_�A�N�*[���J�ˑŵ�ջ�ɯAÃE�.�½?4?]�!]ԡ����:�
00���+A�{�ʧ�庺޺���#��`�z��o������<�31$ަ��/X���y=��A�������Z�M����X@n3ZX�@̫}��O+�)���~da?��d��V$B��GY���1SL�}<�r����k�u��)�D7�E�5RW� �-1�G-V�2�YV~�w�[h4�C�X#(_7Y�Z��c���-Fzx{�S�������ZCh��؆'���V=Ҙ�R�A���q��jw"Đ����*�gO�(�*�q�&Q{��*|O�W-�wO!��Ӵ�O�f	���O<��)芵 �c��r^ׂǠ0��S��/ˤ?tbXQ�_a�\ŗi��0��HN�Bw3�/��=���oI�Y� N>圭lS�y:���� c��3�ɒ��0���%��owb����O�m�;h�JB�����������LG'T�Gn�M�����*?��W%�P������n���]�i���KghW��yh���Ѵ�q^��}�(���dL�;�ǕNņ��A�wGG�GIH�ّu��h# }�\�ֵ���?�TT�JM;LX%86����VG����m&i��\��ۮW��t-��\P��g<A$U8I�ѡ n1k~샫��V�s�H?���j	���_-H��K��p�v��3�����Ex��?:��%�����Q�3��қ�TcJ9����閃�'����;��_�|�&�y�)����N��g?fjÉAVۂ�A�&�q��?t�e�!�a�;\S� �E=D":R�C���>�5'x�6ن&���QQjG���/����H5: �/��]E�CÈ����p Ö i��c��}{�1��5	�V_�3gEp�γQ�c�4��� �v]�6Z%�=���N���@{���7:
���a��������ߙԧ�����eN9O�H�W�q弨������|��'��;�T;�!5�ϡFJ	��"N!�R�T:#r_�|�&B�1z?P���9VhS\��E�����э߅�$�8��J�x��C�q��c����O<?eoF�`���L�|4�>��
8�+�P�b�-G��z��E4ӣQ �6���#j�/��c@5�`Iy�����0�Eɝz��E:!]��]T4|��Lip�;�s�G���(9��b���A3��J��"]�֋{˴L@��Ox_:|�+�e�R�9���?����#u��Z=�w$Ju��"�,�������=�E0��G��$�9��ZZ���O��n�9������	v���z #��8,���!��P6ׯ��.�>����k�}�|�%��yf�SH�짰I��B� ����0���Jv����VA��$u�W�p���۵�c��^13����1l4ubr�f��:���Ư"(�/e�By8��~�"�<o�{���4�����8��P���>{�Jy3TMf�Ԧ Ymֈɀxhk���d�<���.3_j��_��y1�Ҝդ}L�z��N>��7�~����m�Z��dfeb�>�s���ߤ���PD�T
&1���k���2:�W�B2T��)QL�b����)�lp���P*�[(���{� #[��B�h��c��"9Ɛb�n�����B�ޘy:��s��΋��"$z������ms�+�����J��Fw�p4�6��$e��x�t} �����K�USaTh�S	o|�@��5ǿ8�v��b�3�7��w�C���`�C�"+�L֞3���c�����M�.rw�7zwت��*W��ŀ/��������U��`��~��z_�>T�	�x�2����'��Tg�/QT��y$��$q��d_��|�x��G:���6�O0{���NP>�p�'W5W���۲ǚS�3T���+��1�����){�vng��88���j���u1r� B�Sr&��Js�<�Ge��2�_(��`:d���a�^W3�(��M�Jg�B5>����F��C�^M����|�E1G����r1B�i�n8�mD�����:��ԝ��x���epB��{�A��e١D����>n�^�eS����c�l捔����ɰꀜ��EAĂ6r��:���>�/��Z��h{��r.�k�pF��C6���S�v�yM��	Ga��5�s�l�Oӝk� >PI��zy5�^��!���+w���f��=7�V�5td*�T/Qs��sh�7l��eq^��d��t���殷Ú�����^�iR��5A�r�
���1�`�u��LrH�A���ʶ�=1]1%;4�po�p���@ܭj����a���e<�̕&W~˓ ��c�q�֕�[�l��a��M����ܛ����O'+!.��Frm1�4E����"�F�	�x��`Ե�k��׮�Y�Cd �$. ^B �r�>�O0��&�NK�⊰*�p�1�У9Φ䬅�����)�(�C1��-<񇌉��I,��K����HB�.���[ 2�O`�Y�_{��9/�s��"H�7m�h���w}[t��ݞ2��4�uL�6�<���U����xig���udΟA̩sj�g5eM��G���C8M}��B���<��sd�ӟl�]
�R�����}���p9q���9��b��xV�� �*�������<�R�w����<���b�ڹ�"[#M�Te��KNףּ�W��\�:�`��Z鱋e;ЏkSWy�9,R^���pO
��k�L1��~źH9�:�|��O��SB�'�c�D�.���s�^!��\Y�4YW9�sUrR���h�.,wg�ϖ���'�o�Ě�Ag���F�~��0�/h�٭ל�U��Z�m�~w�7wA��_�Һ���j�)Tj�8�����f�t�����L�r�S�)�q�inDGŉv�Q�H�u���O�r:F�P��-3|3�[J����cI�{^ӝ�}>������-R�b��s��.�H����X���GI���ǟF0�-��k��Vj�Nt��U�ت~�RC��J������e(Zb1S��#)5P�.�1��i{<������ݣ��@�ۣ��-�L}9C%���!�H�I	1}���j~�A7i��6���"K
��v��пA�����@4ӭg�w�E��ז�ӕ�2�����i:�m`��{���=���Hu��ϿV�+K�R�&���	�Z�Tv�Ls��	;@e���<
B�-�3jF�ZR p_��&w�v�ٹ�4�ԗ�z*c.:�|�P(a�T�a���91ڷD�����1Wa�S9��r!��c�E������ƖǞ�t!^���+�iU>��p]�^릦���֑6�h�A�ѫw��F���>Π�c��	���`&1��NX�2fb�LY6�ǼЄ�r}�k�Ob��X<��S֔2g���lT�׏��^��)4[�c���:O���C;Yo����q�U��\�Û\$�x�V���#�(�*�,�B�]\:��m�aL8�+m�i̢�����1Rܣ���_ڄ<�1!�M��}o/2�\z1��"t�م��C�Ò��~����lwj�UA�O��N�fFh�*��>�^������Aӂ.@Q�-(��ZWC��<z|=A�t{�UMX>>�����!�J�x��"oT\�:�k���#�����^�00��V�b�",߳�Ӳg����\��1K�������+𐻒쵀>�qt�ʾ0?Z���x(�ms�g�G�Mhq��g.C9=.#ΜL�M$ƿ��*4��]z�5�/�LA��[��j����,{��w�X�o�(*Q��;��>U��7(�3�z��f�N�j��������oТ�ʚFw�2n�N
�;�� �`|�������cd���+��H�:�f�7�������T	���&��&�v��}BwVmo��v�$����ϫ���WQ�M�s͗��\3r�l��!�T@�3]�?�:W���v(��t�]�#�\5��m�BUG�YAvc�X���[)�MzwzN`��5n(/ͨ�Fg����+�$�=��鏄jt��Ջ�n3R��^h�,5�{���z����}��{�5aG��P�O4�
�G�d�T���k�4k�d��~t]��1 �ţ%��$�YA�Ո���e��6 ��������@n{\�4V���0�.#I��*J>1�oIdLV)�'�_߇�Z��*��?9�tQ����� /���3�*����L�9��6Rv����GL�:+{y�?M1����P�e�]Ї��J�N�I&ח �<j���\�as��qE��;�u;��V�&��c?e<b�Zϣ]�W��`�~	�n������O $�����3(�=�[ �U��y[{SJ�ךp�I�k9h$���T?������H�t3S>�:K��E�I��;��J�I]���.ԥ��<�&�.�Ht5r�W�@WM�����2�
-��A穭j�K~ ���
ֺ�N ��
�ְ}��*ŋ�|H�~�#���L���y�����7Ƣn�8\-����V��m�΃s(�}C��k�w���TY�=���]�~�8����	O��@�w�Z@w��Al���O�N�<}d�ZB���%G�s�$|�	�x7V||��再θ4�c�[j�;�rt���#?��9��v��^��Z��_�u����A�r�ǐVhZ'���1��^�"~'�S�3%���g��Ttt�x�Dj�u-��~��d�/Wt��)ޚK	�+9��u�%6�/�E	�Ky}�L���i�{8��(�?�X�C����$l܉��nW��?Rf�V��%���TA��lM;5Y�PE�Q8D��ʦ��h΄.�=�L4nTiο�	�(Un
����|' _9خ�&2�-�;2f�e/�M�e2k��-��l0�Q����9�oo1MaP���Z�v���I/�wh��	�*��]��W_M颫����g�m�z��!�37�@�����|������U��t�:6E�0�p����a�s�c��{p����^��:�s��qIs���;��E&ǌ�r�B�}B&��a�l#�����w~	 't^�9.b�~BF�Xl�	`m�i�ϟy�o��9�O�����a.l��$l�/�7��e+�Wl�t#a3 ��^vya�
�q��/��������5w��NՉ*���+ç�J;ݘ�~΃3��CK��-�U|�!���%��i1�F#,��.Y鎼 �^��@���!b%����`�m��8��R��Ϝ�u��~���J<]��p�ɒT�.qk0�ʨ��#�;zz�����C���u��~V���ݾ�0�.��L�2$I�{�N������#U��"�_ƻq42hOx�`��}r�S����g�%3�o��o����d�)�}�I���!Wϸ�ӈ�[�'"}r��!�oGGɫ��o�p@�z�쐋�-"�"�.�l���4F֘���cd]��f�����������$�� �k�Jל�ӴJ
�;�b�;��<-ۢQ}W�|��p�O/��f��NB���׍'i���`N/�X�X���(@��?�禯�%�ߗ�O�,Q�����x�`4�R���p���N����.���!��\~���(Q;L�M���{��)!�,&d��kc(�]6�(��w?�΍p��qS��S
q�P�%W�O��ѹ�������UÊ)<����C=��⡣Ҥjc�҆Dl� �����]2t��Q�{DB��w��}_M�t=�a��!�a�EZ��7�����@�Ùo����+aH]j-�MM�
����lj蝷i<<�]������Vbx˭��m��-X�b��r� 0�C�p��������a�{�;����՚�g��y�L�8ί;��1�炷��S��.Z��h��>�Z��3N����	�3`Y39p��qH�F�	޸hm��㜦��UF��`���3⧈�뤹�n�)�&��9�{I4����6���I��a���_H��/.��<��r��&oq1���W�����99D�c���
Q�a���9�w����~&!���~�l'9�-�ape�T^��I�Є+�w!�x�vS#�|ij�?��~���4W3en��w��Ȋ�6�:�@�T�"��x4����`�
�"����pC����������+�
��B�i�3QA���t��-2c��:�1��Q���1�$����PV,(7���J#�(8��wAk+3�[�T�N��)=��Y0p~_��na7����Ǟ�7Ђ2���!
��+�Y%��{yp�ä�h5Mh��@�v�l�t�p2��P�R仝t�`-6ˢ�6p����,�����w����,²�ǈ{�	���E{���DI<�g��(KJ$#}��ݹ�� ��m�A���V$"�L�@���;d��_�������Q��Ai�L��@�<K*�����`'*Ir����R�W'w����)��$.|�U+����:�1��@��%�Đa�H��7��<.����$�C�'���_; ׿��ĸ�؆��X����&�H/����^(��'��!���֙5;P�aE���lr;T�U��_2�����D�V�YGC�V���0
4�2rn���An[f�jB!��Ӣ�f�-�T�,�Kc�
b%�w��b����߇��C�UK�iA��(��d&�t�X��c��W��..:����5S��.0��؛�|�)%T��l���O�E�6��	��������xWn��#)�`r��E�P��������Y�����&R@,�7ˢ�4D�k�/�T����RXЃ���u��7��p��w��ezZ�L��BD�qVQ�l1����7��9�Ms�يkeQ�0�Q���Ѐ[�:�%��+�Mb{a�9D�$�9N7X3I����N���}e`?�u-sj�L�i�ۃ}'���<0<e�I�$�U�'%'�|�F���(�c�Lz������gI��
{�"3���-�0	�mX�.����.a��鹱G_\��A �(�Th1��(KuTM��5��vv�lj�{���uI����x�T���u7s�r�#�W�N�9�VI���S8m�ow��d�L��J��}�K� "U$Z�Ȯ!</w�)·@Y=d��ͫ@���y�A�l�稹�� �9%���s�5VD��XD=�����7�u������jҟ��M��ʹv'��F�(U}w���'�BvW��ȧ7Ӊ��v�����2��������c�����<��{'a�,��� �F�`�E TI<�md��nvy�qA���dR<�N�A�<)x��J �C'���^ ���ZNR(d1u�Z^�X�N<V:[0�V��4�L��x��	x���ÌG������w����F]�f����#�(i�,�#��o-��	v���7 ���(�,c�~�ꮌ7���o������X_������t2�|N/{y���8<mX���n�J>;9�u�2p�}�e9�`�r�1}�"�j��]��(�G�V�U+�ֈ��8h���?��B�r�!����i��A$��y��ͧ��Q���R�K�+��6
�9qZ:���i��%jp��=տK�,7n�8��y��	6��hR ��K@�v-P�ٺn�o`���Q�+��3!k��C�Tx4�w �M�����j�]�5�)���Gx���\
��2�� �l�ψ|��I<�<�jƲT�|L��<!�z'�=ԃ���nK�c���9y�k}{Rk
j��ߩ�m>�)���i#j+g_bj��#���O��(,��^4�rVYT�˜�c�����Y'A���vv<,�����*�V/@J�ɂ�*T�>�(/Lw�5$�&l���K� ��%�S���W�Y��X��zK�+���IO�ʍ�oo�@ءv�I�%�~
�k]�h���~pC
A<KW�l����(��6�E/��LP��a�뎧7&���i5��S����G�[��np��<��6"�H���D-��Q��.M�$�#6\8�8j��K��zo����́rb����B5�G���B����V/H�~��p�-3;U���ʎv�i O��@r��
�X1v��.�E&�=.���p܌�WUt�EE�=����42)s��x(�Q�?վ�b�9�3��� ���ʆ@�K�լC�-���UWc��þ� �����q�� `���AAi�uYm�ͤ^��L��٠~�f*������!�c�� ���1��܆�t���T�u��4�[�o��-��	�v>�����׵����RJR�͞>E�h3��Q����+�(�cO�|�$��%k뇑��y�9rN�OZц��z���MGW�ҥj�Rc_(A/�)�U~��*�娺C�/�
qc%��_e<��I��m`.��s]�sS����H�cB���.C7�Z�-a(�j���kEy��7��#e#���L�������4-��'=��Q�Ze#, I�QG�����q�����R˸���K��Gk__z��ș�xHЃ�iO�h�6����۪�����r�w��w��`=�+He2ԛt���I�q׷��Ę�ZQ�"Ce�y�+!:?:.��l�z>ybF����/���P��%���f9;��!stpX>�SOl&.7QH�~e�$���Eńe\ap3��lx�|i�;�i��G�4�S)��WJ���{�ì��݉��XZ���2l��ͷ�?b�>���9Z2!t�㬊��5h)ރ�K)4�ܪ����Z�+`��/%w� �f/�۟�T��ո��Xi��<�t�/�_��A�c�<�ࠃ�k�]S�� ��Ʒ	bf��na�Y����qӽ��)�0�M�t����S.��n����n%)^�L�e��z�Bx��s�S)��'@uc{�����Y��4N�VC���F��C~-dm��Gg7�8����o{���+0�<A1�� �W�[T*�TW�O[�$��;[n9�-C�i��\@-O�-])�W��vL�N�q�.wgN1h|N��"��	��+g��WisYb:�O�~de cv� �\ Gic�����xh�nP�e|GC�0y]r�I�Ѷ��qg���P�j����X��:�B��d' u��9b���bڊG�mm���_bF!��F�j�R��t�;Q�#q��N|�|�< `]���A�x���.L�sҥ/K)���~��%k�tȎM\�ȫ�a&86¤�����!�H=⿙��sS����X���S�F���`�eӏ�ꁻ�'��/���@�եΨ<s�i9���M]Z3�ki�W�$���	�w�qcר��Ӭ��o�c�2O�5Q����)^����hw�<cA��Z��kR�D�HRF��y��՟3�oi��8q�9������;P)M�\�!�vH�XSo,	ԑ�X����nm�+j�c�:z��������� izłENX��p/%#��`-��ST�I���x-��̅Cux��2�ϔ�߭(�t�ve�ՄI����&�P��� ��D\�a���ˇ>��*���#w���~���C����@��;bV ���f�L>>�p�Q�EU�m��A|!�Em��ݏ)#b��6�Q�/�S��@�r�B��Z9��9AR����K���0e
�`�4�u޾g��Ot��4>H��zE6iيNI�W�����>�P��7����#���`��W�+����Ik*�b%�X�3��y>'������4�n�� �"%�S��R?��"� ^n��%�� �!����
ʿ�����-�$��6�>,�^�Y0���(6>b奦��!P���ln#��V;�B"�w
��	P��9"gj=�����F]p%����9�y�={ƴr��r�5خ�n^+�� <����U�X>Ӈ|q�.!�3�����TT�!ذ1Bdn�i��
S��9T8��}{�j#%���n��N��VKfJL�a��A8��<9)��IK�^�,JQ�7 ��d�h�I[�Ϫ�R���6.E>��M����ĺ =5T؝��J�:��%O�h(��ے	\9���N��/h@]��1Q���#
_ʭ��+�Κ�Wo�|�]����ɱ�X3��;�	s8Xo�O1s^vsh�Fb��6?�:�_�Yl���˚��m���@���
L.�^R�B��̿l� �1��;<�2!	�h�;�I�� �%=Nzv@-Y��S貱��?���͓aH��_>��gO�Ɍ�����e6&�~'`����|h ���PaR˩٫۫~u���$��W��<�eC^�ƌxOhB	Ƶ�ދ9���3z�(N�|�2�GS��7X�k=�Vx5��\K�����mwޔ&��t�*=�/�'�	v�=�6b����S�|��ާj��51���g�lS��y��9��ǏC��<���viBt�^`TS����`��H�çS����]���q�-*GW�	�G�=��B�Z"�ɖ�=)�:�m#[E9^��w��m�#�+f ������"×"���P�P+ E������#y��m����i�VTxrSe��d����,z��J�:SC�a��uر��k�~n���W�K#p`�y�Ĺ�@I�z��0�˳ݮ]*�f:�5J����=P��ŉ����ßs�BF�M�U�H�1���⅂�-��2�[n@
z�K��F{�N�.��T�kM�'��*���9�O�����p��]Ƨ��S�hfZ�cP ������B|>�D�h�7�%�o��� �r]�W`��*;Whw�k�'=�J@��Q�bbg4��v�~��"����G��b�qL�	��$���,���}�D�өifr,�SY֕7_t��ƌ'|�"��e�����3ql�����d��B�S¦S�":�M7M^��䟰^~t<�D]4<�dtSk�d�"[�N�B���FRz'\��%-� 6Y$�y)6˝mԴ�-��]��k��@�9��')  ��wRX�����j��;��Η.�ӆ�>H�V*����~j�gn���@�Z����������/Ѷ���%s�r�/�2�q-����e�2�g'��T�k��l��K=&<���հ��ZI謀<V�0WQ &�4�5������ ���a��
qǊo�4�uz�B�-��
�k��>�0a"L�������to&����X����x��ph�we��I�g�\������� V1c�֓�cm���{��N?.Fw��=e� �[��}m��S��u1rn*��z 3��&�H�x�Ys&PZ)B�&��m����0��N:ܴ��L�d"ed���iH`a�\Qwe�o��O�#{'��u�RL����v�TT"��tb#<��t���.��I !M�!�k��&ǈ@���ݩga��������;�	�D���4b�g��(y��9�YR�����B����í?�J0�#�%;:%y"6_*��Ē锧�}x��"���~� ��z��$����$/���:�䒷��-�ڣ~�Vɡ'��c���0���C��{�C�p���$i�����G`�f��A35:U���vU�c�.�8*3E�k��{' ˒DgA�7��7yk�#%�"^0�11YCȸ�nmj�Ą�nh�-�\t}�v*�+wӤ1�!6Oˤ̔᳋D�Pl�TQ t�g
�0�N��:�JѶ5����n�"HYL�����񼩵YIJ4�1�A����r�dަ�&���f��ss�g�S�_L6�����r]lE��^�^�7�&��y!���C��&ϤΆo��D{����$*�ߠ�*�v3[�[�KZ��bM1O$�!�T%-O�%�Y��d��%�ԪJ2��l�����)�N��%�]5=���#ե�9M��!��+dc5��0��P�ǁ�W)2��?v}�Z^�V�VKI(�K_&ǀ/�Ϝ�qxF�c0I��?RG��k����f�����5�[�
o�lتv�T�W��Ee;ᯣ����0L��u伨�I2kUai^/y��c�Qp��jO=Kux��O��ki��$�z>%�kY�e�K�{�8}�G� ��)��1q�c_a~g��"����\J�S�$
1�蓍�I�i�k�Ab��2Oi�F>*���SR��� ��9��a^ϝ�E�!�|gy�`6Q/w+���*�p�Tl���:m��
p|�2�=k�q�.^jx���ˑ����.�(Ȁ '��'��y���)=ջ�y'��K��qծ�$���_]]74""��@�L���-��A�W"�i#>����� �QV3e$�K}ȩ:O��Ю���N�TGV�J�ˆ�5��7g��Ŧ�Ա��]���̤V��""n�8��H��j{YĔ���9 ��!uf�>�O�
o����j����1����t�P*9Q��Id���V9�j�,^�=pr�^
e��c��6|ƨ2PO�)��6������p���C���8���W%KQkn|�U@t+)���7&^�!A���H�3q�vU�c��x�Y6m�NZ�ξ(�"s'���Ȉ@
e��W�Jǳb�"��m�r�(Y<u����m�X XX����د`ˢ�e�s�{�.��G 0MZ��J�ˏ����v��h������2)��n?���V�b���l�ƈ�E���G	�k���As#�������j�:jE{I*���#����~gW1ٕ����]X�[��!��9y���\(�<Al��}�$J�tBiW,J�w�q��H��[�)��K����=�,U�u�X���a'�l�K�۬J\-�6/9n(%]�5(��$���,�nh�����-�e8q�
BG�xְΩ]O�Hм�;�v�(��HƦU|�ހ�r8dOMx��W�١1�r/����4�{<*�Yׄ�+�o0��棐t ��F^��!�gk,$�Mh������=�vPC�?�n�iL:��=������`�ZЖh���y��$�I_���s�a���1��R�1v��f'�,(Xz��u��f� ���1�X��s_z���_Rκ��my���)��e�)�!?<�YE}�dj�W�z�E0ڂ̻ZP�Q� 8^
�������e�3�/��5��� ��t����-/��g�C����0����Pܝ7�Si^ab1�62��6w�(���%��x�|�wo�D��[�렁�hBm�Z@d9�"��M߼db#遼����o]>F̼��e-�i�!e���E�z3�ӮJ�G$`AX��c�b��w�/���NI%2�P=H�p�{�����p�1
�6�O���)��Gd��0zNnف-``#oD��i���`�7�.�~?U����.�_��/O�=�sk����,�j7��!l��� ��Ê�[��-�%�A��8ևVId7��	�Z���&x�\8?�wJ�c���7����`�IۇR���c��3b�����"�;�#3LJ+?�
�A�,�PYi����B���2�3^{�=�2�'��p�
���ε7�t���۵��=�Q�K�/L�@��[d�Cy����q��R?=;B���B]A�h)%B�e��8^�MM��c�H��Bq�=��@�1��9��Â$R]��Ev���d$�Nf�,v�g��+�O�&�[7��=f�d�'�+m��'lF��NH����r�~�N��D�\�e��ط�}u�&�w=��Co�m�z��,�)#se�_��O��H�j�%T'�vX���0��na9<i���D��>+L�ի1mW .�+	��P�j� �W�6[y��Oz+N"�6^��C�gX<o�]f'+/��9�l��0��%.�
����"ͩ�X��Y��pZ��:S 7��7�&�UD����"�?��B;�6��7c ��[�Sn4���:�F��%�ZQMk�*:�*��n���X��P�:7m�`UL(0m��#�}Mԙ҆8>y��\���� �-v@�<=Y��̟�Z6�K����JT�����&�@�)�%��C�����;C;o�Y~��s��US���a���2�exj9*��5Aa^y���ws=��R��3_s�( �K_��8_m>` X�)�L@;^u�%��Ռmo97̜�|āG�T%U�����7�86`��t���du�eӁk��P�=624�q�p��+`��2���jYo�&.�n��p���x�R%�@�fo|-
9�q6���<���|�sY�U��"H�x��<��@�0���fG����6����ٸxV�0هl脇�$�'����p�a�q�����,0�A7	9��q��8�$$�5
�'#���A�qZjkWo�WI�0م)^�rׇpSr�����ч���_my��sD�����Nb�5	S��%ս���4�m0.\��[����y(�>���� �M�l;�
�'�Xx�!+�Tt�拒���\iI�A�d��(��'"���j�"�H�&���i��<5Fa���C���PRx�NT{��%b�|M]�2���21c�w<��O����М�v&|o�N��� �/�g@�g�rh��!�U栴��v����Q�P@�#/���gȆ�vVg�ƺ��S���YT��6	�V��s�UfcǠJ�K��4B�
q�LG�Tg ���v8�k�ŏT��g@�f��!�h�$�'�I��'л��V[i��}V>?�n5�(�x,��׷��L?�@+ө�
��,�Tz}#�vUj~��u<3�l�B�3�%�>=�]x~j�5���}دꙶ�
I@Z��%z�6�\�Ë�9]�?}E��lׄ*l�Lp;�iΝ����ǀ2�Ͽ]laB|l^!4�L�Բn��WO�n��Ol �\)�@���4�3͢�?��3�"����'�ǝz#S�&�=ݿ�6���6�l	K�9�9l�{�Q.nB�D���1ȿ)~�*��G�o*����Q�����7~��V���bc����0�/!�����)��L���#VA&M��@��[��:�^�.D���j Sѕ���W/��e�P��̕��9-\��aQ�:�.��N��$u�F��7�Y�ȕ�t�"G:}ƣ!�6������,h��f�)�`ct�-��@�(��\ْ��f��_d«@qҕY�[�=��e�a�"��סfݼdJ�őI<n��ϕ���<�cŌ�c���A���1�`�w���7y$��3�]t��A��=�<�"I,}f��'$M/ �E=4��RgStO�.�_���q_�K��.�M�/ǔs��j&��h�c�� qW{/P�����u��v"���?���{�L�L=ݻ�2}�p��,�����7~���Q��s�
a9�@nKa�H���r]?��1cz��7�Y7�B�o�;f0B��`�`���i��i��P0P
������CbX��(��P���\�Ҵ���^��*�bɋ�+�ȉ�ك��G��
�����ouw}t�-#���`�sd_<\�&l�n|�SF-"�W*�f�"�H�K����a9���š��[�<��|�Ó;���I��he��Oآ��9�G��SUL�}�_u�/HWAii��lfmoA/\�3�r���(�u�TS�
_����9^_�a�^Gn2� �	�K9�JN%���q��蹕.o>cU�L��Ӏ�4�O���O�d�Ѡ��Xع�\�j���6z e���3�aA�lW�Cf�v!�y'��N��Z"�]RcE���R��ÆQ�m�����4��)�0��ƚUe�����de&��&�q��_��n�w�O[��,o���7p��
<y�O�
��-��Y�t�M�5��.G��p��F�cӳ�*�}�M��H���'2h���+�o����9�U�2�I@顗r���J��f����[�9oS�=�\!�^�3h�>e��.e��?�[�P^rğz�0�Ʋk$)b�VA�6E��)qָ�Q�����ă��óꏰ�B. ���m��(	e)D�I3�k�U��l!H�	~_[��yN�D2��҄��?�^��˪�Ә��[#yP8��nA�l);�C��
����	ywO�s���Jڒ$�4l#���(��y����|+YN3��"������.L1��2d�����͈^o�x��ǰ*Ҡ}�O�ጫt-G�a*1O��J���ƙ��(�L��S}�������!���m	-��C��\f�]��g�5)0q� ��e�3�J4G�ϕ[M��N�Y���?�G�O�O���4�59�9yMJ3C��}v��)�.��.P�k��i�s�>.
ύ@�.�:�&� \����%%[D.F���B��]���i��m"[�겨�t^�8 #X��{��*�F���RHZ��Ƒt�p���* >R�`�R��;��
4m���	8��^�G��@�rS�%��."Vs�mƯ�N��aK�?�e��#�H�UL"����eKo)9�Q��c�l.��wE��=�K��I��
+���9
ӵϒ����]������k9���E<�`xi��F �27WO~���B��b�e�<*��x��>]M�z?��vb���i���1p�"7W��jl~|�Ɖ���L�!��P֔X�,L'krB��-�@=�������I��l�%/W����144=)�>���D4�S<��.�$�]��S�gF�?�ċ��S/�T|�5��.	�{b�{��TMhTι4��T�M����ɸ��q^��}l5�.�Q#؎�7�Lq�C*��2��1xft<'Z���i9���Fwk��<e��xN�#���������F��ܻA����D%�L�b����9��
���N
�W��O�S��XϧqaĂ���w,��Rh�(Z������	���}�u�m0Jr��]��W����$����xb/��)�Ϡ�W)��ӈ�*���U�Ek��<H�d�~�l��Z����!,1��m�:�@JZ�����-*V���c��_���4y�r�������M �R /}��؄�U;KT�a�$�2��0Si- ��τ�Xv��
3v����Q����d��J�oY������︹�A�Lmq�-mpV��.��{�(�3�{�����A1G��k� �|��bO�x�����`���Y��.M��;�{�W�A�1=����.�W�A�'����Z�,�]�Q�'�٥UȀ乥��ҧu�0fK-�J��A��qnAn�4̃G)�����M]H�$�|�x U��=H� !ܽ��7#mʺM�?x�q��a��{�}*��h*?��|.��W�x�ͅg�r'�ř�����˾��[8�|���*���G�;������rq[���n�o�B��/1��9��]t�Ja-��o��� �P��m���t͔Cc�O��_�an�|AuC{����W�n�]�툜�~	�QQ:S=1���Ѕ1�ƅ������F�%��YK��$-Y���.�<У�w|\'ʭ}���Q��N���'��A�)���B(%�*��1:��Orݰ5��i��׭��r9�x��1�{$�/��L��yZ�j�>��3�I�z?��
�O�A{��QQ
 9Nݦ5�I��)z��:���(�f�(���f'o��J�~dP��Tʓ��j���������):3����Y��:�G���zdu����Le����I�a��ޏ����km�it%Ց;�8 /�N�t����GD ��:A@ ȭMݼ	�G���iV!�/V�y�8�o�x�������FNl#yt���=����"���u�S�y0.�f3�� �Un^+mܗ�#�L�qL��u-ow��-_���t2<D�,ݲ����B���Y�J��`(y�y$|
�(/���2���ex�{܍1�`�q�Y�k�'��io���&��~xj�eKa�n�E�h��ݹ�[?iz��w��U��\х#�
vA� ��%|��g}ꪠ�@��J�xMr��J���n�M\����#� 0���F�>{έ��6E�B=�l@�8l.g��� ��g��}�	�r?���b��Cx�9���8��QB�&���h��O��.���L{�=n�U������SG�Ǥ��t�y���@+{�؂壦���y��8�ɢ��K�rg:�gS4=�V<�9i�
~#4d;�fV�V\��H�Y��bĞ�ɸ���,ml�����cm�N�΁��m�|��,�Z�l#f��$�O���ϙ�2�E~��*l�<��e
w5�g�=�����M`sTl�>�Kۖ�[穟��9e��{H�^\�ϑ�#?������9Ux�̜�
|�^ˮ9��OX"x��\-���~��I#]���7~�в�=�w�&���Ӣ�ۻ�3��m|)�
�|
|l��6*O����l��2��7h�h^׊#o�q�Ӄ�;�I��/렃(�$��ٓ�����*�������#�cK��P]�/�̔l��i�eȽ=����f�N�j�svū�M�55c� _2b���e���Seb��}���\fQ��I�K�L�M��ʓS��~1��+�}8��>(��䒴J�Mś�5KA�UD�. �˩Y(%M��oP�����\私��.��b�	��o3�:���)^R���}:\3Q��Ψ�!��V�%D<����ga� I,�Cލ�A�AO-ձ�|s`!SA�WZ'yv��G�޵-�5�6'�ɛ�qBDuJ��q���lJm�DmT	?�y�GlNg?�/�h�z��v�K��~k��z��g{˳]�G	L��ҟ���3�b懣,HG�#���O�U�|��-M��L�n�\`l{�W�7�Ȓ'�*�e���~0�����ؼ������#@�������Ϋ�������C���Z%�JjpCnQ�ʾLB���L�؉�q ��I��[d�#�c���Q�)/�f��K{u��I���I/Kq��cj�<�+���R�_�����a"C����G��v���Hz|�)�.�����y�T-ri���uU*0�U�s�vt���CSԸ)cS�k���u%����5m�%9t9��13�wp�a����.��\g���s�KY@e��H*���/Ro2��{i����)A��n�I���-ɼ��{k�@�N�C0V6�y]��O��W�?�ϴI;|s�ibS�m/+0;E���x#�q�N݊׌�veԲ���������`�3*��&N[����jz2٧�f"v9��Z�t����YU��^?9�����GT�`��J2yV��3Ӱ[`s���!�aAL4��8sL��c+)���j����c�3��##诰�!�>����t��1����ܬ�*�E ])��qr&� J���|��ckNS�#ՒA4���p������>��/��ThV�b��x��r�9���%(|��yY���Gy��h�a�|�N�����݃�_�m)�� ��	����"��P�'\:��t`�p�b;bКe���X�$��;D  :�[q�E�[�D
L*������E\��ʸ|�S6d�M/�Y��F;O�`���}�N�4�{#}h�����_,���+w Ow�~��?К4.��<�wl6��e�Rx-���"�!|b��O�F'O���ł��R-S/�s�vH,4U��Lz�k�OQ9�*�7*�M5��2�v��DɈ��s��=�<�
5��~V��8�t�:L�f�M�K��D��F_�D�/{1�&�7-�pHuID���ҋ��"��PQi���kSu��0����U�G��K0[Q����ڷ�>].e�i�T��}����[6'Ϲ`hh����C@�1����v9آ�^˴}�L:��!菭s� �����x	���۬Vx�qB�&Xi�+��8#|�H�0D�g������\Eِ�h>�G�Z��UZ�͠��� %P�q�:	X�,P�%�N�X���C
Uͺ�l���K��BuP�4��ܷ��DTF44A���:�߅6��>0\��9]��.n��W����!�\�җ{�N����N{V�,u� ��(䒾���p���c�M&f�|%�����Srױ �A�c��
p���g�(l��;~c�N�r$��E���b)��T#��%������U���o�e��`<T\�����$����'��A�j.B~q�����j�61�꒍������E�x�C�:�i5�}bcK F�.FV_vc��]f'�3�v�L4뽏m��K�F���̪��C��o@�Wy����W�"9Q�FȨbF��Yaޖz}��G>�bq&9��a��fj> �%0�H��]d࿔a�{t���f8����]�	��ݖ�DZ��?*�*.R�b�cU��Ãb���b��$V��Ÿ9<w�eR��cV�
���k�iD��$�[�0�(UPY3L9@#J����A���x�$k�M�0M/s2�0����E��_�$yҜ$��mmb��F�Y:B��:B|.��ŏ'�����Kj�����̺��Ǯ�kiZ}z%v�WMm&8r;<ȫ�����B]0��F�%��ο�����*�,�5���X[�t���n�.�"<^�Z��z�$��i:�A=үS/�v���Zi��ɓ��I�����y$�=��B)xf=4�1塻�7�a����!���E�m��B��2��Ut����������Ev����[���,�E�r�Z(:��^�V[))Q���ObsC����W����,�=�v� �!�X��ߖɋ�$=��(�@�E�~=
�C2:ϔþ:��>�B�W��~��	��{ GD�nT�@B�H�=>����ҍT���N�8��W��E$`�9Í�/��P�W��82w��q�П{CP��"���Ѝ_���&a����~?�q�O��tи����a�UJ���E�
���R������Q�)������d�'��2:ezΥ�*�7i5v@��g��9��a�;vfus�5� �*s�A��nW7��������Zr��E��m�U�qL�O�"<^�2��䴺X�͹EF��f�A��$�s�S��>Xlquv��}�.v�	'���B���/X5�e�o��N�� ���f�vj���?`���$)|i��Gk���g�9�'0��s�Zi��gkf!�C��-�Twh���C�xk���A��0i����l������\��9P։^����3�&�%0��1��AN�E�̢8~2���s��v����	��^�I��Z�x')�����#�t,n�_���0��Z�]�V8b#Tƫ��Ɋ�V�e@�vʕm�����B5wq�?�9?�`W.lO�~%�sA>���~ԹΩ�yQ��S���W��I��kE˻Hy�a�)q�v��{���{��>z��G8|�7�	��P��KN���f[_$�hzS��,̚~S���Bȏ��m	�x����;�ep4����m��
��IPi��{�d��{A`J���$-���5/՜{���A!3U�}����]Y�J����@C��>���5r'��"��'s0��.�Z�����i�Ѱ��P�w/��J}�5�c�T�"�nÄl�\��T"����e��R�X�_>�m��k#Ⳟ�p��w@H2�Q�!(��~�xI�FK���W�h� D=6�;1�#�(�����z�R*����T`���Y���%��P��,�0/q�Q��Qg��Gـ&^@���t}�ԣ�Z���W8�_�8V}J�����54�_���20��t�"~�f}�^�ٙ-.m���ӥ���l�4vY�o�le����1�BCS����hy���%�+d+��?����\�"%R�qi�ح�������cx���6���Ӿ[M�ߢ	�2ȶ�./?�m�hY6t����]�4)���#-ϭ�H��[���Tjz��+�I�5]	���ȴ�m'\�2Bq(�̔t�:k|�����fT>��ʦ���	w���j� a�/�0����-���əq.'9��;0K(�qZ ��6�8J��J(7����*��>t5(����� B��U����	�)D	����Cx0�t:š��#$I}y����P�[�ˡ/R��*�P���o��Pj���<�	Z�z�-�¦Z���XO��6����,ø)1]�.�Կ�XK���0��$o3#"$������jNMu�W����:���t�	�y须���T�T(&���>O����j����fJ�Jj�-�� &�^�X{b�C����[\E`���Z�/B���$�)�!se~�8��e��k�#�&j���4���/2�)�m/V5v`k��,LFB<t͡����`5�$�����(FxH	�&L�I�ow>x��J;r��P���	,��@H��A
�jI���U�N�.ue���R�*q#�$n
�t�;q�X��.PӴ��\)RI���<:EāP��z,<��[O٣�w�kbV�X=�e8�WF�u�Hlj?�5	�Y,Vz�-�nC����#��O-^�qm�TQ�fR�b��ZX�ͯ�k��mf�x�9��J��g���A�j������'��E����P���y:МC���� +"��51�&f����1��/����'�����r�w��ȣ��������!9F�~���z�޶YR����b΅�o��2h�NU7	}0�i�c*�/Ʈ!���)`|,�q�\�w�N�\��N��a{�7CO���_|6)"*�[^�P�a�'�Sr��	�n6��b��־'��κU�n9��mc���K�}*�> ���)K��MǢӾ�r�"��x���4ю*@I�U)�'�y���^40�ϧ"m��E@p)bHy�=��U��T���?̈�g��MHv{�6<�=퇱f�۩��p�TR[X�-䌙���H~�?O�F ���� �\t����Ag� F�wO���4M�ZYD�?�lq�-(GperqT�����ڻ�N�K�2_µ���"������v���Gmc��)�o��g���J9���)�i�n*i�d���<��T�l��<�EK$���(���v�A�[��z���sQ�r�S��a璔���h`t��9vY*�����h�,��;/�l�70��2:�pH�b�x� i}�md�������V"i�m$S�Ĕ��"�-.��ȡ`/���h���8TK�t���8�ْ�eT���҉��F�Ǫ��B���7lO>�z���}�5 �h�	w�d~&�y�ǠD�����3�h#Q��P������Z�i�}P�%m�A�0;� N�S�;Ft-�T�gE�H���9<�濴[��{��d�<�,%�/�0�sJү�2�f�Bc�߸P��sC�p�MZ���~�2p2]L�"QXy���	�P��#����S��i�-v楰��k	A�b��S��u����S�%y%#��'�al�n��>�+"i>:m+��[�F36+81Z�.e�Λ���kʺ�i39���z��:��w�n^�ߵ-��(<�2	��1,�L[���4$NL�J�6��iG�D�8��si����6Ҏ��a��7�A�g�_0Z�E0iS7b��dǄ�م��i!|��Ԯ�?��OW:�(vrL �^�`���P�x�E��Y��85/���r��݋y�W��8`[+�"��KMOS��}���H�@h:�x�s��D���0��*��{G��:���{D��H_���V��3�s:�,��Y|��A�SW�5�^���q��W�ߝr�k��6#f�@�ʥ��s�u��ɲ�v����r�[v�>�1r�2�~r�� P߀^U��i0�`.�Nfm��v��jH�p;����B��j���T��j+��ϖ��
��_q��twO3��9�9T��}!�`N 7hЧP5�飱, h���@�� "�0�7z�l5���n,k��o����j���Ռ�G�+��N�o/,�,�:�v�⸭�i���&ڈ��HU�V�]�W��d�GMD�߱�I`܁/�Z��'�n�?`�y�Ƌ�����⻻��E8*v��G��pI7����c�P^1�Dr�T��x� Fw�7Ho,X���Qs�}-�FJ������]���j+�l;�(a0J=$o�F��$����.��!H�e�t��Iq��3�
�:�<��T�/����m�"��b��~�>E��O��5.A
�$�n�L�1��p�Í���2D%(aXf�LԮ�/<�)?��<���#���x��L��Hd�A�d�ix�)�:3�a(8�:�k�	C��)5.��������Qxp�-~_t� �\���p�E{���	�M.��b��Bվ��l-���Ni�y�LIU`ѳ5=V$ʅt�y\#TS����9#�K/�-���_��*ϛ4��J��<��1j���1|�,�RaiT�2٦k�������Y0G�Ḛ7�����4�թxϿ�<��}����Zf��Z?���YF����_��7��U{"P��3��4$���K�"�y�#ݵ�J��px�v$�vzٖ����\R���l�6=E���H|hA��D�W[��%Mж��k�'�5#��*T�2ż4�¤�݇{��Î<.�D�9T�w�*Ds
����`�J���u	�:
��M�����B�mMp��仱�	���_���Y��b��Zh16����Yyo�-��}@�\?����Le�B�����á�"��G�C �l�v�$Fp8��Ȓ��O���w%�����Ocfp�c�2�F�v/���ݤ���.}���5������+����̪���_Ł���뤤5f�"�"�MT�X�L�Cp	;��=��I�qj����[��+�{.g�����y�3�ͳ��8?KV�k�����X��MYѢ�>�UQOf'�ԧ��*x��FC�c4b�_b�)7A�f;��$�C{j����6�Þ�����o\k�ԱNu�96���e[Q
/�78	�^�����t��[ˇ�y����.5�`��_�QW�g�6�n�ү2+6#7�(�H�K�6�8�=���~<�u�Ny��0��+�z��5 �+� ėې��վ`���sZ۔!���P?s	�bΑ�L�(�+��q༛�OX>/O�*ɶ�[���2$ A�����V�t2���h�ׇ����� |��c�\~�~(3�:;��(�*��5����I�%�/<%b �b�3�P���{�=�	[��&Ga��АJj����柱5��t�r�1�8A?��>ܤ~gK�kmYQ�<�LHQ���;@>�FyE�i�i{��UN�2�v�ly�Ŀ7���©"�aёj6��y�#��{;L�8�C?�J��1�.��0(�|mgҽ=�c�y�0���i����%�뱠ds��zJ�/�%G<!p�D�Z�v]�f���v�u�S��]}!��5kEńҲO�CX���<o�P;�3��u�[��4���k<u���o�����Brd�q�%������U�&�S� #���R�`��q� ���"�����hg�&j��̓f���̸RE�C���L�z[�1�]��� �^�C\���tً¡Ӏ�����WIHEy�+��Sޚ�tJ�^8�z=|�(�~�����i!Ԁ5l��0�	J��m(���u/���'4�*�,��S:��ذ0]�@�$�,�;a[�kl%�tܴi��jb�z+����Ό�P?������v�g�t^<�Е�a���:�IJmBs2��DL p�x�U�~B�F��M��2}ڭ�Y�7(�@'E�9� �[bF� ��(x��f�'�Do<��zl�I���U��1�XTUp�E���´��})�A�T�# �����p��`����'x��Z��>��q�.%i~ֳ�x	�nS�襐k�3s�\�:��Y�}/�T����2���) ��m�X�F���_��,���m�N���sT	]�e�j=㒚[���ΜN�q�9�1.P�����=ą���#<-�����n<V����tj�W�[=���Hܩ\Kiy�R� [w@��+�>S���N@�!��?n`<|��"��;2j;���*�A'���7��=̩�ϔ�+�.�bLq�=�A`�u��(�`�JV��*%[�!z_�����l�QA��w���^|#�Cg���<�Q.a���ED:��f�i���E�LQ�����j� \9��SB�p�B<�	��#6 �t%YɡK�pq�e|%WY&JS���u|z��gP.w�D:��
����b6$�e��pkf�6�3�$�f��X�h*��~�ǤZ�:2t�wR���A��B�BI5��26��,�� �i��-}�m��gs����ȼ�y^&�
 F�E��6�����(/�<�43��oGDH"v�`U��uVܠ�����P�ri�+�{̳Gt�)*���\_�P$���
�P�(���S۱\���⁕_�?�4:�A�/�~���¹I��"rDh�.5'γ\ĉ���ކ�"n�Y�-����m�њ7��P�Ƣ�3��H:{,p�e��m�w��� �'�%̄�I*r�\�.���@=����0)Z�#�L+��X��׌�׆���&�|�Q�I��L�cS�_D�B9����6��e��/����Fc�)	�e@�C�S��t�P�h�n(���*馿�~��"4a�D)P�7S�dl&ՙ͇7:MԠ�?��_�ę�#^s��:�.���\�#�
P�`�����Ήh��b�é��i�\����m�$���x%���PT�C�Y1˙giYqb<s�Fi��\<�P��_�o*��8A}�^��Y�$t���Ӣ����l7U\�������h
�}��"Fuڥ���լ�V�dtӜ݁QO�q襱`�7��7�T(LiG(e��YL�
�>�#윈���-d#&�i�5��9p#Ϋ�Km< �$����'�-��ђ���Ĺ��lr��8p�"g�s�����B��y@k����7�X�����]�Z�wtͦn�z>g(��#]���_Ő��b�ᒳ-9j^�>��/�zT��2¥����e/���{��Xb����6ţ�����=�@��AD��5��nbH�x��6�~j�KD)6~�C��@�:��~�*��H�Hw߲0L˘��N�z{��߾�)��R&�@؏�aX���.>M�b����}F�����#X
nk��S �/�.��X���G|��%����XW�QR�%���<��:��K�XE*K�F�it��O/�����v�U�6u�����T����S.�� g�"i8����]3hOr�
t�a�R~�.W��G��+��}Q�/č�)�&/��y�"�紐�:�ps��g���Y�g�]'�������R����G1δ�M}O�Ųi�@��$���K�K�%M�&��l�r�-]�rf��9�%�&tѭ�E"�sRH3��
��~'Cv�9t�T��fEw�s�^=4c��hT��H�Hv���oީC��T��	W^7��6���d��B�ӱIa����Y昀�EWwM�a^N&8CF��=z6D$�Q��)�>�y	���x �ΰ`
lG �-F���\P�ŝ%�u��K�;cQ��o�9mڸmYC�1�,k1�kE�5-1�~�e =&�2V�J:��#���LiN�����ݑvݧ���B�&�D�5f�E��"d.&����0ݪy�GƓ��!������h*��9Nt��P/�C��8?� Om΢�ĕ𙫞ۓ��@�8��<�@�:}D�J��-|ܽ�z�v0�oQ��x] ��֟C�&j97B��"$F*05{p��:W�,� &09�O�-yf���?Kj-�z7��MƷ2��I�:�� ]Zx��o�b9 
x�%n��F��]+]!��I֠<��։t|f9�~�U��)����Ѯ�՗�&/d�
?V���@;�D6q�6��ky��2����J�`���
^S�W�MGP �����Q���7����4��:�6��E�w��b-�������{��̓��K�e�r!0U
w=�9���;���'˰�z?��$�Dh���DuZ|W�tiFc��vK�u�@?�>f��1p��u�ְ�	���p�\�#5��ȉ��;��J�l+"��_��/��!/[K�ɒ�E�6Б���V�ٹl�ɯw��UdSӌ�p��!�c�Qy__!�mx��R9��(�b"� @L��b5}q��"W%0Ct��|M�{�;ܛ(�Z6)g�H��r�֦���_\�S��g�^@���D�`B�0���	�T�=�(�~$%�/></L�@/św�Ro�g[�2v��n���U�S뵑��&�+	��Q�U���>�s�]�$q��)��WƳ�޷OFdx�_��t����Q��T�xج���@?< �W�w�c0l�*��{[�R���,��+���8h:����F�¿�[���u&4����]RG�ު�����/���w�p��<��Ho��"f��/l�K_�<���#�<�ۈ�1��
ֆ��<j	`��U����$D}p�?��3xZ���)��BM�Ga����5��U���4Rf�������x�*��x���0�n��I���QN>�S�^Efc5�w%ĕ��(�m���\D�ePh�zuv�r�����h��I1~;䤳!�h�:�=����'��FXP7?x�����b�R1���(����N&��ѓ_	y��c.yDI���� Nǿ�{(�<�����&�E>7�K2 >/
�L.�+Uj
�����(� ��b�z�3�	�*�4����x\��B��6��4M��JɈD͜��������S��J�Q���(�أ�'&·�	�$,*2�Dq��$�e/�V'i�9�G���y�
>޸q��I��h�x�t%-�$����
�G��{��!��:l�G�WD�K�n�-Q�08�>U�v�R%'�Y��'v��R�h�#w���8���ٌ:(�|O{JK�j�$g�!	~f�Hr%���;Th���KL٤�Sc�t4s ��(Q�hV�	��G"��z��g������::���86�2s|-�n��l2�]Gu_�Q����/�wh2͋J�nƙˉU(j����V� ������`
�N�uՑ�0	68i/D%��<O�,���SIaO1��-G�T�Z $��1� =���&&&��b�k�@@l. a�3_�7{�H{�}�hKVb�g<��3C����2;����֙��`��Y�n�s�-D�ZY��Vmv�@�L�*�Z��꟧$���:�/����uL#��qG
�B��PM��;����>��+_��Cs��Ԣ��ãa�L���ķV�XgֆfT�N�=���ʥ܀۸R���zi^zY�ś#��UqH�NԔ�J2Ub�:td}	�5�&G{��@ ����*�C�i�<��!Te�~l�y��l-Nq	��K�w�:�4b�s��X�-cBCQ��,#d�ľ��x3��^�.��V��E-6�N�Eo�Q����Η��Vfz��a(
{dE�u��7�����ѓ�y!�m"��Qu����ǳ����|��Z�c�v���1�_I�}��Pf��F5�W��¼�Pc�!w*�����v��o[/e M�=9檡��P�i���R3�e�J�v�D�k�N��A�=w�K0�'h����n� �}0�H�rt��呬�<�>~r`�N�P`���s=�������ξ�	�^}/�G�����Re!�+C���V�rU�6W�ps�%���5��t���C	��Qp��ZG�	iX�ղtL��#�P��ez�����SE=e�<�޳���=[��{��f8��>1E�a����Y��ŒJ�H�{Z�0��?|��UEA2�,�5Z��#_��6u2�3��DZbt7��z�	R�z������t~�Tv>v�*�_���iO����AF1d+x�����E�́;�Fk';���i$0��!'v3B-΍�QZ������������Aѽ!]A�7�����3�� �{w
#�YQ컬�ɮ����`��fg�\rY�k�]�+���gn0�Ͳ�q��
�Ut���"�v��\�r�U��	!�9>ɗ4	?�ҭǀ|���P�:C�|8`6�i��\��,�i"�0�č��!�R�����U�S.�Yඪ���-�I�bd�Z�����Ǽ�1	��W�W��Qh"!i(k?49�/O��UkTwh{��Gc3j�w �1���z}]�LUX���[�#�RP�~��z��E�c��`٘Ov��7.�:�S#9u'�T�'�[n5�в��܌B��&�uV���@�� ��BGT8��]ݝ.[��t#$����B4�g7���t�2��1-��|�=�������h ��^�KQM��'�A�����6_
i%�X� �ffl<��n4�* �!��&��Q9bUǑ�ވ�i�S��8i%&�o�G/��B�p��j����ٓ`F~b�y55Ӑ�g=b��ψ)����z��k��`���/r҄k�kSO�������/����{��a�\}D�!L��:z�����^=l��H���g� m�o�pC2Kf���[�bu��+�5�*��� �2_:��WW���!I,�N���2U/���z9J��~��{��G#����-�qa�Mc��hg�{X��P��&^j��<1DT��B]�����\D���9�S�Pr�����'�t�W	��]e�sTeN���]�9�8V�� E���h'�Ѵ34R%DBim�y����-r	>n�"��.Ќ�w����N����6i}��.t	�+?ow�)��~�]F:<�ъQ4�[���LM��a_>��/|V)&,�?�����Z��ԢW�X��5�E�s�7�E%m�"��*J�
�T�̾�^�"ꔬ*Yt�7N,��d}���4�u�1QF���@�&�.���(\Ӥ��D#��D�1b��tЁQD�����yM̜�����M/���>޷��;VR���u~ւ���Iʘz���ϯr���1w�!�&3q���.bI����x��ͤ��j�R̖Y���r�Ta_���&e�D��"�X����#Q��;�9���>�:�(�����j�3\�4x.@��N�9���1�I�@6��ı�N�"r>�O�x�U>�2-c�X*wwx�S�os�'e�d����S���%��*�m����3�����	���'������t��^��ڇZ,���X	�t��R��.����B y �7e}$M[�\���m!F>Ǝ��Iw#�/�B�g�X�����u�������7�Ih��ǖ����Ek�gH�D�Rv�
{;?@��t�2]���)�O��i���������ǌo�^g��irT�0<��,�)��b�U�$�L��H-n�O�ai^�i�|78���':|űh��8�!@?����]�g|T��<ᴮ����y��+��1�d��4A����w[ro˗�̀e��]Ek��C���Yǣ��S�{�����^D�#�nڰ_y����_t5�WC�3�w�ed� �HqbO����J��JK7-�_	��Y�woy1ժ��rB�^�6ք��S��r�@�D�	����W�����
Pˀ���v�j���j��t���Ϗ���L�}u .^�-�hV�p�w��na�d?ј�ɣ�	3��5��R f�,�9$ĀI�WШ!��G�%�GIPg��$,yɵ� .�?|&/H�`����ҵN;W�L`�kE	��1���k`�D�"��n;��!nZ.b7�ms��3�m��Yȭ��fQ�N�}�Nۀ�3�
  K���@�0���ם��I���}쌴Qu�T��ߏ i���I����/Io����s���Y$�!|{�O�`g	����zj4����!p��<HT�U2)���N�Y����&~,�ߗ�^QV�O�Q �ނ��m�8��YU�:�{`~[`E��+�0�M���jx{���:���4�x};�g�[]}�~����K=�ϳѹf�<����595@W�5��&}4�����7j�'*�h]��h�.d������=�J3�9�$��n)���>]�-A���-�1�:V�MĬO��MS�����1i�͛j����ת��L�����?.�{/i��]��b��m�������Ժ�+'���(�Egށe�B898�\��4�C�
�}�6A�Һd�v����	<�a��qk6He��Mh��X���'IbE�9�W��:O`K�"�+mi��?$��a\��LMC��4K�yJ촜��Iɟ*JO5��;�{0ƌk�� �db����M���!�o��Ė'�N�7�T��|��Jg��7�\Q%��s��@$�_��A~�p��]��,ꙛrYE�S/����U}��\��y���S7�� �Ʉ�{�H����D��~��10$�M�,���}���Z}����SY+��
a_��MB-�v�Z�q[0u2��m*=�aD��>�#�2B��7�$�����^�6Z鬍L�������S����g;��1��K�!�(�:�Ic<��0�� ���,��1k1wz��|�jT2�rE�;��M��ȇbr>NA�:;����H4��S�$����x�g��_��dy�����#�8Z���)�{���3��6��*�Ä�H1����M�
lK.ϻ7��ҭ�EU�#ok-���âE�/�N�Q\�E�@\���-�2��PK�_E�;��pG�V'�%i�3i��w�z�0J�xӇX/'+PpK��	ZX�H�閎�,ƀ���۞>v� �8��a�-{d1��$k1?����}�(*�k/M��#���k�D��Jh1w���ƹ���p����.//f�xE����9r�	��^!������Íd��e��� �ԭ�f�R�7��.�{�\Ki�ܩ�U��g�Ny��IGe(��n,cj��w�E�=J^`�U�b�)[������Ʊ�$���9��af&�W�r��02���#xΗ�d*�U�R�j(Ryޓ�>n�ϼފ���ځ�"�
y��QHz�����LƩ�����G]����QO\Q�MGM_��/�@a��1pt������,7-� J��%�(�&���S�sv���єc
��hb(����-��������tV�A���Ĵ�ȴ�*a�~���HW�hu
g���S�V�����j��Vɬ���hYAf���/
�S�����k4��Sj�o]ƹ`s;ZwDIs���B�.����6�9��K�1�Ѩi�!w{5�PE�����sn�j�7�T2���͸Z�UP��>�X�X�%fU��Z4���������'�������o@$n6�f�^"��i�|	q��L&ܮZ��]
8/�>S���N(`�
���!K4՚>:<��9: ���R�0��+C��Y�1-	 �nZ�m������`���e3�ج�	�j�j��?
�SsO�D}�����0�ɣ��� ��W��آ����X�	�C S"��Y�� ~&Rg�Iu)șt�d��&p9aF� �D�d~?�d��?��1�=��%5�J�-�{ͦ}W)xb�m[w@p!A@h�ws�".CJ����*Иs�f�k@7O|�n���D�������n��N?�ۈ���� ��fŝ<QK>��ӚN6{��ӝ=���(8M�i�!�BA1�ҵt�X�p�2B�!���2�C<J�G�r�mٷ��4�L�s����u��'r�������O��֞u<�-�>3d2IK���rP{��o��E��N*P,��}7�m"2L�X?C\q�hkxe~*�{?T�1�nO�N��S���ė��X�L��yfN�R���_3�`n}�q�7,'ei�n����C�v�)'��$Z@� �(@He�d�	E�؉N߼�������l|#�t��xy�6��?�'�wצt����ϝ�������T第Yt��h��|�BC!:�9��<�aٕ�,ٛ"Phq,6ܤê8"i�(� kT��xO�����%Wy+�2MV�HT�2�n���|@�䳂�'��e�C��g4l���s�t� sP4�t20C <���c�U��0Tg����Fh����S�z}B##JE�L�Si���*�-����;����7�E(��5�0�QͰdމn���F�A#�z��G%�Մ����dJ��7.kkī���_�"�E��,��}b8;�[=���2�R��A� �֭\���s�d���F��;=-�X���OB�`M��ς����'��1݁�CƛR4�a��NM�Ǯ��ý4w�ՔR�K���669���zXF �=�G�0q'o_��M����|?��a�>C�a|B[Y&�X�.���tt0�H��iB��[�no�R뚈2ɴ,��������c_��`E��ݒF��|R�gc����g��$�hS�&�sA����T]��OÁ���NK��e��;�co�{�;o	�Qs{�/�'Q=m�P�󃴴f�Wxoxk� Ә�9� W���Y��ѷ����`l�-�G��z���@r3V\i	Y09��d9�2����yqO"[U��Pޝ �_>V��Y�:��<O��-��{?�d�fk���?�2%�.�PH,qd<E�L�e�f�y{u�f���`����:ΓbS�'�]��b?d�Ʊ�?O�X>�(D'��dZ�n1�/mU1�W�PK5���!���Gf�@f�<wǕ�X���q&ZJAUzV�7���{�'$0��'�S�\.>k.w��h�#�HZ���U0"�M�g�[YY�[��`�bRⳇ${��{AVQ˳ؓ+7�m��9����T?�a��G	weN��H���{Z��>ŷ�ʊ_TV�T�P��.�iHqʏ&���vE_s�q3�g�sX8%$��A��i�	��w�*p	;�w����3�~y?:Z*u�1���Q�e�VR��s/���
79��7�Jݹ�y��:xM)�:^�4�Yw��Ӫr���{�6A)P��jN�P�M[�� z�q�)�)��;O��fD<���T�����0E�ݣ�A���M�0�ۚ�bЪPv�Ȭ��:��f���0�E�B�Q��H��gHrͯ�~]ߑ��8՞7�ֻ�l�\HՔ6�D��L�[����{�g>���>0��7���ۤb+XpY�f�#u XD�OAD�c���w�&oy�b��ca��xvhX{�/g���ݒ�����2����J�?��=^o@I��	���篎��k*!��^��i[4����:��2�0�Ȉ��c ���VH�d����y����Z���=-"]��r,�b�:�0�K�%����"!��aSd����z!د����� �E�"Z� ��8��A\��!�?�&��JD<��\۽Tc��J9ք*I|�k�,�;'���X�7��7�#hf���_H�u�ID�3����兯9�zl�Od�C��6�ȊO�Q�$��$�;�0�>������v�]y�1���NW�toW��#�و�����W�y�������'dA\#�~�	��{���.�R��׊�0��!�QJ��gq1}Vۢ�	nu�I�7��*�W�P��޻q.�Y�O�(�f#����f*{t�mc����^qo��_u�'5��ӢR�)�������OŲ��x�#5N�����7<�����s�6��f���fH�u7N~�:�-�`V�4G��$Ee��p_?�$"�ƈR�;z�����w���:��HC�I$�Ԩ�֜���:�G����ۤ:b
�()5)��Y��C�_l>��RJ���_�P-��{�c����W��,�V���Qbg)P�`=�!i)�<��������.޲@���s�c�k/t�L��Nx�Fަ#7�s�̒��!Y@�Í,zFL�\�v�'�{�pWd�K��K���+&Ζp-��l�������٪� �e�WE����kE��.�a�`9��7zK7�K]�Z�y5d��V����#��++����lbN]�w�j*���!�����	L�#!.3x��/�ul����=*���r���G����|�,#���.�ń��'��I�Ma�x���Z�|X#�r�6�����]�\Ĥ��EB~�Q�ɾ���0�r2��c�3�_bS����n�9<68���~	0��_s'Kt�Ӌk-���┕�B'*�� ~ Bl���o�B~�R^ߴ���x
}�.s�易��!�(H�J�e�t2"��&���ںqPoP�չP��eF!�WbW�)��T-	�d�~��N:�f�Vm��"l� �a�k����{���� W��P���:������6l?< A|�q��j��v����ߗ#�����@s7�f�޲P��8�~��a�g>�-�Z�:�T��ʥ��9�K�S.8�-/��[��t0��]P" �����>�Rh$�Q\JL��V�u��ޅZ3���K@�
6��DR�D��r��\m'��ߍ��T'Mᗥ��>JP��5䃁����`�cj:9��óDC�]H�����=�����4)��d�c�j����"�y�D/�ii%7+|W��d
@�W�Bjq9]2P�@;d0��M#��wU�4����?#���Ԝ1�]Ab����7ʣak��w�Uy��Ʊ��2�a`�j:	���V��� FA5U
�2 ��I՝tG-i	_?����@�����T��~�i����	���7���+�覎��T'u���Rż�5sM��U*:�nc�W��&1]��3�&��C�v�=jn�Sօ/����A�C�lU�� t�l�
W��:���>� 0��J�$�-�`��z��r#��a�G6xڣ-a��Q�#��C`@_˾\�)C�^�CFz*/�ɂ�,�Y����2� V���J�԰�Y02n���No�"�}���m����&W�{АB��GP鑈�I��NfU�l�P� t���t�c���.���/��3�q���e�.�k�����$�j���g�Q��.����ܷ��$���ـ�~W�u�7M��������(􄨈���AF������i���-�&��9�йg��e���z�[�r�ޭ��J ��AY�K9�]~Kө� U�.el�p
�u%��T�Ni��UW�@(��*2���GM��1���	�%��FLc�*:��fG�H�{l��UmJ֭y;���=i��X݉��+vU�V��c�`��Fҭ��3���C��qV��fE9=WyJL���WOa�;8���53l��^7�~lgߧ3���߳3zB"vfM�&�P�"����ط#cYZ�Y�R�4U�?�����-�pF5%�X�ʵ1�f�r]�BaI̺Gp���L�_��w�-�d�2��<�a��iv�C�����J3DzMO����yy
��>���lNCD���ݻ�������k���]:�#��/�g�lC�CK�=�E���kh�^�2,ͩS4�^�B�	��K6�=9-�8�q��Z��ψQ��zr�L3k��탄`�+%�Ȏ�i�BᲲ]����C0L�nN�)��
�v4���.��ZN�w2U^�G������`���+r
0��4���a�>5��z����o�{ޥ[>:���� \��W��K�B�r�eKԞ��ۼ��y��eO�=զ��dp���k렶�� )���u;����F���E�5~���f٣�BL0T�S����v�V��=�&򧒖}�H�Nq��5&�{M�B*����G+u3��S�����.���`.5���8�q�J�Dvb�,r�}@��֙䎗��C��~gK�)uN��~m ��*1%y\�Fs���3k�
5G�Z5�۔��{��c�x�V�[�j���2���۾�eZ�4l�6���nx4�S$�C�	dt�n�`���O_��C��ȏj�׿&Ks+K���w�Q�� j�Jα�=f�S�%�?�����8���h�j�"�G~��	�kp�y�*�t��]�� �
���i��G�����v#ܸMɓ�%�hc=��2*�D��b�<�։ �`��6�rYE�}�AN����z�\'�(Oۛ��m�!-�[r��X���d�H�ȩ��dD�0���dor���~'gu�М�n�oడ��T�/��ޟ#��I��e��L]�b��`s?�IV��ػ��X���w{�`e,8-�����2�Q�F�[���v�`�թoʰ�D��$l�9���W
���}�ۭ��9/�C�P"P�f{��jAT���qSq>	�~�d�iȰWN���@G�H �ȥ�꫅E;��w ��B����`k�P��d�V���'R�#>������|���/=Z���xY۾G������(ۏt��'
%Ak�>K����uυt�#A(��r

�p�x�W(W}��+F:5^�̆A�5�@@ϭU��@���!@'s��u�r��Ҏl�����E�ڶJ��g;F���E��pHA��W�c�,M��>����:7�8w1�,�Z:zL���!�Mw�Bm�U�%�]w|5�ƹ*#2|�,v�c^���\!�XQ!u�#Iu��~?���Y�3�}M"�-�� �G����$H��885��,�����^�,����m��Lgݖ�
�d��6����8�;��~,��t������1R����I�,����W��Z�ƟZ��k+��t�P�6=�$���ijC�P���
f�hlV<��cv��~~�さ�|�Zx%�a;��%���:����1/��2N�5*~�3zVA&���Mɴ*��!��>��-�IzJ-�HwJ���bݩ[�6>O��;>�N7/k,FD�����,�k�>nY8h9�J�O~��5HT�� �Y^o��Q󦶙Nޮ��%EbT��S@��ר�P�UM-�D���ՁW�$�۲��߫li#��Ӧ;ډ�LU�������C��o� �ߚD��-��J�Aۚ	��h~?L�8�UWyh��{���b�I��VA�^��js��=�)�1h��]H����%��� �Ni� B��_�iAV�ǊTفxݞ �X�<��X�aUP�><�j{�԰RG�6���O�ӊm���_o�?*�'D��!������954"�>��gIi���	�Nl��1���x
�}��U�s���$�xݒ�[�!I6���E��w��ڸ
�=��B9o5�k=az�2�{V$���������]�<�"�\B�}f.�!�
�����g=�/��i�JfN�v�5N��_F�f�8��ֱ�V�������6)Yc�D�<t��y���kݓ�"����);����{~Nd�{��4����<~�y�!�yn�&i�~��@K9lrY)�rЪ��AN��ͦ��!ȹ��Y�A̼��>�q��,q��F���if}9�,���Ls'�.���`FDt��
�c�4�^�_���&	4����B2,[��_�I��6���R��q�~b�Қ<!�!����P1�^!YVo��/��=����u�V�����!!w5���0�9qI{�+^�g�W�|������]���'��A������_Ag��.0��v�>�v��Yϰ�hF��mL욋6���Nh����5w��2c>l)���7g�b{��?�&>��U���[vz�Z^�I_����3��@�hl�-PiɅ�3��ɓJ�x�HL��aXQ3th��`8�c��)�l�)_�T_�5�EThEqp��.�_� ��Y�#nj4�Ƥ��X��5�L�5|K޷٬=S�����R{ˬvf~I=Wn�Q΋����Y	D��Is�����>28tKt���� �+�����/9<Fr��$�2/��H�v�mwt�@0�#�-�<�4�q�AαMn	��x��~�kH��`"_��P��#�fI g-N��/�v:z�ˇ^ ��d�L�����1�Waw�a���b7��)�z�)$VO��x���,����pH8�i�<-T��h/��6`�j h��W����(T����kKx.��יB*�١��9�W�l���=��b����h��NQf���8jҪ�ԝp��Z��z %h-�X}�r�ش���P�T6?�Rs��v���&�Zu1�~&���9=Q`�8bk=[]�?dz�ҹ��p�����rح/v�K�$ؖe��^�%�����S�$E�Q��d�s�*2��ф����]�D�X�mHTs9�?�L���k" �!ޒt-�N-�5���̣A��ć̨�V�J�/��<Ɵ2�3�-��P��������hD�=�p�]5���>\kV���l��BW�!Y���[��FJ�c�ur�m�yuZ�$�F�f��9��C�{}T�[&�&��}ʿ<�Fڲ���?R�5�v���8w�}s�#��*M�(�"]��9�'k�K�ռ�\e_�m+^�-�o�#����hdӋ��E�:����--)a̿���>r�)m�{�M��
9ۊ�m:Eo$��P�>��dk5�觴�U!��=>���:e}S�A8Gz
 ����WC ��ݦe��	�e�*�2r,��D����}���#�i�>�Ѐ�2��+`�O�QY*����v.o��w����7~�Й3��`�S�wa[�F�ʮ��հ��(>�|���&�䔿7=�-�T��"�1�6�ۤ�W4����!�&w|?ˊs���CR���(Fw ���6)'Jnx�������+���˼��[�.��w
�GW��%�tz��d��ai��ߑ˄6��fU�((k���G ��u����<����L��	�>)�Vj}q<Lqz�D�j*�9��Y��QW ���уz�B��3��!"/z��勉�T{QS	��m����g�?'��孷�ޮ������cX��.ǬC�����'EQ��M�e��0?�뵁x���k���7���??m�V,Pc� �TZ�R�z�2�k�O�d�����ŷ#i�RYʹk��\���U�h	�`��q^��|��<1���)=��a�j�Y��9��s���r�7ڪ)�Z����Ǐ4��Ҝ}W�06L�Վ)�psX+�̖\n�]1�Hf�2����0�Η$�l��q�݁��Ē��w{"�u�F%�
="V�@�9���Ss�4o�o9��6`�e]������1獅A�C��X�"T�z3�śGt����Py�s�j���K���aTHd�gC�;^�ҫm� ��+�W�m�8^�F���+ ���y���7ђ� !��2�3F+���/5r���Xڪ��Ԧ;�#���{ǔ�1���� �"�6��Ht� 0xB�+�
�:�Ď�D�\\U�m�`b�PY���${f?�UwJ�mb�sM"P���'m��@a��P�/u	��֠K��[���#���S�=���0�Q�G�L3N����,%Q��2#�Q2�IyU��g�ţ���*p7���~�{��~-���'�h�+^�����43�vp��9Aѫ�������/ ���і�Nѿt�bt`h �(�;ʟ!����y;��zu.'�+���Ku؁K��Tr6w��ْƻ���B���d�B�f���Jny5����1�z�i߈,qŤ��{�+�x�h�R�Z�Fq�����Gp~�!�>�-�[u2�����2ǐș���Л$��}p���k��L32��V<�T��p�����/eșZ���+�HS��Roخ����0�<\�0�8mG�%��螛�T9;/���Q���2�(Ə��^�n��S�iJ�Z��y`;pi9�«���3��wfճ=&߶y�ksJ���cbGC�.pA�F�
�6�E�J�ݑ��2��,�>�{�p.���c��Twz�@��w-S�KFNk�v��kz�>�&�+)Z-l�fk��X�p�� 4�Z�b\(��_!���e
�_�7�<{�n�Cs�j�E�?۾�x�+.lp��w�8��23�2�նٽ_j����(�,�eB�Z���	����`; �r��4��!�Aɶ���j�rSj�����?��,
Yɐʾs���Ϳ��D��;�O�^�xj�|J��!�q@Xfa��m�6u�LJ�YD���>����i%E5g���y�8��c�S����Bh�m�ǥq�.~5�ݺ.�d�]9�"-!Y�uI�Zw�r�̺��ͤo(�-*ʯ�1�Huv������nh۝/�:NS2x��w�r%�|��	;7�n"l�DG��%�iA��m��8]��&�ƔqC�g/�]�r��Z��$���Yj�b ��q~� ��̨�����G'������u}:& �{��o�I���=�`|s����2S-y7y�˦�H�b�����q^M�똃�Sճ�B�^�z}J�G�����^�Z=�PA��B���jt��u�ѦQ7zErBp6`���i��Ja�D�Z��?����]�Y���l�_J�N"�_��%�%�Y�(p���A����
]1���0.J��}T$�2�O�}3`5]D�f�e�`��h(!�)"^f%\kϳ^:P�=&��
M��0K{��bI�������=�g�A�ɊsoQ��w$(���{��4�v:+W�ly�0������`d�I-ݻ�F>����K�]V�MU��ߔ�͢�/�B2�������g�cg�)���,R?�)���ȂtU�}� ��,TrQ���,���RvW3�Q�r^G^�Řo�)H�fK?�L����p�lC��Z��H���p"-*\�[2&�w�x
�Y���%�ⅱ4�+�m�r�#`�ߔNX�J���� BI9B>k3�{Wt}�V�x�.&D%�����u�������M��MB�ub�8̉<��H����k5~��C�-�!����a��v�D*�|_�:h��ͅ	��E}M��{���MR���h
�c�M�	,5d7y�OƵk"�5�^Gr������{�@x�<�����m�3��ٸA5�<��kB�t+��:��6�����.��j&s��o?:�x3��y0���}U�l*)g������(�~�@���S!���� ����uy�4M������>9�R��XX�1��F�^Ћ���V�;!��d
Z�\��:�g�/�	�s��έ=!|,:��]�R�B�p����7�V�y��Wl	�u_�v���)���Y�۲PMW;�3�b��^���4:e����@��@�XN����0��~q�ZQ_rDH>��z�#@��8��ɇl|��DZ�:���BZ�όUՍL�JG�P��2�� B"�ٸ���:Y1�F��7[85����5q��/��ۋ	�
�[><i��>�����K\Z�bq�l��2[�s�CYy�#�"��v�M���uR���7}�~���d�#�QCzn�Y4d�9.�5 �E6��rVԭ�tA%)ZƬf�q�,�� �'q(�8\A���Z��w�Š�do(p�J� ��E70���`�;b6rj������:I�w0����0G�����h����u�����O��E^��������`�uٗ��n��ج�ݮ���sR*��?.���a�?��@�QAok5��=��Y�'����-$��k�6�>��>��fc���^c49��<9,�2�ߑ���#�P�u��)
��A�����VYR��ӌ.��� @x
E`�y�u"�Qs�)%/��� t;���3�	0�#IR�O��$v����.��f�&٪�n��I�L�'��j����r\�(��Ѝb ����񪽪Q�4��=��M�h��u�|ר��:�W�����0�ݙd������}C��o<[�u%���d�GF�<Ĥt��˴Y0S�� H��ϔ��B�.��ù��Af��Ϧ�od�+��?'�o�֬%]����NZgi���;"�y�"�b��@M���o�{�c֫}ɵ�9�"���U���0��2��!59�@���^�B8CZE�h����T���t����P��j�X?g����U����9�9�&�Ik��>��NX5󗍩�d�K\-�����
9[c6^Mip���Um�9_���bP|�0��?�fWͧվ��) F�;�![ ��h���؛�������`��5��N���>o-^g�e([�[NO�#�����LOs]���PΫ��)s�l�|~e���2<�#����+@4V�$H�,�`pB�*@.���Z pL��u�D9�X�(�x
��o���]"
a���S
]xݱ�%n��&Aςՠ�ٵ9�2��E����<��
���^A���?�����u�!9C�>X�� D�ӯ��/�Ȏo%����82�x���s�/��x�7�Їz����x����y�:��T���o�1�ﲏ�/Z��	�[!���`��^!�]>ɐ����z���(��3?V���]�͂(�DU@4[��{�/�C�t�}M =�J!���[V��K�L�yM�b�s���Tk���1�Q��OM.`�t���{�ʫOŌs�}l�d���fUs���s#.�Z���c�_"�P�N^�kz�rY�o�Og�m�^��$[��0v�L9�K�
�Yjr(�S�_94�hA"\�`�u\̙U��F��l �;[z�4������X1*� ��ʨ�i���kl�Qdb��h^��P���zs�zD1^�-X�O�uT�u�ԛ���"6�!>�o�ߚ��v�P�D7$��h<%n��vK��=D��8=u��;�p���+d�n�މ����K/��d���-)e-����~�m]O��.n[9���ψGzo]#wPm��%��v�Y�|��T�Ђ��7�_#N�y�����0v�>��B�Y�x�߳wwx����%M
����^~u��m�*�2ȕ�!^}��4u{�nwFF�&Iv�F�l^�*�"�'5�G���np��[�i@f�Z�ɟ:�Z�w�BN�ކU3Jj�'Ս-Ay�1>e���g�{�+ww�]���^�-o�dp�dǼ�Y�)���a�%Z��U�ȹY��}|�o:#��vg׹��A'x��Ί�ց�d,7����-`�BA� ���M`[�UM�	��VEx��#�A[�� �}��M�n��?i�zD`�[Ȕ��,p���d<E�J�����"�����?4p9�-9o����4M*c5������i��UQ*2!fM������y�����ͼz����'?�Ћ3�w�"���=�<�b�"��1�й����+���4ZD!,"М�0,vӶ���P7�i{܊��^�BG ������Բ�澛�0����L�_Y�b.7��x���Ȼ+\x�I1�
�zΙs�C����·�ʦ�w2=}}�M"�p���Bf���謺q�3�2�B����53�o����i�B���%b��u�9�Y���V)�S�5��P)g�H3���җ�E�e!=�gK\�`�2^�����r1����H��J��� �:�E�]aP]ؕ�q�"km.��ܶ�ɒ�"����:g��ɟ\� ��]+&��y�
'�@�Sq�d@�*̚zA���(6M��4D^9���eK�y,�Mv�۟��6��l��c�X��*�t�W�h;wQbn\��x_WY[��>����Ԇ�M3d����f�i��o��k'(k��� �꫺avLj��%Э��6�Mt=��_V�Pu��!�&���/�_j�~��!'T|�|�j9=�eej�J�"ȡ���O��o_�ZL����ƁN��f�|k�n���^����5����1zL���.׎Dp����<8�{��c<��Ƈ�vs�~�q����]D�`>w����S��1���`JY��L��P\sk���E�NMl�bW2+N`��;|�FǯK �N�*���+�����#8a�%���g�V�]O��i����_��5��;3�ڙ���^!��%Q2��6�򒑹��:�o$0ZHX&��!�s5�S��0$l9��*���b��	6�isXj����MNc�֎�{5��Lũ��Dކĉ�����m���Ħ��ع�Z4_ܯ���[��}~��@nYu����<=���E=�o�}ö�Y(���\�f�b(�	���V�1o�k��2śn�0Pݲ�
�F�;��0���ʡ�$�Tn}v��V��P3Ο��"��q���`�7����d$,]�V�mn�rnp��]*�ypyE���'��-,���)NI��D����Y�]m:��b�hOA"�KkO46��V*�rV���x$���c!<�A��3g_��t��]�S�w�Y���	�6ኽ�"[&C��71N=�E�t�7�n� ed�
��,!=�y���7�,����L�f�ټ��]%:l��A<�T�<�M���9������Me+���[b�{"���_��'4V[r��Ru]�<M� "W��\�T>_�l�t��o�M��-s'�9|y+��@�B�?2��k�ET<Լ(vn5�8��4����Rdʪ2z"�א��1��s��2C�_t��U��� 5t��Z�����z��}���c��D���{��m3~'E�^�YKۧJL�����kR[0^ b�ӻ]9�Ɩ�:�	3,('��x����LY �JzɻW�C�7i�ԆG���K�WGc��h���*��=��vmb3X4������;��}/3a����tv�(ʪq̦#]�u�70�	ɡa7�w����nm�[�%����q���63����#�ot���c�e�r�������� �`>�%��Pp�S��z�������!��$9On��<�`Q��)P�7]qw(�����'����F�0�DE����!��ܼh9�����{�c9r����RŒu��3Ig���U��d��Y���$4�y�����r��U��og'����`�� a�3%ar��F��ɰ�iA˷z�p�e$~��>4�#�rR�W�*��ӼAO �x�y� R���̂<A�H+t��� ���"�PWû(qk&�y��66m��)Poi���㏈d��TV�uG]\K��O�~��m!4�p��|�S5�@�p(��X� ���a�\F��g�r�R�_��������R�m(E�K��p^�s��A��nU	>�[�'�qT����Ɛ���T�=��C�/A����.���2��=�F�i�s�_�g�X�2���Ü��;y�0G/�?b��)�3$SUi�l�m<�� �;��\`���m6V��������rg�q	�ƥE�۳9rv3��+��O⛜��(̓�}|'9*/�Z�Vۢ�������U�� �R�pj�=[�x����9Ux��3wÖ���E���
���Ɗ��u]|��cY��⌚�ŗ�K�E���P��,�����Ĭ��puc��u@�ݗ��7ٜ���Lv��W��i�ǣt>�&t��F�Ë����t��l����)�;���nz)����;�gy�ƕ8v��MN�80���Xe�gR�:|���l�(�ǰǬ��:vN�j�*.�y={Z���"�x�6��s4�as�@��fd��!pvbD��N@�9r}���l=ֻ�|�w ���(í�G)���N�]5�ys]Ŧ|2�0������o�O��V��Q�����=2�R����R���P���o�h���螨�����mH����u��\`Ԁ83Y��qٮ�\�n���8��3�q�x9��9���Q�Fo*����D��ҧ(l�T����]�� \��0��ڽ���pRo���*;,Ev��^{���S�|@Nv�g�b-�ø;N���c�)�:��ʗ����'�&v��K�+ CB��̀Ү�6m8q�7�������|X�܀px@��؇f,D<ЄCZ#%�u/wwk���7�3��#��$jwX���*z�j�Ȥ�(���2�i~U�m�T	�H�ɬ��xJY:�v������թ�"`�9���o{XG�7o���N���vU�5��tX��t�? 8y��(�d�:A\-W�	<`^*r"f0�+�DO���_3���Q.�v0F�	�v�:$����2M4���H�Ӟ������>����Fcp���q` 蟷�輣֠~���[w�tHҩk��nA�W������*(�!�0`ww@r�Q���R�P&�׆��wa4f�h2�9;�,�_���
q�Mt���5U�V/�R!ا�HU������G���~�Xv��qc4��f�k��l�(V�S�Y������K��)�.e��*(�u��f$�vA��.x�<�0�� 	yD���?��$���aF1�-�2���VYg�<�����zV�FK���J��j�Q
�{;SQ�~�z�}�삈��� ;ʩy�8�8]�,(E"'JK�J�'���r�]��۲�� �/���wJ��f��C6P��y9+�~'��u*���]��?��ӧA���(@���etG�~��Ha��Y��5���6�c��X+�C���}�a�\����,B{���XY 	G��?khq`�b$J�8B��ݯ���j��S��۔JYD�`�%���ԫ��1��"�KM��&�mPW���]��o!'K�����7���Q8�d]�ʶ��0s�)3$���_��2��l�7h��m�ɹz�"/l�"���t�*p� 5��$'&�l ���mS�T[�zk�C����H���.w����I�ɴ��	t�yt�ɠ rb�}������u:2-��@���<��/~4sbb\|�}a�ޑ�ZmSb�/�9xw@���#�{]%����1_,��Omo�)�P�|U��D�ݤo�g�l�����ŧ�y�غv^EUI�Wq�C����W��|+���U��7T�D]�DB��1�5X�T0�h$W�GW��߼����᫽[�!,���r�k#�<Z��8��A�N�F
'�y�ZA�Am����m�hU3G�%F2���e4e>�S�ZH<���5��Z;�#g0�_O�����~�n�h,�Y� ������ٿ��@����SN������'�*��D+p����)&�0q�!���B�ڷ�?
>D�_�o�)�x���;i���a���'r\��������0f��P?R����x͖PM��IG̏�t���hO��F����0�
�S��T�AT�ت����p�l�l�A��;�	�,�2'��#9�^��v4��a�!R�����s���\�>�H<,nȡ��pg�V�8�ɻk��!��r���׉���K���� �2�1�{�߲��?�3����	��@V�o;���ޥ����ͯǦ��
���}M�Y����B��C!���{���l�Y���l�Y1K}�i�2H�k���Zm�e��^~��-�{%�3��VjW�3��`:r�@W-�:��,��t^�frW��r��"g�G,eb@,�H��	\׎��p-^�{�
+�Cqu.0rbq�����1�\njb��P����˵�Gf�~$�>ҷ_�U8�,��pV��
��=%y�^[�@�&�r�[�����Ϗ/������q1�z�2��誷@���#��]#�2��	qXmڻ,{��{���QשKs�#Ŭ컀�>"�왚�㛖y7��w�GĽ
c�7?I�O̢�z�~P��������<�ƳO��4���A�zb�C�~t����<��zV�|'\uE�Ov�#���DZ��u�]���WG��㈻�Z�`�I��
#�����V�K�Vh�
�[��Ӧ��P�b��*���f����� 2�l�����lhCpz۽7���i�Hh�ß���5��	�Պc��Bp򶳳?пXG��;�y��ɗ�X/Td�ZA�4������X�Y����s���!��������\O�%�xQy�ְL�Ō����+h���j���qP/B>����-!p�G)��0�� lփ��Q�Gӭ�&��]�UM_:`x�� ��C�Y	�	S�F�կ����I�ϗ���c��@O�$\�E&K~s�d`!�_%юÌ�h�;�+����h��۱�>�%2A$�5��h>�.r����c�h0!����@Th<�B���T����Id1B#-n:������
җ��?�Z �*C������R3�PДe��ެq��s��~bB�%�x�)L�I&��ҵ�f��S�"����-�ֽGUO��D��|�A0]%�  =�n���dR�����׬�h�g�<k��Ғ�\vC�)n���O�h����+�՟���uPUǆ�R�9`�<X<NQyK��%ٿG���V�7f�'F���'�T���2D2��jC��ǳ)��H�҉��:"�D:3��Ok�eЈ��kV�za�7ʉ|i
힥'�\��1!���<��m��4�<:$F!������1!�ion� �)�I.�!�%$^f�5ioWH���U�hf��N��zCh�JmTxe�[2˄�IC&p��:��͋l�"K��vo�J:J���z&������!� "��%�<���taT�.���C�j�¯Ɗ�4��XA\\��e�j�
d27��Nѻ�1l��s����}�zd`,1���K����B��LX�R)W�����e���j����^lgIӟ�J�]����F啷��zW���.����f��^?Hl6��<=�ҥ����j�[��D���m3�b�Į��|��U`����(no�Jq�7)I}�گM]@�&�/6V��b�5�Q��}\{������tMzH���"�p=��o�B;����T��nԎ��/6X�A�G8�eS����.��[�_�ѕ�6U��� �L_���-"�J��8&f���r�m�>����o�39�L��y�ϑ+�t�b4
>-Z�}�c{�k;� �����YK.�)Q81�	�s����J#��^M�Ɖc������,N8��hj��B�<7~N��$"k�S��k�MJ��)U�8�/�F�U��3Lɒ�Y
C_k���K�4��י��K9��3�V�WKOW� 6�@�X��d���*y�I�ӱ�2GE��"�	���E�B��q"�|�w�q^?��L
��c&��'oD�;8��6�_/�òoj"�y�JĄ�l��=�͚���w+h^h7�Q-}ʆ��US�q�^���5�!�(F�OR�/�4��bXѺ�/׿�k5��̷r�B#W��(�Q���4���w=���[ǹ?f���z���rigVv� �;�Ϗ>����t�۱��W�.%�	ҫs'%��#�<+}�O��a���ls�9�z����T��SE�?ξ<^�ȷVǩ Q[&����Gs5H�?�F4�_�tB��I	�m����^/�{�"1M�C�����U2���͗�B�_�^,�O����-����df�4>�A��W 9:(�\:Xk�"���s�\��`�����|�#31�%�+�����j��b���]w���q��kӪ����Lc�^�ϥ�-)h��i�սm�^=�f|i�r����2������q�!�v� g�������k1���Z|�f�%�aAx��H�܃�)��J2أ�z�^.���9�Kdv���K�hS����ZX�j"�P�w�/8�㑏N>&,�[3X�[���O�"��Tj�����
m�g��S��\9���1�2x�^��ժ�A!놑��h�ޑ��Wv`0��sW��,z |M��Ȓ<�M�@�/������_s[HM'�BKݦ���Z<��~��(�	Ei��
(���TR8S�
���Z,��)�����o�������R��&���~A2s��g����[fK���*�4��7`�I�r	Z�FG�A2!<~>61�~D�au7�@���*�F�R~�[lڪM�����'�N��jQ�)-�=7���:����B[�8�.�#�������r:1B�_0��z�1�!r|�C�οlE)�)Ip)���0���z�����,ώU��:�:�8t��3Z�j!�iS �)�U��]��������1�v�$����8���s����w�O)�?|��}�\Dp�b�kߛ�E76:����C=�Qn:U�g���������?@{�H�'%e6�O�����Pz��X�cgʊ��x���*u�� M�+�.8����vQ���t��T�p����{����zT���?�ذ�a�)���R���o{1l?�3^���:��T��L�?%V�ڣ��l���
u#�0*8.�f��4S�8�5�>�Ԉ	�ěQ
5� ����x!��/�p������b�x��Q�篲�ܣB�o\��8Q��W���!e(p?��Tq�el�*0��8������Uj,���/y0���;?� k`�!��:ӕ�SA���UP#��z��峉e�]è��� T��!�����Fxl-�d��;�T6��8�6}�W��,T��g�~�nYe�`l,f�<�pIf��$�c͐V��P?�bi���z�}D�0�ffĲ����;�]2�����5��my�ض%L��b3��F-�w�w9>M�Ǣ�����(��Lvm����_K��WV��]a�Cq�uB��X�s�XI�BaiM�0��0�A�pr�}eo>-��-��T���첯��g����d�jc�F�;w���O%h�r����v�`J����2N3����4)KC.=��Ȗ�7���������s�8�^/�y�?у�����,�s'�/�@s����Ցvc��� (���3�I�{�$��i�<� ����b:v�W0�̡ԁ�7�H�<ؕ��G�~�ɽ�pK+�f�o����<�X��T�C����)�`�ڙ���'4�ºX���>�6����?czԫŨ�@u�n=&m�w�i����R��H�-fvj�~��$o���w�C�+���$j�J�.�~�e����v'���	���t�2~��U�T�ѭ
�4��VU���^��W�Sb��,ӵ=��6�2�
"[������/�W��,�����?`Z����._��n^��}�9yp/}�1����Sfu�l|'��F���Z�+��A�s"�W�ZF==7UO���Z�DkX���B �� M�ٴ����[���p)*X?�1'�	zR�� �3v�"р��3�C�2����a&���q�H��z;�{{V���}t���Cu��'�V�CC;5i�7"~�?�Zd��f���6�Z~j��e&}�R��U��R�3�i��y>CR+Ԣ�Uy��cI�M���',۠�g��&�Ob�Z�w�Z����."�ɳ�~�*�h��2�ˑ���[�oD�<!��9����fk�9��U:8w���3���N �������m0�T�27��'�?�	x�"&��Ę�KF�y[9N�ӎb��N�5���~֒1��|��r���[�Y)*?$���_�������@����Fh���{�L.���_�^�!������Ů/��u�u,��t��2��o�Ĝ�w��3���B�Tn�a"�ay�,�%���ML���t���9�љ��K3�[uyܪ��90��>X$�O���@���:��B"o����(%<K�H�eȡ,��
��i=PT�"� �s.T���C�6�nI^oa������p㣰��j���o��ߓK_9�V:/"�c�wi�}�;$J���ƙ-�q�c��]�W8�=���O񞥥
u?u��n��G�#�N��VGy=��f`@��ZP��9� l��J2��:��p"��1�в��Ɗ�hqqc�t/� l.�c0G�˸�`i���E����yR�2�7-h�ë�O/�#���>׻�[���{8)�9W�j��N{]�[+�R:�ŝw6�N��N'�29B9�ax`kוp�u����$�����4�F"��VJ�u��:}�ɕ�Im_����2E��?�B��HHN������_]��
�=M��摏�s�C,u�Xn������Z �,K,ew�Yw��q�%+��V�䂫+��5Ӵ���Q�BD$��M���3�kU��e��60ˍ ���Ӥ.��P�jO�r� �x!�o9���,�x�E��y0{ǖ��}/l������~`a�������Պ�
�o�F#0�z!�M��[3>��y:���ch8�d*�J\9Yr��6:?r�$�Tg���=�e@ԫ�J�('1W����;���ɟ����u�p;n���f�"<��r���:;�!g�:I2�Z�����v������RO0@���D䌊=c�P�?A��ew�̼����T��.�%�+4������rc����� �LVb��~w���Y��)ѩ3ĨD�w0�4/�B��25s�W�:m\Vy�`�:��:(��m�	[�4CAh�Q����d':P�����/㏓P�{]��x�Hq��u��7�e�`��c[�w�3�G�e[e��J��2��N��ʉ���l����>��reKl'qU�|y�ӕ�6�6R3/��^[!��``��;����j�&��l�~�.�e���^��4 v�ه���grȴ���-��d�햓O�nL�z��>ʩ��q@�M�G"��P�~FX��(��-�0NG�`^��;Բ[$ٹ�Dj�FV�] ��h:x�l�!ЁΎ�ueOr��H���2aTS�X��J#�6]fM�d���:n�g������l.@���X�h)4� �4�Wa�����.N0UmC�E,���Eј-�FS���! hD=������A�+p�v�#o�������.�k�����-�v)������\q�b]g+��|����l"^[H�:�q�)q��G�\R�M�b��z�S&��g����md�$U�=؆�c?=�R��\2&��¹&��<�D�����hv�i'�)������/���|�į�Ņ.��Z5� ��Q����⬲B�.�=�P���ʦ?j��x�j�]�H����]�́��%�cf�`�N�J����:z��Zs���On�3.ij2�7ـ���H���aN�MX/,Y9�n�a���P��8)� %?y���6)7Ƀ���?����E�/���BA�%ܚ� ��S��\�q%{槶���>�:�[���ю���7wJ�1C���T������S�qm���U����L�l�|��r�N~XV��4������[���0��$���ތv)�iWZ��6�1-#W^��G��(�S��.���16	�TZs<#��� 4c��ʹ����_���x�-q����������S̆���$�h�p���5�_nu���P~�E�ZrF����^]��3��l�f� �d_r�H����{�]*n^��ՙH�GHh������0��Aև�>~�T���"-�|��;
H��ұ��QuADr{�����5� ZG΀�G�Cy��sN��0k�m"�]E��N�����������:��N@���>��	Z�º <���]㶀�����:� �t/lsB�2��v:�n�H̕@�u>�P�jL_��y|���/��,�?�"^o���ٍ�F@�PwF��QF�Q�-?�bխ�G�}*�޵��������g�*���۟�'����D�<OlA\isP����PP�%	'+������΢�C���K�4��|t�7��p���JT�5��c����� ��I�~{fx�S ���>h�v��.�-ǁ�rz��#{L��0��;�7P���c�x�(���y]����� s�/5b��ؑȞ�sX�U��L��&d�:�|�c��N��5�%r��qW��K�ɂ�M��#&h�h܏���8���I�s
�2�z�60��
�>j�nj!� ������b���	��A
���.~0I%q�����+:�0_H�m�&�,�;I���k��*�q(옑z1��Ye�/X�2f�!�o8��D~�ʝ2�yV+���#�fȴ_*�P�R�(cq�S߄�+�v�+���A�is�s���'=�=�c����Y��wvs�r�eh����RS�&]1����
��m5����dW۷ЙS�(�Rof�,�d�"���g��$���-�%	���{���)��i�@��������	���]ˊ�n[�����x ��M��R���	څ��h�� [ܶ]�H"�,�a9��jw��@���G/\�4�I�^�Lt���|:�#G�tH
_����m�����b�)�紎FFZm~v�7�Eh�)�t�j�Q�tʗ�b�3ྏOm���%}�����Y*�t�e[6���ơ6`��:V7����P��)�,���Jx��c!�Z>o�%F�;��e�QQ�_Ul�ޚ�����\�'h��#ø+~>E��<r�t�Fp�b<�!|��29 ��z��#B
;�@�ÁA�En~mN�3e饳�6�i��I��/(%Ю@2�;�z@�ؓӇ��Z�R6���n���'����J��tKvm�iӦ����X��hP�Z�Y��J��������t��ͨ��9έqC�r������ϻw� �re_R0ٯ�������Ý�|;R^-]k-�ҒVe�T�3J�X��6�U��Vn0�.E����2�4=�3x�P�| l=�Ly}(z8Xh�p���ې�#���ΩmT��Z�uH��!�@�mIYS(����O�l��5��ʗ�Eܷ�q�M���dI�1�[�Gt���A����6d�Xc���Z�qP{��V�`��|�חKt��v\��lلF7��M3�Q��R��m��Dy��z�76�/?����I���m(by�ї� Ɓ��c��L�4\$�C%F�RI̤�L����<[�	It[f���}��Q�;�>��A�& ��5�}���z��O�)M���9�.���n�F*��)�g��WW`W-%����M��1�b!�D}@�{Gj�{����{�ޜ����m�Mk!���oU�wYܠ0�%t衎�|9��KXU�ƮKy�L�l�	3>:Go��e����IΗ�xjz I����%�m���w4hЂ��`b�������.�C���&�IO�M�
��)��U�$8�Ϊ��m�X-���l�ªx���#۶;z��@'b�N�ל�A8�x,wi��]�U?�������m�l��c ���#�h�x�Ĉ+�����K��9�����|��:�g'����'�.T�_����a3�&Jz"��]B�X|�@w�����
?g��*��(��N�
�{ <��a&��*rG�;����[Y-�p��*@�`HԢ\v��r��{!�C�-n��幉q,3ىd�
�n�R���/�KB���H;�*f�����9� E���ӂ��/�U�xܠ�Vd��������R���i(�ĝ�U��P�<�|�_ 
���F"�~�M�������W�dީ$,��d���$�7@�I
g�WY�,G�N���9�Y�a#";"���g�F���3j�;(�8:/i
���k�4N���M(�:�B��<2O��uVA�]�)%y8D���yy�(�
��:��f
֟����vM&6���V������D&�7^t�+7rJ~���1ڭC��k�_/O	�}ov �������۰<����;t�u��M�3h������[In/����KEO���-�����$�HE�j�p$�4��m�!���5�T7@�	Z���8�m�һ�D��;����x�aCS����mo��U� �#��IJ,�X�S�6���
�D����I�MzawT��^8s�ʏ@Rk�?d�d�r��<��7H�h�>��xa�Vք?}�Y� ��<�'��S<���d�%F�� p3�\1.��
��\ ��� X�Dz���>�2�>��1�N�c��O���W��$�l�����7ȷ��5���%w�"`'���S^�ϖ�%�_�"�t$M�x3��Σ4J��* �E�������F��ph1������p �q %_�PS��&���k����tn�N��|��-�0����e�x�U�M]�5߿��$��2w�t��v�f����Y����]ўD�G�;�Efo�|���z�:G�a�9CqReح�%;�ib��F�no~�����Z'�9x,�t�(�G��У	f�Ey�۫��)a��:mb���T���X�P����LV�t�DR%J�H �� ����^��Χ�\csCe8���Ec�bm�KQ6���-�x&aT{{�����2P�����]�D��{*cm ����czR���m۵/�����<Ÿ�����M����M���le��1�]�N"��ل�����b%�NO)�)|T��N����1��^�Y�n�����F�;�	㔗҃k�G&��9pFαk$!C�19kmG���ݞ8����m����}��"KG|�-�D"��r��]]�_T�{1��f�Bdⵥ��L/������b.����Y�7vT^����tq�e�D��;��oJ�H��n b��n��1?]�R�9��rf�c��_j���>Äs[ߙ0<^7&ͺf��ϐ��R�����+���Mf���{���W��WT~��0_0���d�M]1�qcR|����)n�[���#ʽ�� �dIuP���lěb�|�=�#g�1��s�p���i��|��&�t��j<<τ$�Ar�O���� D,�`�2�]? �ĸk]��$Ĩ��=.���~�������lm�}�j�QՖ|���g1�F]�H@��a�w��3�m �/a���F爽5�%�\-*\�4`_�w�Rn�T"��mP�NY�N�� =3$���f@�Ebc�>�J�
Z� �O�~ ��
� [e��9]_چ�a>��f��;͈�_Rc򹷡�G��-tiB$��p��2���m+���B�M�^R&��$�o�\���9�T�TU����qj�3�_h4V��I��N����}�Ս��1�G1�h#�;���9Z���� �yHP���t!0�ٚ��ǒX�����V�9��{��T\s��֦I�l&VFtL?	�O�ݒ�� @nHU��*O8��-��@2j�u5�*��g����뒿�n2�Z��ܒB��Bҿ�v�tYN��bF��U[Ì��m��M���p
�Q�e�g����'en��Z��/j���Eg&�'���ڲ�j��Z���Ç�U����P&��D!&��wi�x�yo,x��ƺS�7�u�Ժ�a����L}Y�����&G9���o@h�P�s��O5sT���������'6�Kt�=�!�� ��:$�g<�������ƮDܜ��G�K�r�>.���?�U0��3��T����pݻ\�8����7in�D�������G����vN��)T�컻�C�z������.l�RL��E��%���UG�@j�QJ,C֣�ye�G^\xT�������)Y]���?͡�=3!Mә7�$L���e���z�p�?"x!���ke�X(��t�-��T6�a�����[;��9��&bK6��m�����q�/"}#F� 	�"�h3$<5llޚ+CQXG��;�ڌ����[��[��Q�w[d�OI�u��������)�0sL�3�6���k���}�g�V�p J1�Lժ���i�L����%	S^�Y��
������#^�����<�ǈ�L�g��n���{G	��(j�-����X�����=�?����@�T�[���M ��i�bAY����d�n���6���~e��'���v?I�d
�ɓ��.@�S�v�96�&Y��(%%Iv�`��^-~ x�.���W*����ni��M_t6��W�X�RPeC�x�I�d�B�레���O�,$yO�3$5F����7�[�  ��02l�8�����2��%'5U[��D~M����!,��b��[p�~�Va�E�M~Gg���ET�~��d)F1�s)�!�׊K�g�G$ۓ�Mq[�g���6�U�u@�j�(:/3�`/ϜO��<�+�����	
\�ͷ���RSb>Z�p�%v,RY6�[��6�v��EZ	j:$�7��t��rC�^ǳ=�tZ��������C��5��橏���%U� Q)�$�A��D́�3��T���,�L�O0ƦC����q@��I�5�������E��!�(�j5�[�z\[Z�v�3�3:����֧B����D��Kn�6�)+�0<�k��C`l���h�4�A�����PQ&��k[KV���^�#i���9��Ú��{q�Tr�@e�CWl��6���f܍��V�FV���|���Vxz�_S�^�S�)!0
UY6LV}��B��9�/o�+�%oR���(�$����Y�c�%�/��-:���*ע��A㋬�S76����0"���d%!4Z���Uϼ�辙s�r��0�!���+��0<a��ܺ�R���O�A�Q�%ǯR��A4�.]��9�t��b(X���!�j�fx�RJ���iE2��0�Ur�Ҧ��yN�'�<��;e���W����B�g� ����}���r��1�m��P�������p04��\��k����)���p�I�5�������;�N�� ���8��$!Q��Q����Q�P��$.�j�L�|%��X���λ���j�wSxl:wk�J�'V�)��2��Y�h*����O�(.�v<?v}��I�\���m�Y��_��E��P�x�q85�W&9�T5'`]hZ_�@��0���M��)�Ә�L��]���w�ӌ�3�U��~x)J��i�{<��ؽbI3�b��rӑ�L�-ɵ�t,�4T�gk��&l�"]w�ǥ���2
~�\�������:Ōn�~�wo_��;�b�I.�}9��J�U%���*�	��<��rw��0����"K��0/,�}t�Z� KqC�pi`F��e��ߋ9����It*\�a!�%��Z�vM�m�Kvu�#���M�#�V����e�~��$	59�=V�8�g=�FA���4��%hu�$
�k.�Y�6pT�jC�����	Y2�bs�'�ظ�m��SX��c�M�tR\ݹ毵����m|tk��9�P?�����F�S@��rD���qM�y�v�Y�M�� Jn]fM(Bj��/�)�B�N�'M gk}���ʻ�ͨ�ޤF�_�-�S���ɒl�4s�+��%b��N��:Y���4���|�p��{�Awa�)�e?XM�ޡ���DP[g寱�;��y�denw�	w�ˆCDi�SV@֗zl�x0�숺K9�х��9�
�����0c���1W ^m�`F�x���u�Fߑ��>^Gwc� A�,�{E�sü��󿃍؀e�=mp�?&J�t�U���m���U�A��Q�b8�,H�8�u��|�K�S���-H�ʄjX���]1���T��s�ۇ�{������9��aU��"��$�OM�lLr���x���g�08���⒩M�9���6��:��������J�[:O<n�q��^�Q�vS���a�s�,PȆ������{ˇ�C�//��A��a���S(��72��%�{P)}/�%̟ؽg'��9�W��K�8^E�hx�tF�1Y)6g���,<�x�TV�x�G�]ż���)��69��i��3�D�}�F�b��]!^
�Þ�Aׂb�lkqZ��9����& >A���L��lGm�1RLEj����5y���>�V��z�*C�T�"oGD����X�1}��5I�nJC�CnA�|G�Նx�!%7�9��F����x���Ę�g�z��䍩�8�>h�E�LC��.N�K�)>Hb6�፯���T3���ќ��ˣ�{)�a�ύ�P��=�n�N�ن�nA������-����'� �j`�p4�}��^.�"4Td����q�bK��V��]hX��4h��L15�����M�����-�U��)��1놈��i�5Mp\���j�\�	�V�7<�[ʮ��F�n�ܭ��I����6��ȥ
�l�b�H&��,����ӝ�{W佳�{����͗:6�צm��D����I���+�$����3([�٠	���_�s�m@�;�hq)v����䜻M
��5�t���8�
��rGa���X71��Q�ȯ�t��$�ŀz��LGu^��V�܅?���^g�Kt���٩��8��M�������xY�A�*V����WZGU7�}tc$�N�b�H�]5,4F��h?��> Gz���"~�a�/G�r�r��Qn��ː��)1h�V�#Í���b���Fa�w~*m���{x��_�O�G��H��ER#��^������O�
0��ƚgo?+�g�����m  b��P��k�Z,7'5�u\�8�-��;/ɌO�gz�~��Z�D�bö��J����(���g�i��u��g����W�V������MY`������V2Y%H>obNǞ9�n-p�� ����`�-9cA�QC���6�%RW�$�7E ��H|�r�Z����G���&!A�q�*dai�]�`�rI�K�N���l]�Vt���r3֌ؽ��K*�sA�H����˹�F�-)�Հ%�|��3�P�  ���7) �(�(+��[���3� �V��[��"��cD���� )�s@x�,z�&��E�;M>]<a>b�A���u���{T�4yU��8��9����s}�g�7�{'���:������5ě-k��G�`��e������^u@��PL(��<��;��:G:�c�?����x>j:1�� �Dy+���m-�Y�¶�� ��5�4)��7��E�9&gx��.)���
���7�}�9K�\�j�.�q�6"Ė�3g��&aL���/�(D}FN��yL
�I|�vY�8#�
��^��{!�̾NZ9���V0sD��P�xnJ�2㉟3�p��9+�5�C$5�5�7��f�=9*�'u��h���� �H�����J�fO�}v_3���@�ۧej������1ڦ7�W;%��}�|�	��9�G:!q�/���G��6@h�p����\��a�t����y���g±�g�>��xMG�q�'��_�j�K�3Or(`��l�4�v/���{�[���Ԧ���c��߆��y��t7l��oz3���=]�<5���o"�z���\�8{�q���4�h�9w�"y�m����,�ڊ~w���g�T(�ݓOb;���dL.{�C��~���H�I�:�Er��s%zRqi�a�@�7����`����:<����2#=�js���bL�VO�Z�r����OI�C�H#x&�.�Ɍ���Lo����L�o6}U;lN��H7:к�0ӳs2��h�mf����1U��ae;����(��m��qYʼ獪�<�%��%���Z;*�W��)�Z\�M���]_��sg�����i�yK�H~��r���X��aR�U8:��P�bչ:��8�ѫ��צ+~9(�:��`�|T��j�g=�
�_uE2��n.W��6L��&s�4B�6�b ץ�L�Yj�z���Klu?�%��UPk��_23޻�ؤL�T���4�YFn�s�O�
$e�i�nP���(��H�����X12�=����x'�D�gЦj��KN��ȶ��m�c��<N����b[��G~���'�=�Z�J����[2|�k%��aI�#�nf��P�>���fu!p�]����+=VEEh륹�a3avC�hw��k�n��������㉨#�{���w��\l�H�s���n�C,{N��:�"��8{��?X��`��В�q�!�?.	�Ж1S"��?o�0w��9Z���&�Tv�vH �4d�%��w	A��O.�	NB���ϭƪ=�Z�ssɒ-�DT�(�R5��i �
C�K���HH�~��w�����`�H�[,��?
��#76�{�z��&P���g�7�}�$q���xq^X���� �7cR�B��V�Q�>�C��H����Ή�,s.����*�d.���@V&rǩ��yIȮj�>�d�d�'��W;�}�D@��[ۨ���r�H����C�s@�k��xCaxYSd�^^�0����kz/)�%po8���b]�r��7��!�a[�	ϱ$;�� ۹}�=��9����f�A߅�Z�Kd����}�&�3e�ųE�(���j �h���	�H:�&ӡ�-����f�yk�<Sa0}\�}����
3Ƙ,�ڊ�����o�	��z���@����E��뤙Ƣ[��AO��P�gA�I���)E�Ӕ��5��B>39{e��bಸǳ==�̃�9Pr��Vvt� ���[V�@&rڈ\Q�̜pkMu����_O�QQz�X�#��΢$�x*�8�dj�vҬ"��=�6c�.1�)}%��=K3�l�X�҉�����K"a��7z{����q������>?3,0��ؖ=��)�����4��ۑ$�/�����w��D/H�����s�zҫn�s���>��#���m��a�O,��m#Qmy��a�b�m�����m��y�1�J�L�#~~^g�r?��H�{��C���Q}"�]��ӽ�:��מ��qP�G����͙��^c�7_A����u�OeU���K�ʖI��{3���
�u�4m�g��"�̠Qǈ�%�f��D	χ�ث���^�~�Af'��L��q���p�k���a��3�(d4�5��5Z�����p&�U�l*����.l�.Vi��k~V�G�HR�|X���ჶ�4�LX��W{�9��9����\W0oc���o�����<� i�Z�n}�rV�A�V=A>�g�� x��M	�*��9D��#�i�-�����{��4�8Oq&������B�|���(L��b=��t]��G����ءpI���O�zHYܶ
V�f����������Y�>7]M�3���A��|k?��C��}H{�U�����Q^}6��Q%N���߄��,<H�s}�v��/����Ȩ�]tr��gZ���~v���Q&n�^�А�;y0��D���<)3!�c	őL.�ޫ@������!�rY��矏��ڨw#骄�.f��n�Q�i4�oK�߬���kš�y�!�;���¥�D�w�fWv
�&��Rc�\�&Ki��D�������9�m��GO��W\۠×驹U��_%
O���n�4vG)�P3#4G!�HԷ�����xcwM�v��Pb�N�����ͨu�{j��r�ʖ�^Kg�Y�5Մ���Ω
 E,�Ƴ��5Y�|��b��%�:�i�G�b�����/���H�6Zz�o�+7d\s/�Q�XOS��Q�9<{$<Xo����Q�T�����,�q������2���Z�{C9��2=��&w?v\�1?4���ۓ��Z��,!yi��lRU��7�n3yBA'��i��,�$4D�C������Ʉ
�E/�<���la ��oJ��g�������i���:��HO6��Ú2>=b�Z�GĜ����� ?�Q�O�$����8%ռ[� q�o��D8�V��u���چ5�k���m�r�h�#�T�����2p�	������V��;>��[��G6�i��:�B�7H[G�h��c�.����J70�����s~�L���f����zp+�ؤM}E1l�I���H�H,���'U�=!!�9$wuQ.���#�a?��6���}���C�_�w�H���ݭ�2��TĹ���+y]H�5�oD��u�����^&�>�t��w�ˡ'	b.kJ$����U+ø6�]h)�c��1�Xq����]U��uQ�ނ���}�VW" )��j�Z�{�Ї�[�ݒ�o
Y�8:�2��_2|��$��ùJy�)���S8�i$<�mSЋ@=r����7�ޮ&���x�����`DA.�H,�~�:|�#t?�R*�C�2z�����p9�gq�ev�RN��*F�+��z.޲ko�/����OC8���;��Ң\�`��
^c*k+�s�3�����"��nq�� g�BbbV�Fj��,���tc)���G����;A
X�<�j�Ԧ�nm����0�K��x�g0(j��Ŧ�2\,�Zϋ�X��3;��M��0��,$��ʿ�,7ωMf�0��݆2����}��ӹ�u����7򀳀��Ae���"�U>�wY��%�>�r�<S��֮���2:��r؉��pW���#�sS�>��	j��l�=1b�Ռ���������S-̵P)�H� �s�=]�i�s�,x�k)�5l����ˢn����)���?��g�ܺӂOP�%�&���!���dq�K�Za�h��~�������n����A���)'�҅�o2��Q�j�5N���oKf�e�����&L�$oe�3�e��!���k�����]��(�qܮ� ���O;ڝƨ�x��<�J�̠4́����Gv�>�HM�R%<�h4���4�ES��fbAV��MN�٧�X��;)82�I��f��Ifq/k�,e����Ý�7V�zT��ӗ�?ń��+��"�����f[�g�|�����=�˝i���k���)\��w��i�eZK�8kC ��Q;�"�S�#�Ʃ�����#ɦ��?ЁP�:�6{'"���u�	Z���_�{0{=y�oom�ђ�5���*�E�߃��"���rVOH���u��|�W��xti�MK}���	�~����)�U�v��A�	ٿ4�+�}z��y�MKWp�5uw;ٖ�dv���\�$���������kU-)M�yY6A�-3e`����ە�qig��=�]��p��tm�Cß���kķꂟS;����M2��V"*�(�]��9��ҹ����	�Tm�DX;�ua`����v3ܪ��m���(�{�\ު�>����&�Ɉ��(ݜm����q ٴ8���g;]t���}�Eg�v~�'y�E����D'l�
iχ�	�4�|�`?:-}��`x��]��v��eJ'��K��2�*A~���3�&���!`J;���w%�0��`�-^W��s R3֝�R��f#W[oXh�.�pҿ�Nꚋe�;b��-K�?�?�|'w>X�x�aY�eٶ��Z�9R <j���i�^8�|����C[����G��	#j6����LO<U�U��OM�E��LPf%�SdK�˽��4
�����v�z�8�� �;�Rs�X��+{�G�Z�����F4�����h�pY���˶�5�;�D�A���;r%��3��Π���UEe�>qv2�2}��q�n6���DR���P<ǡé ��2���-��R�� 濱��������<��}��q �G�MݰxeV�t��q���o�C��l�$�b������5��L�%��;������Z܆�V ��j��Oi�K+�W��K׊��!y��%�7�CW�lO!�a�%���Co��,=�*�	.������J$ީw<ȔE�j*J��T�n�����;�7N:on>p�Ӄ�o�ha/����k�Ŏ�����e(@��^gR�#��<����֢��Þ���8�)\�VHȟ���l_���C���7N�!Ƅ1~j|�fiV]��4#N�-$"L�4*�s�-t<Zdԯ�O�W�*zS�>�N[���k�����:�X�~y(�m����v��KCTjsӍ�P���m���G�
Hfb������1#�Vk�A�>����́J�d̽���A����Q���+��]'���U��o��W���o%�j����0T��E�ҡ�Al��ĸ����� l=I�Z��#n{V��Ls)S 4���]ܧ���ɑ�>��]���V1�iwb��@@�������,�w�f���aoՂ�6Bc oM���O ��>w�y�ܸ%� �p�w��Mx~$�m�J�.�Ս���\��!^P�������:ƅ �+����Dv^$׃�LCFF=E˴��=43����O%�
4Ը��ԥ�$��2�EiS1�Σ+�(��h�f�&$��5ꨭ�P�ݴ��nw{�~6!�@ ��'�e&�G�a�~<	��.b��ʚ�^��	a�X���n^=�#Fb,�*�Oa���`����U��+��R�y��<��=�B�}6j��w�;�wk�-Gm?�.�Y�*��Jy�����%I���>�-nR<���Jze o����]���$p�Q�F��$>N�9.�2J,�%o�v�o�z�<?�e�Χ�־$��%qJ�-8̫����'�ԼFi��ϗ������\z��H@��ׂ�}(�O�Nq�޸d~����Gcϲ�D����G<��gZF糣H	���K�8�X� �C�y�7Oɮ���/�oH�j��Y�X�Y:����/�Nmƛ;��6z��1���t�Z{����������D͒_�
��5I:���5<�K܈�ŏ�`��p;ʸY���vM�,S�&�7X��<q0߯�{%�YEH�ms���I������`kp�^����=�Y�Kg2�<���="{���1IF��K�90�y��l�AL|"�3Ï���M����U$<�W���?��6��n/��Q�riڦ�P�Hm�5Ĺ���##Ĵ���ouhcLo�6B[��4)q��$O>I��@��&@a�fp����	�`2�g^���+�o�2������7U�&]Z�)�"�QR
y�0]���������-,�r�R#I�$�K0��=֜�4�=�a����{̪�o�N�&;S}^��}���M���F�k��/$�ӆ�L�og}S�����䍗�`|��h[���Ȼ2��`8���Lw�N/V�E|��G�=���:"�R@�,�}"�)#	����d��.�չQU�=vd��Jyy��~�`���G��+��F5.�됥2_m]V�/���м����X�. _ܳ��z#���D��Չ�~��E�T2�N)NIA	�٠sI��p��(��r�U�z�9�R���۸HY�5M�3�u�0�	!ߣ�s9ƙ$�	����i�������b��|�*Y��3w�J9z��f΃ok�a���pL���?�ˣ��>dA�y��ͮ".����o�����ж��,���K�(�5���k���<.�7ܑ@�"A��@�������Ig^�.P��3N�}nʩ�aV/"�j��u�9��5�3��o�d��Xhۧ�Ua��O��k:5���&V�"&YS�{]�$EDkeQ5q}�,���wI{�2�L��� �Q��4��g2q5)KXw��hzt�ѿ˔�`��l��g����S>�4�~H��*�d&�fN�����F5�Q`��C��l�^�<��3��f?�j��e��/p� �nL��&o�e�-����&첞�y�Yb��(�n�ʐ��R���vm@�=�����6�#�d0"ZJ��@��Ĺ��?h����dKH�I�.)�e;����2N���!ם3�漘��m����V�1�|���sv����J+K�Hf�K��p�ψ�nje���8@~�uW��N�ɖ�yRk]�HY�(�L�D�=�O�]�� k5�����7\�;��\p�؃		����?96�����߾EJpX�A�E8��4��XT������+��Z��Ld�P�$��������ZC|��jn�� ����xk�z�݅����&����rW�4_  �Rj�JY5,�-1M�$�i�`޴�6�UO��q�vh&�7�ͦ�3 �Yg9���J�S>���Y�J,�IbבA�s�*V+�贶����w��y�R����|"�s5���4`GV��_�y�]��hfVԤ��KzQ=��T��M�u\�{n��%t-�W�~�r/�Gw?
�4h���ۯ8�2�p[�)7N�+��)z���O} k΁�j�e6�8�~�ܚ��a-6E�dh�Ѣ�\ә�Ǽ�����}�=m���2�&%�(lFe��
S8����@'��^[��Om k9�,�'�$o��ر���d���c:�9�E�v�8uB����^���o�[�N\�y���z�g[� ���L��ķ�u��@�B�����z�ɤS��`�.f�G��Ȃ-|\�������Y:���);Q(������������:�������n�B����cV�v�>|���,p<dG��y�/`�HJ������H�%��/�~%����B�Ws�i ��K8�w H���`h0O�sh�_�1;6����-8�m�"���B,`�h�˽�PsE!j��yh�I����l�|=�#q�ƌ�`�����'	8u9��G���D(���~Oб��G}�IJ�C�.^�/P��8��'�4�����L�}¸��mV����,�� �	P���{!m�t>�e
xI������G��7QI
]Lz���'�C	��B�vv�2�b;R�����:KH�hH�Q'�#UI���z��C<+eDu��{Z@w92cz�C���կ:^9	Z3ʅ~'C9���f�9g�l���d�ę?����Tφ ��>���v��<��Hq9�A'��������b��W�4��G�.�o��`���\���:䯓R��UƋ����y�F�)���D�^)>�4����Є�l��%�@Xo�%�ޔ���> `-���n��0�{ޖ��!}!`N��&��;�p�� 1bvm7Lb^ �(�{�<|	t6a�hfw�CjqlFB5g*�;^jЈ4�t廚w�k��J�җ���Bz��T�����1��*N��Vl�Ln�cF��SP4,Ң
m�;��P��i�ה�5���
���Y<�n*���~¶z+
g>��nN��M����cπ��n��F�3�!?����P�7��z��OY睂��>�COE�y.n��=s��O'E����+Z.Q�7U��ܮ���ҵx���H�BdI���`�
I���ҍ��� ���Qd7�r��n�O �Nxd3�;ii�qS( ���V�Uv���3sW^���^}B�lơ�F@�$���TͥT��d֞���2�r���(3�a1�}|�;f�	A�Q|�c$5�L�$M�Wx����Z����LAɦ:2�v�i];-d�TͷƼG*L�W��Oއ��cC�9�*�����0�F��r	��-/�xHv�ʗrP�^X����q��⒱�9r�i��_Ó\�� �=|�6,�ע]A.V��3V�L�K���I҆�Z��0�^�fRc����.���}M�(�hMY���W�V��g�5p،�{���M�[mE���8-���FG�/�c�N ;%K������V�O�g��,W����������Q�6�>0z���D�>�uAU~�3Lq<O5�=u,x?��VT� Aa�<�S�'T�J.�c��f^q)�x�Y�ֆ�n]p,��5�W#c��C\#w�<5v��=�k�Є�j�,�K?��U��N ��
�j��_�U�;{+������fˠ�z9��y5�d��lA�����cp0�/����y�$��W�z�B��� G��pZ͍�ӓ�JɈ�T[����F��%э}�7^n*@A����:#aki�.�R%��;��|�o�vtqW�y�u���w�3��g;_�u�0*sʊo�4�2����c��N�m!�/��Z>�FL�{t�s�Q��'2I=}G�%k׷$��s�~�7	1��%�x-)bF��YU$�ھ�9����Xy����,��h�~��݈XH���o%0t5CѪC&��O�S�e�����hkd��m��7Ξ����Î��~�Z_�ω����;!��W�� G`K�ί��F!Jӄ|^�������d�
�ֽ�@�0B3��~���A�r�\"9�1���4F���
|y��P`�A#2���v�N	��oIҾ�I�� ��
:��ľ��V-;c���_!SY�	-�#�I��b�ᠭ��x2�kJO��V#Ӯm����TPϛ��eNA�rV
z�}� )he"����w�����T��;2�BGuwi`�������	.u�	o4��h�=$���g� �^���G��{1�.�Ƥ����ћ�ъ(wq��e�6�-�wsD;���@3Ru��Qy��s�6^-M�&����O��I�C���fZ��+
�xq0��T�b��Y��00M�V�4�0S:�*�\���a��,��|�'YtgS��_�< ��rm��`P��=F��ydB+?����x��_o�G:Xqc)˰O_�[G�^�+���F��yQH�)y_��6�/�,x-u�z1�p���	�4�^�rWZ�^��M�0��oGY֡^Z�q4�/�>��md�I�6z��J��E��<�Eڜr��G�͹ӥ�[��9c��`>Q&L'�3���E��}Oהr]�2�E���^��t
7��Z1�3L��+X�X�8#�����L�!��'W�