��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+����=n� Lv���:>CQ����̛޺�/�,�]C	�/P7SkT��V���0>�܏�.� Ȩ����O���c���(�����6��ƂY-oUIx}��]d ��� �D��W^�xȚ���Ml�2�*��9�����o���E?������@�.��zx�=r�O@�ҡw���.$ǧ}���)�1������L����q*،u���D�l�/UGc.@�'��bI)8՗t͇I��E�I����G�T�S4qN6C���U�"$�ؗn�RzM9/%d����Am�&�*��, �&�d9�\��G�S�𭙻S�F�
�c��^�"U|L�4��:0O�a�DT'�Ck�����r��y�s�
��ꦀ�7�E���s�z'�Sыt7�NQ���5>�t�D�b����,oL,���mP�8̾Kn�1���,����p@�̷A+����?�%�f'�Ѵ	�=��;��]u�ք='C{o�1���FEb�I��YA����:B��Ο�����5U�ͧ5\>A�)�����`�Ế[/��{����#�-~�*|�/�#t�z`�K8��(��	R^�c ���������;	@w"Œ�<'��Yl"M��k�d�qĬ�⨔ɵǱ[Z* �7CoZ��u�=;s�6�4
Y��lNP� �h�K�sN.��5�<��f�?��_��]�~R���䜖�$������Bj���ө@%:�
�(�\q�K��e�j>�$�2ϯ�~^��͌�u����>�
y�d�5��ft��_���I��}�'#�	�!��j-�%�4vf�2"�A�y�{ݞ)��[��r�ޮ.��k_�	�׈����P#M#0BW�-ʃ&Kc�O��䙚�U���2�o
�~�\��*'�����qÐ_�14��*��O���0n��吻{z��mQ�,6��|k���N�4�a#�y �W����Ρ9���j�0T����ο'{{4T���P(%g6�>TK>��@��AX�<�>��U����~�vDȋ"_��z>+l�:���;�� ���`���A6���Y��`QPv@��m���r�~��m߲��z���#p샒ѯ��D��џ��V��m��Zv�R:���>g�YSn��4�c��$�k�o8i��+,S@�����R�JӜ))q��vZ��������l�����6U8.%�~�2�������DE����v��:�7��
���|M��u[�j�)�}��Z�*o�|��i�%����3Z��X?8�E$�`|w�����R׬�M6	&��=�n�P|v�i5ha�e�Z��+. o�p�qC���Rc��pR�Y�A50�#.Oh^��ɒ�sҗ����/p���̊�������<?aVY��O:a�Ÿ��	e�'���>k4�L\���΄ 0��{��H�ֿ�R=��\��vw[�]�嚿��}�ؗ��������H
�J9"�0�ۧ�B��
3J������/�b�x�� �2����C��GpM�c��?\J�&��d:n�-̌��U�T��Ш�|E6*\�X��e��?|�ς�>J����@��b[H�b�7K(�0,�#���A�Kq&~��Ж���L��
��{"�"�8�w��ǧ�d��d��:�]lJ0r���Y�e�^i�<u��+���h�I��Z�e)�W��	���`]��mq{B"s��!���3s�;�o/��E����(/ڼh�O���fIƖ�?RM�79�l<�t���K���|b�s��{
F���Jrj���CuzBbwC_&45g��eY�w�<o/U��ib�C��`UM�e�^ɒy���v��v���h+6H`,q`��8���PS������t�M��QAD�\N��S�[��f�B�(��ٵ+��T��"�ƮX�6���cj^Ɵ��3�p�4�(z����|.'��JD�4ad��pB0�c��b�R�}�� �J~ӱ�?����IF�L�t��s���ޅZ�*B�J>}��Q%��9�*b���<�������Ǭ�����f����}��c]��i���q�G.�. ��[�{<vX����lwh�����uJ�#v������}��l��ʙc+�>em	刖�� Xi(�7�.ש3�����<��~J6!2