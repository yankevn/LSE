��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K����i���sFbu��:vc�s(Y�x6��"�K����0'�^y��/�����_����4 �"�����JF��N�)��[J_�K��	ϽZ$�\�_��ǽ�������v�z�[b�C�6�i��˳�6�ڀ3�2GXG�v���o�Zz��}7E�
�R6����n}B�����;����"��z-��{W�� M��v-�2��ʞ�����ښ.���8��EJ�r�Kq��S����K�E�Ƥ��Ŭ�"ڃy����*������x�}�8^�y��2M�Opйٸs������庽�[�8��q���n�4�爉͹l��o�@��0F��	=�&�E2g"W'����]툼> u��Yva�.x��9�r� ߁38��v43�W�d�ؚ�Q�j�{�P.��I�;���khI�I��e}���p�`1�O�����P�/l�۳WF��0w<=v"�a��6j�Ζ�-p^� SI�>ff���\~�DD�JA���S��y7W�~-^sr2�&.4��m}��ZoqBG�� !S�,s`pUAOI>8�YO�
�I�k���i�rڮ#B�b�UҦZ�QؽIo�\�O���,�	P��NJ4C�MvDZΐ�t��NN!"N���,��Uh>�f�d�/"bЂ�Rӳ,�
,b4�o�[u�1��I��u��'�ؿe1�k�y?~���K,�}��YW^i�����ή�쿌�S��`�/И��LA���וP�� �<G(����T����},�Ŗ̍m)��VL]\e!��v��r�cH@]�ΈB�w�Ȫ�aXͪ���}����h���K�h�Ef'�8AR����JEU�mA�k��en#�[W|�'U��tY�E�d!{�'Č@
S�cM��qpEc���S��5����kˌo`93S����Na�d�)/��Hz�+B�_�C`��3�I�f�����%9_[���1?j�qJ���J�(ߖo%d���$L�꼡
�_��*:���jQ��A��B�؏k�?&�A�>?ȵ��TS m[Z��}�&��Y��>kT��ΘZh�Z�?��})>%4b���?%��eʆ���*'�M�K���y�;�}��%�� ��Ū��H9e�zp4����3��}���q������Mu�]BU�Y�I�%3��x���/(F~��?��஌oZ���`�nX%x�TW��dCܤ��ҿ/�B)~����jT�7���u������ގ�N�
�pNT;DV���pL��HL�9*Q(ct�t-l� 8�]:�Ƭq�|���d�!;^o���WC��͓ϡI}/U���T+�xk߾�Zֳ�)����9a��OzQ6R5�&�,������fٯ�ەTI g�'�\Ô���-N�wK��X���Z��/��L�@�6��/({qq�آ�,�We�4_�c.��al���(�LS�F�F�"y����!�о(M(Y������Ν�[�F�gT3��'�?w�Y�����4�FfԯW��kY�,�M���z�[)z)���<_���N�G�Y9��T����X�0(alw-�cO��^a�)�4:6?�z�UT!�e}��{s�>uǫ�HMp�_[@*��l��zq�@h�����,�4�޶�E�q�
A��lt=р0N.�n9��F�2$��Hr��������:\\[ٮіn5z�	#�]a)?����'���R�.�Zٷu�s�*�k[[&��RHw����r��v�9B)�~�B��X�^J�4FV��l2<��SKt)/Y�)�㹫P����^d6��ݞ�.���,�u�����i�Rk�;2}�=�U5�[�E�z�b���0�����\@�̈i|d ��q�Q���$��rm1����r���M��m2)��M��3D�\&9���#�x��Y�p�(���b�毆%/|;��n~f�-?����	t�$e^��S"i�]1!����R��1=�UĤ��&�w��( �Pz���,֒���㐕�ZIj������9@۩��(��ĩ��b���c�#����xss ��D�5k�RJ���ό((�hHA5[�ǘD�ZD�@�a(hZ��=��{����qjNeEz+�w�bn������ ����&? �X'R�>�J�#If�(]P8����6�a�^�_=��_�8ے3�7d�%�`�c�h�HQž��0>R+��;4�ӣ|jՂt�;��0�R�r������)�֎�{ү�x���[s5��>�ME��_�r(XpT��?��.97�T�|�Z��'�4�2!޽�ޒU�"K����M+� 폶��+��0'������Xj9��;kDi��DC��(���@�Ph�RAa/D��K��D� �T�􍮻��ޫd/��i5n�V4�q\`Ypif@��:4�CC�'`��0�����a�Z4���y奕����%�
꧒21����/u��=�dމ{�C�������-fD�U����HT�?Z��!;jр��j�gl����ᔀ!c��x�Ua�Hb��@0]+�X՟IM���k��?(�ea�s ����ͣ���:�D[4c$�XP���/�$��_u�ؽԡ��
���$7���D�%�yU�&(���u�ң��� ��Ъ#h�r���F�x���Gnd��da#�b4T��:Ȼv5Ue���p3��Q�Ը|�hl"��j)��:[�eA�"/��!6Yez��$(j\��L��a������L� X�V�b�{l׹B��C��]
g���NE�G�^eC�:��"��c�A���5]�@�R�.bQ\�#ء[G������Y��j-b7&�N�?4���p��sdm������tS�Wc��#��cE\�Do��*�@0JU_�����H��dT�}/���b[WHg�(�;w�fϩA��i�t���ھn���©u.ϡ$�%/V�����F�u�?����)����8g� C#��av��Į�����}��ׁu��0#Yo������W��+���2�0��!����`3.}}v��Q� ��B)]A��ҁ]g���A����$����
�I��<e+"x�t�o�K
yk��.�j	���\	�-w�JU���7s�������S�L��d��>S$�o�/�����vV����@Z&�Տt9���wG�Kn������^%�?�?�8)E��Ξ���KU��rS݀�퉍t����	�RP�˔9��Aui�ֻ�)?������A�oB�6��M�����T�2d9�Q�����0IPg���=<��n�t���_o-r���PZK��Q�.v�X��6�B�j�pAd9��s��Sjצc/�x���г��g��
��5�8c���Z9�|&ꏝH�u�3��,�vo��U��!�X�4��>�Q���#ż5uHT�(�0�֖�GI���z�F�cZu$�z������hM�3��� ��`���K����y�&~[b���Y�n:Xڢ)�9�@볕�$J��Ю&PKmݷ�LF�o������b�8��oQ`���/hvQ�oZ��>>���°ll�ظ&��:aτ�v�/���x�H�}��-��.<-_����V|	�F��D�����˴<���9��w���G�ꡏ3�rC&�}��}\��p{������-��RP��]a�_|���
��a�����I�޿�L��O�|�je��4��D��v��%Ci��k[)�.�� �c�[53R��;C�>P��3�v��s���:��s/��Ў�V J�m�	�<~β��}���05�F+�mBm"�����U���a�w�W��ʕ���a/Rڊl��O�]�WdI�T�����73���"���c����QP�q3 7`��C��K��6b;ri��O�֯+[�[K���t�N
��Ѥ�3d�� J�YD��"�X|�P�]���u��bf�qT2Z��L\n�F*v`ߩ)�+L|6��D�tL��L��%X�ϳ����qAH<��D�R�H9�6��28�[U:l��X��^��`�摤��o%oh'jd��\2���A&8�o��ΧL� 5gL�'�f+Zg��|j�N 5��<$w��8�WG�끪����yj�+������S#�)%+ �^�E�u\+'�L�YW����&v��*&�BAHsH�x�!���fo�@|tH��b�%�=)��̺t�>�֏8�p�D��n���'�[e��d����GN����/y^l�!�iz#��/~��BcF������k�2V/-<=ʎ�>3r颰616J�2�k����L� N4��4
S@zӻ�QaT ��{fs̓m6�ۛ�ě�M�� !F�wid�c���6#˯��v
�G����X��e����Q��AT��SS|?d��s�GNA�S��mCRыq2@���r�a�=<�l �'M}ҔB�'`��݌rO�k�3rД�]R�#PS�8i�uE����ߕ��a���E��J��Z(��E.��`N�P���?6���R�{j���#6���94��^|�����$�'L���3<�BZfm�>(�
���Ԕ�H�Ā6C�ڐ�=wN
�JZ���x��MW>�v�)d���ǲA�ӓ�2$΢�)HU߅LJ7-�Hn�5����/2�B�a�uY�� l�#$�F?/���3�UA���|a �:p6�o�Ή}��禣.t�s�[�Z�_��$ɍ����Lь@�(��9m~j!�7Ml#N�H�~��KjOAZtB(��Y��Cz,��tܺA��ǂ��O"�p����W�!�1�������7u��+*2��.,�oJ�T�U���T?,E;�x��AT�R�$9��Uh��_G+�7��_�p�C]p���t�P�`| ��ڔ1���z��?�jZ�z@M���_�$�^Ay��)vc%{䛱T�4�{'�4<B�Hj�Θ��c���=��T�U1��T�?S( [���Y�%�ݜ;iv8t"M?^�v���v)/r�=-VMVÑ3��,s��Lu�����q�݆"���q�#��l��������Ј�&Z��"e���8�uO��:-��n�M�3l��^�}�Cq#��6vQ��JԶ��&�<��;SU�S��Y��z�[j���r���*�N�oDL�i�/w��:.���t!�]r����Ч�q"3/f�y Օ9��/�^GU�D����t��2���.H-�yo�p��ױ�TR0j&���Bж_�fD$YԆ6?���c-q ���K{>�˰�w㢆SX�mY#�b��<^m�V^6s_Oh�(��z��`hƷ2����׿��x1f�`�G�[�[T��T�����ɭ�}�Ec�z��3��_��É�!}U.'fuc�EP&��@_,Q�`pB�]?��\�D�\�ǌhE����|���ZZV	�'���C����ꌎ�~��{�m�J�;/G�y����oQ��/&2qy^	�;��ퟭ|�۴xQ�xP�Wۏ�\�S_7Z��D������݆��l�۽vgCzH��7a�r��¼Μ�����M��56�����c�����JX6Z"��^�o�����b�f���$g�d�V��i�����f|;��>��-�=u|�Ӻ��X%�U;I���F����	FF�,�:�玭�g���i멏��B!큦��_��%���'A"@B����d�.Ě��V��z)|�>�zv����+�����\�&�#���5#��?%Yr�E������q�!���s����*��;!?�Im3	h ����*� ��I�D{�$��m��Κ����Q�&(f��I���~DDS���b[i�qn����ѳ�-������fD����.��7QS�ٯ��
Ҟ_m¯����ӄI��:��2���4[B\NԆ�W~D���c�O� �VG#�>p�!a�GA�S�K,�T#Q�����f]>���'�g�CfI�0��%Rݚ���Gyg:h�om�^�����8��F�I�&����Z��5�u"���m��ӂ�T�@Q�bu����M<;�@]�Nm<�?	��aj�֖PZF�H*t�q���,�\<�?�A\�@T���j���Æ�w>.�zIuS1t�S������4)K��u���h����-�_�ih��Uf�m
�|���Yg�F�Tא����E��#U#�{���J���{B�j�
�@7�7b˓0����(N�_D��I����HCV̧=���>$Q�5I^;#a�5HM��u��j[���m`�U�i)�U0��oI�3��l.�V6e�Lr�p�M%�O��Mf)ϒ��b#�� 8�H�u���%Oq���7�n�)��5�����U���F��Ԫ�C����byo���:tI ��J\jÇ0�Q2:�ӂ���;�|UL��r�d�DȒ���'u\!�U����I�H=9�΍}��4�v�)��O��w�m�FU�q�ޓnon�jͥ�)3�����7��Y�Mb���w�sW���B�ٖ͂1B��m�.7q'�Tf����r� �F��&���,�b��CL��]�	��1_`�uax�$deVF�̉0Q�s����������o�X��{k"��Y*T���*��<G\��Tw�,���-[_?@l� �Jmb����'C;E\��"���+�,S)��)sN�ɺ��*s�}�4ͣ�ë���d�,x�����Y���u��+">!�[J��jx��c��~����7�8��R��΍���hs����抝bȺ���h��3o� Ì�<Y������H��Ǽ��{��{�c�A~ۖ�O,���;��#�.�(H�ͮ��yc�lC>�}Ҫ�%��� �G��p�� ��o���˴J�G��Q�*���KG�C�.	�3h�6�R�ee0X��.�6i>2��!4�1���g"�w�'���z�Z!�� ~�s�a����#>9c ��-�-�aY��Fq��t�y��K!�e�&ܗ}�	�x}����u������,H�X����L�!��a	1K�V�0�=WrȲ�-�Ui[Ʉ� o����6;�ux��^�k.�"�}��K0y��" LJ�'�!USc�a�E^��^�n1����Ό"�ȶ��] [ڀ�a�@���&f�En2NOj��sX�9��N�-�'+¾����@�Sɉ�c-��a��*�=J�T^�:��xμ��U��jKT��R�&ab��FL.�"�Ґ��nL1���p�G�)���𚁿��j�C-�CՉ �8z������u�b�$_�-A����f��nx�/Jz+���9YX0���@�&:2�h�׺�E8i4}0��Z��Z���ja��j,eї�r�e��8)����B.��*�pV���eEME�^3�hggî!Pu�n7u �3���߆��Gϒ�-� AdEb �$(ߕƹ(�ւV�d���H	a���A��Ȋ��R���8�����/8|e·(���쓛��J[�9�Yأ7��V�3G�P=H��,?}u�@zL�.��̱^����t��G�+�;ԞmOs�bHܷ�V���w�bi VGs=~)m���Q������	�)��NVf}���!�� �	��U;�V�"��F���6I�&��	�*Sxr�r���{��%���29�y������p]�חv�3ZnŶ�/���8���Jޮ�n���@�3�3���,@�KC�?�;"D��:��gU.����f�o?�RA��޾�Ou�OWAx1��V��6�7��%��@y�砸P6�Mxӌl���23v	��M&1Q����Ei/�,�x\�AgU�<�q��%�fZ���	��ʒ�Ϋ����Cr�C�7����d�n��(�mm��vg���F[J���?X���&��s|^�[� ��ϒ��鶵���1��[����;�!C�&g��S�(Y`"IR��|�?u�A!?��w�Ӄ�	�hm}�x4����j-���ݰ�&	s8�'v�}�N�bV7��'�/O�b�x4o
K��_=��{�6��!�����^��(���F,�~dp���f_S������0�p{�;#��_�}�5d�dܐ]VT��8����g0"5�H?/}-
�B��}D�90��d�-Gi�/�?3	i�ͫ&�2y2��roU~� z��6�����"v��z{Q6>6iĂ9n	��*�^ɸ�1���N�
M�G�q{s5+b�{��D(��>8��?��4$@{�d�,en����xz;-3��������P������r��Fb{Ț��K��Y�;(��T��Ek�����k���i���+m;�>�G���wy�M�߹E��:i��������-rN�ǥ������>^�#A+o��q�9��h! n`�A���{O���n��+�\�/_� ���~��h6C�V�F���%܁������?��E"!7�́r�E�k�@�o�g����з+!�JL��*�l\�Gѵ6�j�A��UT���,�A07:���R`qJQ~���������WC'���ڇ8�A�6��a
��kG�f�HJ`@%�\�sW��fUȗ�"a���I$�3�=����+R��1͇gy@o��iy|׻K]e3�0���y�Z_�}��4N���w�A)���`�nAF���@�n/������k�R0�V�;����Ḧg|�<�x����P��T�e$d_�H��r�* K"!��a'��5�VXZ�=�2���1RL���۵"��_��$l���p��Z �[>��~��p""v�.
#kP �E��d�"�֯�g@V�|2U���D���~g�cl�S��v�����l�M������R8DQE7+mM\B���N�s٠�$�M5X1�q0��[�!�,�M%��hl���x�C\���<�[�oܛ
O�;�,�e
���������B�
� 0]=#�֭���K�Z��dĜ�靁�)�P�2�۾"k	�[�`r9#Z�^�TEu�!�����=��"���>�?����uKG(4%_7����W��@<��Q,�ad;��",�A���Γ�_SB�Ѹ��o��J��yS�=��� VD���msK��8�"}���#R����~�m���I��qv��W|?w���Ϝ��w.��<F#��0����zڥ.�8O� Ǫ���I|������@�D���+^ �m��h(���񦮧�9���t鳨�iQn
�?z��q���Ȱ3�k>0z9Y�~�S=l+shm�s�Fvs�B�`ah�R`0i���Q�	�͇UJ8]}�Í�����.�M׳S9�=�@"z_����&��!��&,�߽�H^��Ò��1=�j��:2�:��QPA���C
Pp|����v���^��brd|��5Xc��.~���[|0�����b
�������G��j��V�3 ��}�1�v�.�t�$���m���AvB�O:�r��=��'[}���� j��ǈ���_���̕EM��{�7|��ښp�F��,���s3a�3�?;��?A(y���@Å?�K���v��^\�=
�\P��H�$sn�'N頭�oJ8�;l�0�ٸ���{2#;i�Y2/>c�u�f]�M�۹e��?�����Ζ��5I d~�<����/�?�+D�6LZ:�jX���m�X
,Y��#����w}��Ib�x��}�[�����kؖH<�r`"�!��퓠Xe�m_G�o�3PI�E��`�e]�j4������%[\UH븏e��9���J=կ'��=�*n�1��n��6ݍ�M
97lQE<��+�,k�he��ƴvx��vF~p���4��ܻc��ݥXv�L$;������2���a��$�x��[x���n����T�Y�d՛�7Y��-LT�"Zn��,���}���hy4!�\��S\Ԕ�9v u�l!�|��ъzp���k ���ѥz/�����$�����#����al�����*�Y��R�5rX�͞���}� ��B��v��P�Ic~̉�-�d�
	!k�Q���u)v$��)��Y�`�o��}|�L�J��4�ʅ���u������.��R�n�X_ȝ��Th=�D�bGC�$�3��`|-[�X�m��0�}�Z���<�� ��n9G�	�o�OS��X���uGs���U���	!2�g|�I�S�>z]�`L!�����l�К|�__�RM��+Ѫ��D���0����v��͑Xh!��A��_!�H<���#DQ�ބ��I��"�M}��wֿE}�d0�27�_Q�>�;+/.*P<����K��㽛��A�O�k#�;���.~=3Ն����>��[A' ��k[G�:e��"Yih�c�u�Ew/,n��<��2s|�w~�A���n3{���].�.��Y&rA0q�T�K��u�֕�w�A���8�R�  � �v_����(#%GԾ��wRE�7�5��J�����;�W?֩��5���Ac��@�Ng+����:�F	���1	rK�/sm���̓���a�}����૽��w�{&�\'��Dw�P����S{a0'�)����x�^����򆵉s�7ڙ\��[����J�\�a��͞h�z!��_��W���?uV��O�_Ai��$����cau��椨ܦ�K���Ʈ������C�Z'���GEs�I��ȿ,=>�%�OV0�^�����Eb{gf�*Z�;83�(�?v%`�[���n���N۹]Z�*;�����p=���u�"��WZ�`�Mkn>]Kn��z`s��-��9�@���5�����t-�Q��_�@@�}�H�Yz��o�xe�����0��D.CJ����eF��KX6��b�1۠�Fޡf��?g�W�.s�?}K瘺��r�j���XF3�"B�Sv�-���'A���{>��I����:w�?�����K}�i����5t)�-�j1�VU$*_fJ)dKE�b�!Q�(���$�I�է/v��R^�#��h�n�������]�^�����??�|��m���NM�E�b��̸���<��^�
x_N!9��Ѻ�˴R�,t���!��S\��]�Yc)��ZV��V��}5�N'S�%�H6GY��߈����p��jR��0�O���R4O�Y����z/��Պz�������,
�zE�57�v��U�cO��{H�3��W��M��GPq�������Υ��	r�W��m����o�	�E�1�ӆg�����b�x��o�-;�=�����p\���z��E5��z�b�Zhe�.	aȆa����-���32
��LL�oF��T�nn�F�������j���oF��?����` :�jRA�Ey�M��?��+�(A���ŌO��C�X��V�hk�X: ��^X�
R��G_vU�Ta��� M0��$$��ݍ-9-M��Hm�v¡k�`��hOA�xP����k�#9IN�I�8r;�ys�ߚro	�2�
H�����8J)1{J���]'�<�$[��i�I3IY�B����-zN���P1��J��K�71<�g2�t��a�N-��b�~I�hp�*�Ƿ	���)�WGK�L������|R�� �CH�`W�Q�n�Å�ݸַh�����]�Q�_=�Fځ�"S�1YB�G��1b�r�h�#&�ZI���C�~�V�Xdps��X㞦3��i�qY`�A�R_4|��@w۝�p8u�BD����@�Tm���A�����	?�����?�#�詣��P�WQR3^��H�,��8�V��ن>����zMj*���A
I(V�p����Vs���U� ���<J���]�B"cO��V���I�7ǫ��`�Կ��qC~��_�H����*�J���~�(u�2�4�<tI�G#���ߗ�/?C��������b����?@�����6GY/����_��P�[x���i~�V哻k	=uE�~��)�s[m].���4�l�L�5�аؾR��d�FQ���O����bo�U����C�,,���
�_�?;��٬��������g�nx8O�K�尃D��#�R�zo��簾*��,�fv�w�K��I�#��U~R�9��0��QY��O�=2�1�n�:��s�UHT-G&���J7*"�řu��s��vbr|.G��@Xo�h�6�v
��ɖF�A�\�E�%�a�m�I'��� �5��b+@�D8��"�T�}�4H��
���|[��i��{��$PB�;�*G�։&��
�A5,z'x��a�L�q��_*��6v���T����l6n�5����ߤ"�_�E��������P�*T��y쀲2�A!R�$�z��G%V�>W~�U�F��_�X__��~�u]� d}���f��^�0�b1�g��(����8�[�d��&�_\m���$�%x�7L~�p���B� Uu���N���n���0���Y7���\��gH:���ABI���5auP�:�1�=���=i�`B�қ�K��!
Fe��� C�q��e�޾j���Ƨ�.���Ɂ�I�F�?�5;p�7A��=Mdep�	�q������`~��� =��O6J�>�u_��{�z�<�WX H�uS����Q%�S�|�P6����"2|�a��$i"��^�ȗ3g��8�*O��Gf��a-�'�K��R��y�l��t�[o�G���9m��V�G�Ͷ)�J�zs�d:=EOqֱ�[!Cx����e���zL��
�M�GR�e�E����f�� �[
0�P��|f��[�Q��_N0	�f�����8G� ���#�3�H@�l�iT,�~U�� ���H&C<��N	�4ጮO �gyp����x����z�.O��L���ۛ�G(������L��+}���X��h�F�<c��(!6�e�o�}�"����&iY�ïb`��i�����Qtb��y'��v�Pa�)Z�wF����������y�Ol�]T*��-@�yqd߇��ŉP�F���ܼ\�y��ڥH$D���船6�����53�d�b[m�=%��0������e-$1A�3T�������4�8�r��om�m`B$p�c���Xc�tr�*�3��V�G�l��Y	qtH� Ȅ	|�b�K���k��N�-�u7r���Z+�9��dQA��1��G�8	&���y��_U0�F=�:�e�}	���آ�;�.�}�mi�1
JƘ���^@�� 9��fB�]]���>�p`D�W����`���X��]�J�#�$y9h�T���<;Z^	hf,��^��b�{���Ry�V�4K��Gc��a�6�͔`Rd�g���-�꜉�E��	u.�^t�t��S��r�_��N��h���z��rI�p�����A�D<��I��n����)� ��=�vwuVi]�#��		Ev�
E��CW���B���y�������	x���c����}Jeʬ���J�Q�M���o��t�.�6��G�b��G˺_���8@�`Lޏ��c =6?W/��%_?����#�B��Q��B��Ǽr=���%
�y�B�X��G�!g@�B�A�I�=CO�FN�T*����J_���*q���Dʖ�눛P�(P#�~����*�{�[��JR�3�$XV��n#�Ƭ�������ON�)&\2]�r$pz4	&/�ݏs��4_r4�;Bs�:���鎸���~����o&��F����1�ܱ�h&����q'
��ƇI�TY���~lEl@D�����z�v������:a!K��xy9��Q���tʷ��(^D�F�5K��)0�!ҋn;���>���}�z����/m��ǅ�J�P�n ஈ��̾w�Z,�����-�+��-u���ݙ.���:��2⭍�i�K�������4ꎁõy].6nLvP�"$ϼ(
lⶤ�c�xW`�*|�٫�=̉�;S�	��v?����Jd݉Ül�7l�s�2&����#,�s���~��QQ�ga���� fn���rxZ���@-�5ZH���`,#�Up:��:��/������̢z���2�3WHdWj�r͉:+lv�d���A�y%�f�KҚ�E�J=`oa,G��˔��U��X�"s	�e^�-��P^[�i��]J@l���S1��� ��};S1n��c���m�[�@���d�rn���_���kDZݵ[D�P��'��ǐ�Ī=V��$!�᮸� �'�v��Z��Χ?d�/Y���G�&	�����A�I��W�SJ�*�������j�ڕn5�����vX�t�22',"��B��W���0�0��K��PlHU�\����WGᏎô��Q��uUHb�I��0����Y�����ݩvl��a�pը���7�|M�N;ˊV�W�8��}�p���'u1�aH�/hf/)�\���q��9o|�2�@���h�>�}f*���.HԜ�A����Z����W��W��>�tOS���{�!рʭ^%]�jgw!Z�{��˫g��k���i�+q��0�F�,`C���+��!u�u�i]������)$�|B
�`�˪��p�/��/{0}楑��,�e�dz�銓'�$���N�������dBо��֕I�M���G�����x�q���@$[QE��_0��Հ�( �v�x���4�R��������VO�JUw�nh��1��s,;�Qjev9�/���]����'Ds����k��1MKlZ��.V/�b�#_��D�s)�)�YГI*F�CG�}~�R0-�न-2I]���'��f �>���:��-%+Y��� ���ӡ��r�v�5PO]Ͼ�8��ev)@~Fǡd	��D�{�sϾ������S@[�� I�m��c��W{��g��f��:t*7��Y|<�>��F���ҏѾ� k2G���f/���b������r
�S�V��6>TԍZ�$����C���D���}�k����y�~�tC���.�%��� K��H��NWyW�4/	��r��wwg�/PLrP"_�eNA���лl#����<1��J���m���v�+�C��w����a�����p��2<ӝ���E��F�m��6�Lҕ��b�譠�P]id�hS�d�
��#T|NM�Z�}t�3���Фә�]7R�o}�]=<�'�]�����4��\0ko^=L�{+�d،����ܔ���&��z����)	Y������c�	�ҷ�~TBP�6��/�Y9POT�	ao�J�-ݸ����2��GC�P���L�f�����iINW��e(�%�tqA�;���k���(��&�+��g���}�x5����aB��z��J�xC�(�|6	q�4Q��e��G�ƭsд��<��y'F��S=���E����lk���^�U�h�7Ӱ�C�,�t��1.=�[n�D��ϝ)��*�B�*��~��'��e��$��?=�p�T>5U��_r4���Uz]9��Б�e_H��Q"ƺ�Y·x^lI�O	�M�͒\ǿ��ȁs��8�`ӿ�䎟��U���\��U���!�6�"��D����rnj��KG��B���X%�P�SlO�G�,���w7�+`�����էN,�Œ�e�qM��Q?�ڦ�n��q�+�������H���M��m۵�:m�#���F���-�<٤�y�i׮L���3�j���l��cMS��ԣ%�F˖<������i�Y��ׄ��|ٯ� �N�>+)lH�i�}�{�~Ko�����߬���E��VG�ǫ�2�M�g)�;!d�������N�V*�$� �y/E��3�+�x�ѧ�>�/�j+aZ���@Y��*w1����ÏL�$URγ�4z���K�����"�r��k'q�����Ek�s~�rI��vlJ��i�Y���F��aD����C�|���}	�]�D����[nr��[xߜ���8�L=���B���DO��!*��S��K��CN<4�G�`�����/�4���Q�����٥��8�����H>�D���l4?幖�!����1ְ�:��p6X��\_,��g�[(er�=�avߒ,�������誝�R~�@��;��Y���;}n��{1��_�I��Z)�}�`�i�	��Kh�-�rpd�?1�&�^M�F8��[T�dMV�;G�BPǾf8�*�`{���W\_ ���A�?/��7j�Zd4�w�45+Y�c�~3�5
����g>������Ԏ�$Sl�Q��)�z�p3�"kz��x�چSA��=���&���Z^�zFBΠ�Ӏ�&Wa	���֎yd'	�Ds��m�����!��H����ߗ�NI�u�E9Nr��?�e�i�"M�K����5t3�� ���:iT(; :G��ub���mܼ�AT���r��k�y��v�-��@���BwT���~���P�R���z@�U�;H%�ek�u���F�L����]���0�Ԫ��ɧr�����ە9�/<���ݒ�����X}D�7I�����ƿef���rx������M�ׂ����0�}-�����Т���w��!�8�)�z����hXT�ڠ�lת�Jd�7�Yo�M��R=-��	�`�^w���U@D�qN��~�_��D�v��	���W�E��tK�{.�4��Wr\*�9r��o%&�����n�\_tN��R�΅�&�R�qZ�*[����~ $��&Y��I��D�e�6�z�Kc��1��d����%��O��^o8�_��UD�J��цid����lF����J��p��
��\�o4��^~ ���qZ�D�!��5���E���� �� G��%D,�`}?3�}�^�Ǉ�f�Rp��̛�Vb��n0�Qo��·XX7��W��K�U��&zQ~K,�S#��0�W+aQx|��+qf�~?P�J�g�-�i`�w*v�<��]7������Q&���nS��)�.��1{Q6�W��䴣V�W�>�l⨔s$��O��5�Tq�E��*�֨�׌^�9�縒8�+���_&�H�{"|���/JW���ԝ'���᷅O��CY^��-^�
%����yǧ��;�O�G�]��eWٶ�����=��������0� v{��Mu����A`��t�Ҥ��}��[� 'SΟ�]u��B�Ll&	��m��f'5u��B�'� VȬ�Lm���\��M"�seD䊗��Sf�i�ի ���t8\W����3�Bٜo51K����Ѫ0$�-KM���6=Ar�X�5�kхJ����J/�?���O1�$"�O��^]�%e�A9k��/�S�i�>(uPˈ$IAp�L��Sb(�z��`��;��E[��a�bq>�\��Xx��O��-�{<���� �-P��Чs�r�cT�=���X��)5���t(�m���U�kަ�b�}Ts�&�tЖ�u
}Q�L.��2�C ߎ4EN�a��xP*��	�����>ET���<���<)^�&�R�����81�G,-xG������y{��0S�S�b��[A����)&d󈘟'�;��'��̑�An�ɦ���`�*�s��lJKd��X�b���#�S�
�//l�n��B���$��J�œ�C�����\.��Y�j�p����(�Jg�~U6H2�3-$�}7����{a���ր���x�V䍱��=�I:l3���k|Q�W����]t
�Ռ��LCX;�V�!C�k<��ӱ��p����tgp��e�a���H�Rk�!D����{q� }�f^����T.p���8kk�S�7(��ز��٫p�k."ɓ+GK�m� ��m.�4���'6�`Dz�'�-�G<rNM��AfV%��1�&>����d���2��Gz�����0Cͧl�)L���\5�oUP%��ۻ]�W����Q�?�3D�j�D �臻�D_���X��k���.��0�1�W��j%��%V�5���_������w�Ќ��:@c�r�����Rq\����@(b���o9�`>:b}d
��sL4ܚlc�	�j�'�(�q~=�m�*�p�$z��r�!��5��i��v����(�c	���� J�KFv8"2��b�󜷖�~��Ϯ�A�@�G,��?_�?�}�Z�4��8Ki�ܞަ��6mg��Ax�ٸ�T
���6amζS7�}�J���I�.V@8J��:�s�ɖ�����h�yV(�;���T�U�e@�O"��	�^G�I_��N$�s���"��R=8�s����W�!B�Č{|����W%�,D�#,h7N)�F��A�F�e��y_cI��0��|�M
'���%B�K���K�x�F�$�Ч��I�uc뀵�[�ǋmכ�[�.2�\��RM�NN�c}��u-�(�	"ݼ�q1Z����F��PW\�N��*3��$�����=�$c�Q>D��k�1�88��Į��O���3�Z�w�;�CnPK��h`L�M��y�k�_{�v��!�<���o2�O%=LX��Ԫ0�jH�z���Ұ�����x��Ω�ZI	ӎB����j�� �k�g�2�[�n�����H��FD�'���o1���+6Q�0k6�F$���G�j_љ��%餃@��t�A��(����;*�upSʪ?[H~P56���-f���H�����V>�3��sK�U�wtb���ɬl��,�a
�m�\�������I�>�n']�xJ �D{��&��)�#;���,�������n�I�xӷ�V9�:�!��:�p\���i޷��[�o�钻� ��`���T��^���^��!l��n�Y��)1��U���*(Iqإ�� N�Ggh�Y���r�
	p"q�M�Fx�j�=�9 ��"d�����0�ϑ+��;u��\��P�V	E�������_��Y�v΄ƍKP�#Vg����{j��R򥦧�kK�l�.g.��ה3��/�g`w�Wo-�n����j�t˗Q�Z@)�U�d�r�zJ`]�D�Zo�x�+T, ��[}+����p�'q,��X��NP[��ܮ|Wv�م�^�#b������w oͲ㔆@�|���r�Ty���[ϕ0rS�Po)�\����!|na@��ZZ��]۱��G谇��<���7���D�Q�d+��ZF�?�$�P�+��g>�}�����f�����g���7c�E�����B�c���ᮭI��ɶׯ�Ɨ�h�\a}h�8+�Q ���	���6�\�G��X������EX����C�ۉs���f����:	��*�E�h�(�����6��Z� Ǭ�V����9�<6�vnC/	���tU��V!�Y3Uޗŀ��Lx	z���E<�xvn����5��#q}ڬv��@sl�/ �XX��X�������[E��`�2`�P؁Tw�E�j���LEG���j��>Zm�m}d���h����)� 	�������(�nO��E[�R@:�$���Q߇�o�+f��)�"M0��y>m::3��w{�.<t.���Dvpn�W�+�Tbn)ԙ�q'g�bd��o,�^�'*�o�=#���s.)�r����I�<���9־;�H�wO�/��O�����t�h ϳ���Q�z	����:#-c��o��(���Sx�6�
�yn��8=��=Z?؊�	���²�� v<�����GA�?a]Zu��1��i��ԋ-mD[���ԛ����vy�.FZ ح�;4�:fE[lS� ��q�
Ĩ=֞a����dFO���E=5��?9�5_a�L��M�����f�Y��*vs�C�W�?�	��<%�ůfzsP�$T�<fMxr�29���XM����$(b��f����,�)ə 7p>�:F��nؿa�� p������}����s�$�n~@��6Ҵh-�SG=$��-�j��a�W ����
���NV�:L��b��FCm�+�*ۏ�ĥ�v���͜3Ţ�*��PQH���c�   �"H��u��V���(骀���B���ѵn�7ē�~%3�hG�9u���7u���=�󽤣�2Bu�>ڥԔ�3��_:jZ����F��E)l�tI���ʐ]I6ά!qrjZ�eQ����ɀ���I��[#�R��q�b=��\�="�'O���bz�>�0q�i��h���Ԫ0��a���<���w�;�i���>%V="c$o�-<�`ò����d8�@Ċ_���|gN�jC*j�9*�����qBF�虿�׍��ȧ���Y����}4b��dv�Cm���z;3������t���0����Q1�KI/���p5X�#ǹ�7b(�K"�1̜Qh���D+�� p:�����]-���ߴO)�I��Ýa3/ߍ�tJB�e���ײkΎ�d�y�﬚I����C��v~-c�L�l\���گa�#3�iOp�d�u�q�OI.u�:_�컕�9&^S�9�%N�ڕa�S]V9	�tYE�B<�*,%��Ba[ g���7�a�9
zn��:���3�4@���ד\愸cگ
{vt�q�X����~�*��9���,Gث��`�
�b0F%���n8�&�5sV	�>�������~���_�5�L�FA����J�(]'2	9���b�c�
��M������I��oyⳀ�S�9t�.0�c�"����	@d���7�U#�Mh�8����YUZ?3/��$��s�$�$�m xҽW#��iB_��,�`m�&�t�;�/.T�FW���c��]?�I����Z�L�ء��S_v��A;U���/�T��e��d��kb����۲V�s��7���!T�z�I�ٟ{��@��=Q�Á�Ii䎋��1m:|��)�K-BT�>G���/::�)-Ŏ�8�jkO&�[����Dr|�@�����w~�15t(1	,p�̻�[�<�c{�յ� �%>׏�d����2��.�!�����Y�Y�*�P�J�k�"_�����>�Fw��uMC~�K>�DP��95�r��ad�.CLZ\>�F$�!�]6}g���YN��r�6�6��t�޸��D��:�U�D�.ĺ�M��>Y	[ܑ���3Kφd��7�W^��f1�5>��*C@F�h'M����Ѝ�F�;���g�����b�o��u��q��k�<�h�+���n��f�}�k���a4��#���k��h���V�hT�Æ.���t�hL�� �w9�R�Vӆ]�:�~���x)��]�O��:�c!�2��Z��k���"��1"�? mxh���Ӹ��8O*"Bz�~E�'r8���K��R AD��REN������w�X�A��N�O��i�����HV�'~�q���������*|-#;���\�k>�;�+\�`�'[m�a ��b�bI�wU�5���<J6`0:RHp�������/ab �~�m7�媖�&�{w����/�L���y�s�ʞ9^6AN_��`�W:+��q����w�m����g#�h���0���kկ�́�M*���:Тש���*�[+��/V��
P4�CM�x�9�h�s�����۩�G{\eu�9fƺ6����C����dK��[1��`���I�ht��'Z@vћ.ݵ���`-�⫑��lQ�I�uU\YK��,_������A��$9K�`o=�n�*�h�A�Mlt�ދ�(.��?�k��-��W�`�h(��s�Q�5!�[ل��di� H#���b�7�W;�h����*�@�V��F�^�[���g/�$}I�Nwaڜ��τ4J����P��j�kWfZ��5�#85�����{0I��0/Y�_�]za+�8���o ��O �>k�SUQ!��
Qe:���:8�	����C�o�������3zy��`�_B�������נ��ݳX�K���NP��_��I��hؼ�RZ��w�mz�=ų�����p�򿣢售��1�u(6�CL�=ֲW��f/$��? �xҳ�J��w��?�)g�ŝ�B྅� Z	K���vK�i��Q�㵅���X��So��5\tDk#}�����gL6�I���01��n���%���-��y.�5�vf<x�s �bC�L�j�ٻo���D�m�t�q��oL��ƃ<��NJҸ�ְ����0�s�#�v��j�n�w���ϕ^��I��.7�&5���:��u4�^M_�}�@/gM�%��t��	�^�w��h���Tܧq�AhQ[�Y�"x�b�6����YWə�ET�a40t���0Au�dC
�E:��#�4����M7s�"��u��>��ϟ�՝E�(f/������|v�;�}o%�堢�8R`�)���^���^m�n���N[��D4D"b`���ML�f�m��e�L��T��XL�s���,6��sÍen<bzG��Q۷�7��;��O�/	����*^I;:ck��-<����YQ\��i�瀐M��gOUٿ��f�����uo�h��f[o��T0"�G�'u���ee�E-�2u�0.����W�r�����M��2؟�,��#�eX��-\z�C� Q���-zM�#	�H3|���fsE����
T��J-[��D��*V���Y�	i���Ey���p�)���,;}7 _�{��k��]�-8���?%�J���7��kd�.>�
̷�+f�x��@�/�B�K���ҡ-�s�<K�X�J���ەF@L����<K���1��)<��Kr�or��jug;���.@�_��C�F�.o�^s«�,ˇ6�#tO���R�G�d�/So!z�����ğ�ɯV���l�6�}�Һs�
b��i探YR�����	���L5'�Z��t~�V豇c�?]�t"{��v����:?�Ơ2$H8���m��SN�/�*%���U�[tHZ�	 BL00k�����zV�Z�Ҕb#�ˇ�˺ϩ�XPrޡz~�d\���@��K�o4\�a�� ��K;4pmt,����C���=.*��yD�VE�p�AP�Vqݜ�bN5�u��l��eϳ�C��-�@}=�	��l���-����"\�uZ�F��S���J�Q���n��Y<�P�H�,\f8��uyX]�`�̎	�#N�$�j�ٓ��m��9� �6��]�t/@r{��``6�z�lZ�T��x'	��H��̜S�t@f�eWr�V�r�d��sS��a:�Q���}�Zd�+Lr
�ќz�-R���'C}&�o��咐$G�z<{��k#o3�LW�x�V�co�uwq�0(�^�G���1��l�3���%��/�4�>D�����U�k����{['�fq��@���x�X�^oiH$	�p���}�d�*�v�0K:�EI^Ά�ΉE�
 >����_�����UHj?n<�x�i(��=M��5D{�G
��G�n�7ZL�WWyg��v�cra�2ŋ�}&�Nq�o	/�I��ȢL�Z���*3������S���rS[^� ��Hб�ńﵴ.^׉	���o.wT )�\�cM}�����$6e3�������ȝM2��NU%4��v	�8��΢�F�T����臜}��2�Ft��E	���U^�l�Nn��u�`�d�G�&*O�%�����
���]rw�]�
@�_H��b<������ �i�KǱ&��-M� cLIlpK�)��@�|�L�~�]_��/X^�`�� �ݔ�:P�G�/:��1�`Z�
>K%8o:i`?���[����e�1����AD�
6��`��g����	�:����WqyF�-����_c� ����� �ߖa�K��Z������DW=�����L�Z����o�4���gx�,��n�w��x��9iQn�iLn�.��A�˾��}��&���=;��r�c���G�Ę�kژ-,�!#����z�Z&|TY���
��c���I��D��h	�-G}Xq\�q0$��q�"�`#��$<s�LB����D�p-�>hI���P���9d���ĺPi*�k�`z5O<kGQ�b��X5��`@'����O���Z(�`�4���=��6��Jo�?����H,r�
ؗD�&\�M�@�'b �T#�ogyJ��l�W!�~�N��ն��V��������[���»ˍ>�=�8�2��n[�R8����n0��ܴ�c�Y-���kJ@9t���h�?"S��uG`E��>�No��H��4���2���;�܉����:?�oe7����,Hw��NpD���f �"<�Nz��?m;�oU��	���+�Qpq�CY�����S�1Ʃ�`��RA,�U��f:o(�������7�Zț�DN���Ō˿�L�v��c^���l��X��#i/1��6��f�a�.�s#������ߓN�^��
�䬮'����۶Р���DO��f	��@-K��j���ܾ��ˁ��[U��T��;,�s�iM�km
�7Om��'���IWX#Zɗ0$����Ml�j��:�-fj>���Q럓8	e���;w�ȇW�5+F������ҦP�P�=�g���Vx�_l���VSY�Cεf����T�����F�gVUa�=�{�л��UrB�	�T�s�a*C��o��Yn�q<֘��Z�6�(���� �Dϯ�A���T�Spa4�Ʈ%�\��hn����KbT�qT�ٷj{#�-��&��=�] ��:�9:-� ����J��bm]���*�^�t6�jX�Bsa$�ys��(��(^��z Öz@NJ/T�$���w�Ǡ��G��s"ȭO�it��[m1�c��|�n���(�(�ɸ��f#DM���Ͻ�������3�LP-�kC�����ΰ���V�$���*I����������g1���S`J���p�-��w��E��Udy�٠D���q����/�I�$��|:ћ/�ė7��q�^�|�8Tp^��#v�w-qɺ��y�v"ێ((�#�i�+�m5��MG}Q��E���hJ8�ھ���~P�Tg�;��t�`�b�������(Ko�\>��KtG��lYpu^��G�.����(Wjy����K���A��#���^֏����@q��cZ&�Z��OS���ޭg̖�l�-kv����SI$&��x���ȮC Cl� p#H2I�\awD�#��
��X���]^q+��_AZ�x����<8¼�c2�q�m���4d�䷤i�� �M��.��f����Z����@+Хp��mEtuE!َ�����ĲA��ǘ�$�3�dX_��Eҷ
�m�aɺ]2�n�$;BOΧ��k���_'>Z�_�v_������S	���ކ��JJ������� ���ֽH ��rqL��H���	�.X>Rѳ�8���2Zl�4	&�l��n	��w��ԍ1�����T�d��ҋ������	#b�	������?��
�|���T/E�sHZ�,�H+	A�2'o,�zW���?���U�+ �I `��}�D,��aw�?��y���/����z�ȖS˪Om4R�&�����{��Rq��b�4�)k�gC�om[�˖{ʥ^z4*o�l��������%Įp 9�U�x�>@�o�o�¦���Y�)C^HZ�G]aڝ�6&�?��!�W�Z�Ҩ��潢"D%7U�l��TiK��-���m8�9oM���=�ﺡ1�m�𴪓�; ��a�ҞLR����J�W�g|K������c�}.z;*N�d���K}#����ɽ�hI��A�;(��/�n�h��y-6�����Q�({��Ě����HD	s�_��H�$y��3 �:�n�A����`�7��Tf��e����k���W6�A�cK �̺�9-\�Li�|�J�����X��hx����T�H=�̇,^Ȑdڦʀv��K�e���_��I&��*-~�����]������v�Ԕ��2D�63 ��nc07Y~n�$N9jV��Ai�E�0u"�:�(���(weY῔-��-�ə]DJ9[�Sw���=�j�}�P0p8Np4���1	m��`��
n�&ս� �X�~gI�ՃH9�Y(���u�t���f9rC+j�]�vr�f��̎�c�w�$�ւRӴ���:*{�~&TΞ�S�W����8w�U��r�Ro�0��5qe��G�g(�Y(B�@�L���Jn>. U�u�Gd�dM+Q9��Ò�k��F�Xl"��:1�#�A���Ĵ&�w:d�dDL�Ll:a)�G2�~�h��)�)mK�����C2����}Ė��$�����%�MzPz�£0��f�aVr%���Ub��#I1�욇ڎ�k��H�����pd����O��G:ļɃ2X�ITw��bXl�BA)7%��H��x��Q���\۴3�i����	+�[�xu9��+�w*H|K��*�7�ժJ��JWZ�.�!h<Rq8E��;��#	��d�-��d�fRH=���Q�a������,���Hȿ�45|�F�N�'��21f�uŚ(E
 n��*�GQRy����s|m��n���XX�#sȖ�䕨q��Q{�R_���9϶�lkt�v�����70�K>�����1�K�e�!d�!�Ў0c䞓����r�m��I���!����"�o�#�%�7�g����z�����e�\L�������r�:ua3k��V��ϸ�H:�Ф؊��jU���
�H�'�+j(��t�i}��P�M1"����!S���J����p<|�8�sf��"�Z8pzJ�Y6�!��O?�:e���n/
��w#�-�yU�j��74����&� *Gܰ����=��>�>,�ы�\]���K�!��%�z�ю�.��y�����E�uʘ���z��Z���4�y'�h��Y��+�6eO�/Ȃ��ո��ɉ�$I����#g�'����nm8��k��J�SW`dͧa�apj�D��Ϋ��PK�3etX�l^n儨����ob�\��kl�/�ޞ�e20�er�p����J�����en����H�H'��L�c����l�F���
�i���N��1��0$R�x*�a�s*a�Wa��	su�P:S��8���e�,�S}ߛ��tz� ���ˆ?LtkfF7���-�����>a��\Z:�IO��K��$3j�(��]d���M��W۹�?��j�o3ʡ���X�t��l��ZT��&�z�E�[�fk!������c���ŏ2p��0���Tͦ�LU�#��e#ߌ�Ջ��*�H!�>�P��D�[�S� �U���-�����ܼa �6�n
��}�,�5-<���}{W�q�U���G����s<��%w��P��=m��@�_�[�u1S���bY1.'�Ө�1�O����U�A�� ��4.�S� Ħrln�4k�iON�T?�M��a�l�%0kՂ1���^Q�����l%���A�l����An�.%���b/v���8��j�iۑ�[�s��N�I�����9�ƀW%i���������J������
$b[�0�A�Iu	;���U"���*4f�p�;�t�RFX6�<��1�i��`������8� 5����ޖ��+�m�{|U ٦��w�}H�j�YV
����$���p�iK>���{yB!*�Fh*��}�γo�D�k6]bL��-���ף��W��SVA�7~�fa��q�U����|���������So|L��u���g;�Z����h>���௩�Н1�����t�4P��� � \�י���C���5p8҂5�����i�>��4�5ȱ�0�3JaV{�z��<G?�{�1H�^�7�u�9�L��Z]�Ә֥��Eȏ{�5g�AC
:+�	��]�}�-4�+�z�a�b��\�yx�H;`�	���ދ�f��y��ur���B�0�p�}$�L�#�8 d��Ϝ�7�"|zo,��p�H-ѱ��F��k}��$���D�Ac��K8��b��Jϔ`n�	s�$4��C,���i�X��1��x?��F��j����$�v6�YG��a�I?�Fp�g,��]g�E��dm��[�deU��<[���@�J@H݈�ڧvu�?��U�T��������<��d:x�;�4����2�?u�M͛�] �O�U׭s� �D��S�>bq����Y�ldU�%I��>��hRQ�R�5e���w����h�;���P��ׂ���H�V]+�Ҍ0h:R�l�1��r�%���`�������I�G���=o�f�?��G���spV��͈_�"sx��]�<��j�,X(9�3�b���ґ��f����8�x���|���L����B����V]<pg/�+Q�ܔ�n���Q�V�ޯ����V���)�B�^�M�I��]v*7�E���<v��'Da l����R|�S
��20�=f��M3\^�D;���\�F*���q�fPW'����S�Ƴ����qc��g�@h��6����f�/T[4�������xO	N{�\S��򚺂a�Tp��1c�P �š����)�n'G�4���/�@ĪV3�vQ��uǍSy�O/(-�z���t���rQJ\n�ڐvr�i�區�	�׃��a��꽛>�2�ml��W؝�G�F/�(�͝��WdR�n(�D���E���q~ e*ň_5���G���1�x�p�?�ҳ��t�{�&�uD�Z��OX �~�N��92N�'���[X
।S��-$�m�'`Uӝ�U{B[#p��d���쨸+JM�N�/'� 4\<G^�Y�y�;� �l��7�hb�}����J� z*O7OO�}�/0�@�}��8v�P67��kǋ%ϢT�����@J��v�85[a��.�~s����_�s�%��%-Kh���4$��n/˯��(�}��-�MV�n<��N;y�!�JO�0��&$��3��rG��v���@+1��H�����R�ӫ�R�#7��$پ�;�t��B��%i]t�$����V��nP�>��n��ә2>�'��z�	�Q��2��V�R��^�5 n�#\'쓱�c�S��l���>ȥ�U��ߎ�c}���i���G[�UE��lų�����Duy��z��q����q�w9;Z��YЩ3���<�G��R@����7^���e� T�E|_��F�Tw�ţr���̵#LU�\�ӳ��J��p��B�+{�'o��4u�� ��hn�ýI���m��!��qv��ѽyв��)�W�O�iK���~�|���)s�&J�sA��{&7ny���G� ��寈Ep�f{��%馀�������DWRa�C��C�=sQ�mg�.Mwz�jPP��*���iK�	5��5wqY�5�ȓ,��E�p��{�k87F�_N��I6Z�>���8��E�:q�����0ц�o��ߠ�w#F��*��������s�����Bƙ}>�D<䳦=��+�x�.��V	4�Յ�z�hS�i�9`�K�E�L,b|�`=<Ƹ��I A�Z�f�G0�)�k�0��-}�\���ճe��s'� �xʌ,��u�"�"	p��~����)�'^�٭vn8��!�*>Y���g<�&�+�._�nw�Q�����'���'�3t_=���<����%�J�a��(�X��5� (�?��y����0��>w�q�o��}�c�K���6��ȅ �)&���E�O�w�����t�@�AD��?k�k��j�ְN�l�����M���TE*5�r���c�������v������B�T���W�k�3pgZ>�T'7�����TN����P����b[Ɗ2��c̿��$��p�!Ix�]N;U=�X��[�����)�>E5J���+�Y0�l�?�]�c��I|���^�A�<�k�h�t���a����J�(���g��U�1�1mojI��25�R�|ΰh!�fՌ�s��W�d��/���ehFˋ��	�E����	tޜ�*��E6����Z�	�/�0 ����֌ܼ�����_��t���1���O�R�ȳ�X�z��	�h��N�����-h?�$!�{�$�$�O^��ܖ6��*-�������NXb)tC&�����4��Y�6�¶��򒬅�����WUs�f��b�=,��l"*�Zhsm�BZ��N[I�dX�Iu�e�r������NT��\i��N��GD�SgAE��R��Ѡ$X�\/��S�Pج�����f*w".�yw,
G�ը+�/�PH݊'s]�b�SdoaS�ĭ:��t���l��60��'w���b�0_5c��a̚��t���|��Utf	J��k�I��v���U\G�e��iy3ј�0����'�2��n�2:huws��dD֨ 석���	5V�"�n���-5����xXJ��+��wB���@��a6�T=�!��l���5f��G�!�He����`�eG��n��=/���duh�Դ�����k��m��[�����Q���a���H����)p�\7�)��M��Z8.�b3q��� !�1��J�p̓Fr��2�[��ݟI�3P�K���檬g��#��3�A5)8�MM���>��.4k�O����|�����������d� ��16ѼѺ�܀��d8���� Bl�yG}���b��%
��y��!,�(�(��&�U���?	�e���bQ��'�bE�/8Pml�X�ƝU	B�YZ����#$-���_C���j,�g��~�cM�Y��2�,[��K��V����Z��2�e�3o���E��"ǙJˑ�B6�X�RSWV��3�h<	�""<q�P����ͪ�*˵���H��L����ɣ�6G��Ϙy@�����BZ�1�qCk.ܣt�B\�Bi����Lڷ
<�I��3W3���߫��ҍ��MI$9�s\R����['-Ă��E���u�f��E3�F��R�ܢ����H��5x����R{�I�&��N�LC��#p��*j)�R�T�p�g;����bo�3)�4���ģp=;�C\f/nS�J�<�{�w��~�]�ݢ;	9�M�G��q_D}`�<?��Tj/\� ��؛���X/�'g�,.D/�)��`�|��U�K��4����2�611�G���B|%��S�<�s��fy& ~@Eà�q�\,��qL�`,���}�ޝ�͖��N�sX��"}	C4.I����m�_p�Db_m!b?�] �ڈ��7;;���&V��m�s3DE���}����S	�i�ſ+����M�
,�q�\mR��Dx��D8���=���)�uu�|�w\�F�/���n?���ШQdp$�T��c�%��v!��Th�k2'���,�� Lt�<���{C���R�?#].�O�c�ڡk��6��q�����g�''�f?'yq%��2:�&�sM���ԃ�g��IsY��>!@����,4�nص�i��P��u��'��Q�n/mz��|P:�ֳQҟAq��X���K'�`I�C��nB��&�}���0���k�F̨r�5^.0،���N����B�hUY��$�B��hۊT���?8�n	Jxsh��	��ا������f	�'j��^�R3&3�q8�,�y���+�M���y����^g���SyB׆�F��9��:V�
Op�(p���!3JG��u�;��nm?t�-����]*`���p�����BV6�~��7i�E���,K��$��Q�_D��2��e:b�JnRMh��j\>�
����qz�3��b��<&��`���:�?�ՅQ���@��"4�ny�n�;�6]:��TԨ���#v!I/��J�Z��w03����Or��~��Uk�(�r9FW/��ڰ:�kg	U�i	�Cztᕊ�M#$c���f������s��o�8�pse�1R #�N�I�ؚA��a8�kJU�w��,��V�j߱H�v�h4}.	�_�PV��r�9��n[����!3�C9�5{�yO�u���K�¯��@�~qUA�2���
��H���~Æ���d�Q��٫�~�@���8�p��|�<$-[O��[�P��&ꌥ�ة�����C��J�߯�9S(s�2�&�5�N���N��C� �w Y���<b:u�+��U�0QX1���H�ƘM��b��nI��L�<W�|!E���(�@dB��d��fA��i���o2�w���\��r�D���^��ӫG��-)M[�̤<�6Ʀ.����ƶj�%9\b��ͣ���r:nc�,�*N���a�2+�w'�ʢM����Uɓ�%Vfd���g�c��n4X7&�a�{ �l���7���z�xm�Q����4�!s�f<� ^���8$��<����K�+�t
�����w����ʞv�[��1�s9v&�"�ͱ�6Ը�X̨������S�0�~R�$dr`P_JK�Q��NQ�φw���F��J���v�_ߞ�詊�k?&�����cL�@I�Z ����}�NO����/��r����:�͆n�8����j}���[HŰ�z�BW��o�Y��5�e[йi��8Is�M�5G��
-�}x��+�uީO� ^�b���`,�5Xr��f��h��]��ob��}�<o`���k�:��!�U�?*^7n���g3g{E:Z�&��_���D�&���V�����M�L�����f�J��,6����DFFt�^p��S���B��o7�Ʋ��楘�L-@P�u�� �����mS��t7�VP�hP�0vl�w���ϧ�KZ��P^6�*�\��}�5�S�����S=|�|�>�#��!��+v� �)��e��w����r���(#Ø�at�sq�������l�J0u��1Ĭ�7Gh���R�e�������ږ���c��?T˫���P�E��Ǳ!�MTX�t]L7�ߪ��wֆ�n��KO�Q7���g�xK�aZҀ8uԧ&k�{k�\�;� FN��FƎ� k?���PX�r"��;l`pC֞D��:�Q�������W�mE�|p��a�h)XDY�h=�+����w/��D�r
~����si����p.�ݸ�qUe7��<N����.����u�M����'`s�/6��t�:�B�5{��N�5�	L�)��J��7����t��������[���I٪L�_�^��2kt�����ހ�^�����h��(yQ���@�ս�y�;}�h�*�E�vlNB"�g�·���4�bZ��+Ǫ�L�d<i*����<8�=�³��ѐ��ɡ�8O�e��h�k�BI����`�.QHtF��>nO��ğ�K+tp�oC�c�! �[J4�d�B_��-��� Hg`��9Rhɪ3��D��I��"��{�:�֞����H0�O�@2�ꗕ�R�of�ϯ4�RwD�bL,��h[��.�a���,�un����}�X#'˖�K��l0	�
}�u�"������Z�c8>9i��;腝�l�ҽ��+�>,|�|7��J��~[���
H圃΍Se�rx�OHl=�����Wf�]}�.���O��A,�kW,���� ��̏�]`VZ���i��e�D�->o) ���%�b1{7��1�,��&)6� 4m�1�e<�D�y�vC��:���n> 5oh���;=D��A(���H��d�a>����^-�ێ�a�y྘�ٚK�:�vw�8����\�=���tNg�4Q.Yx� [�Ȁ� �>����i�5�0�Ĩe�+q1�<9p�Me�"���r]�u�k��`i����� �{8�lN`QJ:E]�,��#��r�K8��Ė�FZ@M�-+5�u�i�hd��[z���?�����������)4����=��ȳ�o�*�s�TH=Ap��&���bM��Ҫ>��}�n�N�������n����ׯ$+��x�l�:&A\��M��h�m��H�N&�'�e=��T2��D�k���1/Rk gp��G7����^�sIA������Ü�c�_�+�Y���=��T�S�gxd�.ډZp�,&��2R%��2����8��<�5}ۯ+ˑ��n�šT�G�jJh��7�O�̯8��Qq�ɏ\��XS9���lo�%I$��ܾ�#�k�|�l�)}'���Έ?2w3�a��W¡%��
�lɁ?�*����8��N��8�b)h��XM�R7���h뜅��S���&[�W��+�k���ʭ�=�|���N��cȈ1��b(�Kt���}�6bM�
� 0�!���Z{pE=D��y���{&Қ�ԱͽՑɾ��/�p11��0�7�&vG�+A��,9���EU�oȆ�~K���8SշDZ�8O��ؗ����/��� �~���.�mh .R+$���$A�)��H�9E��_S�W��8��c����N_���!ccl����R@_��{&= ?
��g�b-x#ķN�퀕���:��J6��'l{��)�ϋp-�A� 4�*����c䥛�}`�C�Xw�t��G�V��`6z�� o?�e!��F<����dXYXp�e��d�J�H�u<�{���$�~�M��'sVaSGsÇIp͛Ѽ_�~vQ�@ϴ?C�7�����Oߚ������f���V�Z��F7r�yVB�2���u���O��U�N�9�i�L�_�B���m����x88cj�"�Y0����Z���p��?�'<0�:f�_��͕���+��S����k�������ޘ�`�G��z��FDǵ��7�d�z��ôw=�j1���jB
����2�]� �]�T������^�B2p+�D���Ȱ�H�Ӆ}j-�ZG�B�	������w<;ͣ@s�,i#�|E�1*�Hh��^�l���V�{s'��[T�����E�3���ڇ�h� :N����i=S�����)<�g��Ki+�dN��>�E��g��	���#�)�'-/{��/�bh�\g��$�nج_}�j���� tu	�݀����k��*����������]�jx7���S9bOś���pi /�#0��;?>9P9�4�D�H�ф�rJH"dDOV����N%��޽3)+" �h�Q��*�ʹ�I�A��P�yz�����460fi 4��EXAԤ���e@�Bz@�32�I'r���)8��{Gw����r��]�����e��z8��c�i�����t
1u�'֍�"�kT3?�/>���dF��Z3^z
�4�yZ�Q��!�B�Ԅ�*zN��O������eӮ�t��LBk�] m$I�4���c��x��kD�M��Z�9a��^�T9_}����M�̲pd��9�|w1���OJn޼
�g�M���F�f��t@�A�12A��r�����d<����0Hq���&��:��q-��@��QPog�Gez�	X����`�˖ �U���R���@*�E^"CڐmOɋ�)	no�p�
�,�b2V/��D��]����[�^�[68����K�+ctʂ\�|�Ө���S��7��W�<�~���l���w�(��	��)�����W���Vń�T�]8�	K.�⓶N�&��h-�cms'��9�kl�	*�QUC�"�$}�|jց�|����[�X�y��e�,���آ���ˍ�L~�ꭐ�I���g��&؋�_e��X�@�E��������'��z����AmO�$����عQ% 3ø~c4�|K�|����/�¬
}S�{�k��I8ea�iiZ����?���>��-�3[@����*v_�~�QeŌ����ӏ��Le�Bӛ�?06�)�"t�.��Ek��Q1����b.��e���Ɨ6P�&�'h%OK]PY�uۃ�35�����w��t;��(/x��Y�W�D
�	~�,��(�4�gN�k<\_œ}<�*����(m� Dc̟�YmQ
�L���^:�BlN����#��`�[>���`ża����b/���c�Y�?�pY�	�>�lY.�TEpہ[=�UR����h8����v">�l�����Q�{d=��?�̩VW>`)ʈ:�S��L��:��lcr�h�O�C���7C�&2�=�F�U����'9�1������Z)����_�RK��*$N�^)�"��r��R����M5+����;��\3Y~����:�_�c�?n�_m���L��|�+�o��齉jA�y��������`�_��z�$s�(� �s\9�5Ħ�X�Z�F^��� bfdX 1�Js�5��IR�>b���lke^�ı�k�ؾQߟ�8��uNr�Z�ü��:����@��K��6M
����bL8����k��D��@I%�xc}��#bJE��a3Rxf��fk��Hp�ޜd(�g �5
���rM����JV;xb}��v�<�.�F���w�Ғ���z�p�f{�0POf>Cl��Fv�S�qqT�Q�쩑�XV��t�!;J0��u�~(�'�1]D4}�K9}�>�c�F1����JN�ݐ0���F�]��3s��ᴛUZ���x[�o�PP$[��uH���E����̲��:GQ���!���EB���BK̠��s3�PQ����Jc�G���Y�@>=}�������[��k<�h�G���1���S�6�	I"pw�P�	��s�v�K�dF�S������۵��r{��e��6������2�~Yi�/ag���_p�������Dz�sJ0�I�x|��ݎ};"��F�S����;U\g1i���:>���#-f�dxm߀��	�1����wW>��x�盆$~�H�a��0��7����'���uJEO8�б���8к+J,��U����)��A�������{������`6g���]�"�e�(��i��"/����OG��:��|�_H��a��+Ώ� T
�������Xڡ��@�&[@_Pyĸ[�v0oy׫�S��v�)@��s���b�3`�o�Ee�q���vz�s@���I�?O	�)��u-6���U�pJ��ϣw��Ʃ��W,,bdhmL�??�)o��l<ւ`h� Q��{$��K��W1������ݎ����d|?�u	����H��_<���V[��n�z�Q����56�5-NH��
7���y��,%�s�Mݏ���w� O�Vh��Y�����B���!SEK�E �>;���#��"�w�*�]�Ꮣ�I㕁4)���VѷԂ�W\�d� ���lBDmG�"��7����3 �X�u$8@t]k����}+{��䴎��#'��l��c�� �����'����4��l�g���ZU�5�߿�UX�p7��.�0׀�lxv����w/��2�gC��D*��[�@��V�Z+���S����F�4A��l�Uh�	乏?N���v�@͸��R5
�K���g�=��@�z�JN8Ҧ�,#xS����X�����l��"`Q�B	�or��v1s�� 6?F)2|MkBH���-œ��)�"�𷇏;��˃��#�I�}#�j��N70b�+G,k�i�b\o���?�o�<�+I�6�<���ؤ�\�XL樆���X�Dkcۆ��|P�]8�$�S��&r �,�JG�����͛�}�I
EQ�Ӑ\����y���5�Z�j��#�_.������		i��|nC��0��kK�آ�Ȟ�I�\��l��Cc�֕ո��>@T٘���Π��N5%#8;VU4�9u�LFqϞ"���u�Sq�m@f�5��Uq��|w��Fc�y��K�<kR��Q*��K����A8��D�(����Z毪�خ⮈ �a��e��ksĽ�:z&�I���Vf�'����[�}��6�n�~�x�沤
�D�a7c�{5��!���X�í�5s���r���x��v��֙Ȋ0\(�y��/g�����A��t؂;�.`.�1;~����a,��@��YN���0_r�T�yv�Zg/�|0`�]%�rą���x�efɜ��p�(&��qF����O�[���4��0�|cM�q3nA$\Xa���&�%�\o+=������K�g"V�b��*��OY��4|������f��Ǟ�H93��Di���]p!w�66mtqA�ˣL����S_��v��wbood�z��E�F�D5j#�������(s�s�5����-�$�E��F.�gܖ0��K���@3\ͬ|�n��ڊ���ψv�!}2+!��e(�E�%��R��OR�}�0�7ep�����5>����p褐MD�O���Aex�[M)u#�������7S,��Ǐ��Cb�M�x�U}�����"Ǔ�V�},0�o�����kh��9�a1�����3�~4yl��@ɧl>����U�Q�4o��x�1��P�T�����9([߀F"��|�8�O'��K��t�t\.~n�:��@�c��)��t�&�^��-�W*f���tb�Lo��
�ڗ'GN��j�Cx���)^�H��w��9�vXD���^2��K�V܋����%��Y�2�,��E�n�o�[����\���jL���3C�@��g���U	�J.+��b�)���^Z^�ӎ ��6����8��Ѧ<��!w��g�]�ޛ����9`�s�vJ[�J'3.�U�@4.f!#-���#�A~�5|���_���e���HP:w���.v�Q}�@�-�3����(d� �o��6�e��:���BiL66��M+�;�y��(d^�d�9��0��(u��_�LfR���+�K�)�@M·��kW�Ⱥ�M-�Sg�ݯ�g��$_:��G0���1�N��;흌_� a�����I�s�V0����aY�tL�|�cˋ9�@j�L�7�h��<�-�&� �4$Tw9:�J:�v�C�hsY��q4�e���7u�H�	ۋϑ��eʯ�|��?`��#?��H�(U�(�I֎A�����p�ũU�'��P=Oy��eI/<�a▻��*�-t�KxO�`$!���k���!f�g��X�������y[���UԬs�H_Y�]�Q���s?*�~;�ܪ����c5}6��u����l���B�͜���<_�E�)�$sG��?a_**�^�O����� ���̹/W!
��w�HA�v7)�{W�D�5M�8�Z#��A���z�%og�{mɁT������G���������.i���?����z.<4��y"� w�zz����Rk�.�j�Ч�t�
��m�~'HA͂�_�W�?P&�;��Z|�I� ?,}���c��.��������1���BE<q�"��(O����h�IOIn)��uQ��~�s�{�̚��i��[�(�ӏ�5�{�����?ֹf<���u�~kT^�����<����a$o[;�����@o���B�4��O�f�\�Jū�$��Ֆ�'@�ݨ})	�w�K�Y�Ѕ�jϼ������n]]�/^`�6.�_Df�����g����j�?�����T�?��6�D�{�K��j�+YE��7��&��ǱG�H}dќ"�rh�XP������(��Mk�76��(��c?�CRw�tD��۴��_��`]�:��`~�>V��,�E~Y 5n���V��G0oM뀸���Ӕ ��x��uDX���P�Q*��KjF2�%\��:J�|���&P��~ހ���g��,�-`��%�-3PX���a7��E�f�S�E��5Pq�7Ŋ�h�z�P���K.�4�����<�����3;Q@���ǹWK$a�@ꊒ=���a�<��R�������2&m/W�Ǳ��Ë� :����q|oz{d����w�s]*R���m���1����J�k �nqQ���&ֶS��:�wC�v^�y��Hن5�J��k�@�c��w&�5��sǿ{�Z���fW��R=m����K���S�dR�N5��,�?qg�Z����X�v�LW�W��+ٔ j�U�� �Ĉ�~c��ۇz�F��<Ҫz��f.�ht�C2(q ��rs��L��p�J"W]���Q�H[f��lZ�����;p8צ-J4.CB-���oE
��ޏ��C'�\Æ���\]t�H8�͌�N�`�k������?X����A���wӋ�H��%��F�?�`�����c�6
�4?�*�VQ{��p�V��xG`���s ��x yI)�����ɝ�51��iE�=^_�{���n�*��KZֿ�%0V��IM�q���v��x!~�V���7h|�C�
!�O���w�����l~�!n/{6mG��͋�=�C���� ����]j�1��r��Ŭ��j��VH�e*��mK�b�f	��I���	�<� �m�u��6څ�`���J �Kuv%8��bO�]�ރI�$��ڞ���6��������γ��j���\F�o�<J"6�B�� ���3���ӵ��<��k��N�}T�Dc�jS��_7q5tZVA�8i����
u��C���X��ʜ�{Iy���}ڵ�0�U��B���5�ٯ�d[��e��E"�9�٤�d�֢���x��0ww��Q���?������1^��G˫]�yom��0罩���a�|s�Wn�Hwv ���7�֚�^�t�H��7�-O�����g�1{���m杲W<n|i��`GQ�,�8��������.���(�)�{�6]��]�N�(�Y(=��c-C��c��a
0Ü��@W��<Ρ���w+�R�� �~�L4�Q������zޓ�Po]Q��8�頵٦��FSf��9����:T���G�@�-���O�h�D�d��	u�C��d�`} ��bH��S���2�,\S��Py��I�#Z��ݸ�*�1OHM�w���Y�o۸��g��H��XԿ�@�=.)w,���A�8�֗�O^��l��ý�<D`��x���h�1`n�3��!G��R*���9��c�
O�F<M��}ў	Z�ie�2]��o�[����e�#� �EU\�$W��r�2"$�}c(�p؂0ˤ�D�VJ�Gc��Gg��M��]L�A�g���٫6'Ry}k��:~�ݍo�%^N�Cf�4�lb��8�eڽ���h�àE�`�%�y�d���r�^YGH.�v�W��������Α$T������Z+���T,~&J��p�r���]�6g5�d_�7ë�u�(�>`1f�e"���
]����[}H��TO�%��rJSL�&�M>HB�������f��h[�.x8P��.�p���2�^�4JWM��	�?�k{����g�2�W�f[�I3~����j��3b��-q�=Ň�D����um%W��� @=�G,�t�q���yj�Hf �s,���;>�*L 8H��|��pʇ�'�����x���7�=�������"� /</i� ��kl.��R�@�@�ݶn�x B"vT�-kD�o�O�-�M=ǜv�e�"�ֺ0�{����8A{ֻ��`�Du��Ρt�J�U��3M�4Q�g�LJ�����&���Uќ�xEۤ�m1�I�������攐=�Nb�����D��z'� |#�h���[֢(�M2�stjӥ�z3V�:q ��Ñ|G3SA<S!�U��i�/+��_@�e2@�I�46�8.���v�L�\�VĢ֑�k'�<�i.ŏ���Zy6|��_Z��f��T���B�t�RS�0���&� W�����Od�
�7	�GwO� B������xW9�o��J����K�-��i^���`�3�������P��K��1�*�ET��K�rw�D�s~�]O�Z�V�DƵ.Ǥc�~��3�=z���CG��oC��Q5�8l[|�cѭ���� �� ��ѩ�v/#$�YN���é�fV$�<�%��b%/OV���'Lx���f��8n�=�42|'�@�J�� ��G�J�m�6<�x�f/��_�k^�'�D��p.L9��a�IuC�)?�;�jҶ]%����j�	��Z���0�պ;58ç&A�fͮ&Y��]�&��q�-}����I_&�Bp؝UG��Ep�9�����yH�
5C�IN���������gD���u˞�×{�<��	s�h�3�ޣt��]ft1�ˤC
�r7M/���4W໬{�#!EȈ�UC��6�3t�﫰N.{g&x�&�x��0���"I_>���AH
J"���5�<ܬ��)^�p>`ܟ����h A��9���x�F����*N~B��H
�!% u>��9_<��9�[�����[���C��e�:�K� ���F��o�/��X���	R/�3��z��`�`4�.��mU�Ctx�q�z���ğ�����*�Y�[�~}NTAĥ�lQW{q:U8��xa�ۆA��㟵�!h���&Q|������rN:� �&d�:*-�
��W�C��Ӈ��ƻ_,����F��9��ώ�c�h��+�eH[���>E��c�(A��G}�s�Wӗ�^��C�)�hS�(sJȟ��JL��V��>p�P@���E�R�^8��|Ő� |���k��9��NPqr1�Fd����b��Ǧĺ�Z-�@�_���f��h�ל#Rj}b\P��f��3��P%'~4���S_�����R��Q����%�NY��ei6A�8H��tМ�4��]�?��vU�0b��p�g����l.���n?��ֿ� ��q��[%�p��B*+�X�fP�J��V݅��1tg2��bβMY&ZxL�|�:s<��[i���TM�:o��U����q�5^t����fbn$�w�6Yvce�P�\I�\cD�����V�G	w�U��F���r�8������7eW��#�R:�Q�ͥ�i�k���"6p�hΝ~«UԮ�Gc:����И(&_�K�3�y�^���/Ss!<��C����)����7��Ax9>Q���Zx�y��&7\^)�Fo'�O�:���'|��@P(�� �Nܴ=��iy���B�&�T\���`��q-��n��pz�~�H�ʍ�@�쇕ݼT>������2�L���+�,
2{�l�w�^�!�E�7A�_x�h�_��.�<�1�ͤ�6ƨԫ��X�w�r�OPVZ���*�C��~k�u����|<�MX3Ҧ�-�����gu	{KM�m��R���\�-D��r ײ�ݖt��$&i�w>�R�YB������(�w�*�8�\,�V�"�y~kP8sKcb�)8����,��5��N�[VX�	,4�$�H��x�oG�j�ꀱڏ)}eK&�	)Z�DU�i1�3I��g}oC2��j�m(!��׽�QR%Z���2\T��s�W�k����r��jd�6�_���Jՙ� ��D��y���nk>�k��1,�I�T�y �G��LHZ)�晗�b�����`��Z�G�SA��T���N�S'1�����~/�
�-�2b���3����d���ί��rВ=Y�{�e��|<G��W��+�"xq�s�]���%>��T٥�X��>�YDy��S�\��� �fۀ�0fs�[/@D���D`���-�tc�a������# ;�/0$��� 	�kq�$w��8�x�}��)�HJ\Y�f���2r��g+����
�	�����[ͻ�P euE�ʱ���![�tK�@�̪�m�<�P��)��ٰR��V��(���ݔ��2?۶��Y㩃8�LR��M��0TQema����0s�!����DBKn9��0}��MU��b�A�X�s\�t�y�&�`��J:��M��7�3�k�CٔLd���&fU>�7*�?�����W��ş�|e�ta�h�	��;���"����Ć�S�h3 g��%���;��$��eB��}�"�QZm�u-��!CP��?h+��tM�ͦ	Z���T�A��n�d*���٬�֞F�-����äs�Y��jj_Y����O�ɽ���6	�z�2::�]U}����3���}�Z6�}|Ь2v�^��y�%9R2����}�bq�������d����Ls�w33�:�ۋBe��>~=��_��L ө�e���?9�ڝJP�+�_�Y�f����c����Y�74�[��V����r=�s�=�i��;,�X���WZq�����P���i���Th��+�
�����J�+h��.�|,�Q����USnq#C1��0�l��$i���l�̜O�P���Li&�ķeg�=�Rs��69E��P�w�3N�]�� 3tN��~���J&#�����8%����LW����9�`���%+GX!n�8�)��٪h��/���5���s!��f�}bVG�*Qқ��0������0��cQKґU��b��Q�LH�M[�u>�.�]O�K�${�D���`��q�$y?��͏O�-^޾�N-E�V�|�쪄5YI�Γ��=t3�u��W�}�4�5�i\���~��T��L�����][�V~s�J�ء���@^��| BC��|����޽)���e����+����j3���2���G�>~�^��{���w	���`���vY�}K�#�uc���  `~�1x��H'9�>f�P)7�d���U�c*z,==���L�v����J�M�X-������/�+v��p0Ag��f��ٲ����
ǀk��d~��7x�.ۘV7f��`덹%�mIFY��Mu�w|�,s!������"�����;Zd8,�]�n�k0�h�f׸a��3F�_���C���������`S0�b��J)��
@;��p?$e	Q�o�<�S�f8�k���䐛�۾�Ec���h1S,������ah=F��*�j��u���H�6�83W�p�R�4�#���`H�w�`tba�]`��!��%��V�-�u���ݛ&BO�ߪ�T����W{�V��r�� ���*hp\�~s2;�Q;���	�S�R���ɠp��	`���'�w�$M$��� ΃O��M#������q'͓(�b0�a5b_T���k��UZ�AHe���M�\&k!v #��(�Lڏ4���$1�kA���c���D�H1�Ƥ*5GΞ�5�% �+��ݗ�+���Ӹ(���UJ��C��i b�8�\K�\�T#$�7�4]l�L��Υ��ä�	�oM����?�UgBr�p;|��N��2˜i_w�u��7?���w���_�&�k4���O&r�����a�#�D9P�yX��H#y�ņ�!��%4��{3�~pt���ͦ�p��z� ��J������P���,���ǷO<N�	V1y|�w4ӌ��c�T7��XZ[�1}s�^]x�Jy��7���o`/�cVI�0�ת%4��Oŧ���
�ZaE;ߍC�D�,��d�
��9)\����)�[g��1k�|`�ҵ[nɑ��{�s��FU���ٰ�
��Ӹ��s=>-5�n(l,�R�%��B��TŨ��U7K�B���𖐎��J�	����d��E!�6H'̞��m�(�^����	{�y�ߍ� 5Rs��3�b�:�l�Ѐj�>�|?����w�ܱj��ݯ�kE�h������������9Ьb�'Ψ�=%�È���A�}+HM,n���(�ߜ�G�L:C�}�������]��tD���ʇ����$�\k�jS��ō�R�l.p/��x$E�u 7�sHP4���?RӞ�kN{�Xy�?�������Xϙ���=l�5Bv���PA��#��U���ȭ�c*����CW��R�y}�#�Ke۶ʈ=�[]�r\lA=b�����I�S�@P�6��X�	 ����е��LG���,�>���D�X�� ���j�h+�gZ��m�j�i���^��n^��3�4d1�.�~RW��
��.W�P�;�=���b-X��z�d���!��c��̡>bx���_b.ڲ+�]���p�^�ྉ��nս{����J|(��g(��G��`��>U�+�R�������E��I����(�q�E�y�F�<ր���
0��FL�����z=D�2"��1�E�$�'���gjh�}s1|��B+
2�G|�9������E�t[��S�u]���.��h|���}*��AN�p
=���#���"<�����������%�dBO���sj��v��]b7��k
=��$IN��m�&�;��TM.:^3��D� X��f�tT��1�(��w2:�ȼ9�$�8!�^T�:�n��<>�=�Eg��֨�%eJ���lI&2=-P�TxȇB}TWea+��L7pHp�8G� Y���4R��j����'g>a�eL�ᚺ�Z��dJ9���^��������9H���?�2xZ�[��Oӓ����l=����=�v<��'����9o��*�:�/�5f��' m��_���^���=q��2F��m���o�>r�>l�EEw�
�*�v�����_�H�!�;���@�¢X��wŲ������Ǹ�}c���;�~J��p�W�����a��"V�Y-K2�s.]w��q�9~q����ދ���j��_�63Ӊ'Vj���O�,��l��~���,عV]w�ӏ�����#P$k	�!����sQ�Sp��!{^�e����=IH��h�����e}��T��8GR W�y�0k����rl$����) �G���F�wwK��J2���z�'�_̴�m��7���.4�L�K8*�R�$�۠o����-��p���]j_e�xv ���t��	�5Gp���Z3���������­�i���l�:������'��,��"��"T�S�75EQ�O����F7��AYX%~M����#�	���Z��M=�ɵfY�]���1�B]2�o?.����:''������cZ�V`��x4sHR��Y'T��ў�T� ���A"a�nrԗ9��ŏh��%-���-�M!��j%�C6���M��}K�˛���̒9�
}������ّM檀���,����|}�Y����� Z���h��q(m�B� ��$e���\��1�~��7Lz�ۼrٱI+�ԯ�����$P�7*�6O��w3)[Y�����\*͢���󉒣��I��)�I�4`��ۮ[$�u�MQvG����W���r���@��n舄uԾ�Ef͎�N4����ʝ�G�=�1V
sh����Z"D푩�Z�G����賶f\��hB�L�¢N2ϦZ�9ZO�P
��twM�ä��#��fI�,S��Q_7x,���!�e����{, �PF��fz�F>+��l����q�$Ј�׮2���X��\�S�dQޥ6*�����#e��}ތt�>�����g��4ОJ`�D����ஸ���힪��	���U�t�+E}|u|_Z^Z�1'}�9/Q� �U���QgMOS��9�|Yr\yD��}�����{������d@���z��·Gh��� a(��i������Z��>ػU�p`�}cQ����	A���-�۪�L�DG���H����N�����asx���?���=�ڥ_�4D�T,�!�3��d���d1o��*J�zZz�i�e�[*WW�R,�-{dq���8(=�*"+7����Ekڦr�7n�>�y�w����{����|&�ȯB��&|#L2�8�R�����+�]��:d�}�+|1�;$���p��+��̹�J��Y�²��>��G��j<�dR��1=��޼��{�l��`�(@"�OI�Q��g@hU�O�4�j�9�f!�~���uA�'ga�;Y`�������)�	Gi��閊�����),��=yx�{8|є������t%9(��jA^�W�yfĩLz�py'���K'��/�i� �OXK'���FNv+ONd�����j+e���]$�=�=����H�8Cn�o�Lk$R֢���j�5fC|�#Q��%�o��o� .U�7,|'�|��_�pZļ7�3�s4匜�K}z����S�a~��؂M��ҳM ?>�I�x���klX�c�~�3=١��(��z֯��s��2��V��R;��@Z�.,�rg�F��ct|�C��&�6�k����C�``{�e��Jl�]䢼|mi�Fԥm)D] ���.�3���W��%�F�"۽��G|쩘�w��N�=m�nmᝳ^?�]��Ere�����g��BWN�3�;#����gR	`�q�>�!��2O:�W��\0��*OW�Jt����S�0R|��'�E�!v � X6J�s�I��4 }���*$�����*0?�!���M%�7G2�_ԋ(� ���ܑ�Xβ�FʱEhYw[T��E����W�+E*[�18S�s[H���f�c�P��v������m���n���
�k�[����9?�3��+G��"�U�ۂA ������PE���? �E�8�p(��k���T�7����>t{m��D���|ϧ���k�@}�- �\�:s����$�{;
��/����~�F�V:DR�'<S�b�3�%^o���d�>S�w���>}�:y���bT�{JLɌm�Jj�;�XWA�<�?���]F��}�`�={6�lJV>ݝ���'�M�V�C��^��Y�2��fK�(	n�i�NlT��� E������O�f�*��7�7�_iO0��y#)�o(Z�ʟ�E	3�$(�9Ȭs���c����}��͙��4����l�e2�D�U�nq�#��_��6d0>4���Pĕ`I��eM ��� 	x����w+�O�{���JR0�����Xx2�,g��f`��)����V��N0B��I�rQ��f >��+R�5s� ��x����)��@-��t�Kx�xd~���h�ԩ�����X���:�1�f�����y��X��g�d�S�ب 'j�Hm�LVV|lIޫ��%��W�����M�C鸨zd `���5�p�E�7h�J���N�|�H�� u�zs���g�(�%�J_�����T{&�����[�zou �g����Q��*��}+��0ӣ��8;�,�K�e�%zE�N����ߒ�����6��/o��-�Y�M�����|�=G?f�u�ds�y-K��1[U�D{�ã?;Ou�/h[� ��绣�E<Ś���:!�&EP����h�:C↷�Lh��
LU(ʹ��ᡞ��䥭sF�$�+�쩴��i\ ���p:8��4̴�}��&��Z;u�>F�������S�Y��z�T3��&����,�H��	шQ�Ū:#J��#-Ȕz{$�7��u���» � ������5���Z]���+�K.
Jπ����o���)�Lˋ��S��w��;����o}MV�]V�wq��K�Bz���M�:��A��Td�D�����m��vUZ����gHq_&6AF�r�i���['&Ŷ;,���xF��Ғ2�L��-��� ���X�h��V�_/A�SJ��+��K��ޱ�L?RG`y�0��	F �.,e.����o]���7���$�P�X( �Λ�*�p�.�K��Hi�
�gd�%�����V���9b�o��]���8�B���6�c���9*�^���n�[�o��cUϨ����
m��/�,n����&L6�S5��M���ƙ��+ l$I��j:��\j�9]�]��9h��w����^7<�FQ�^�s�:�S�f�zr�k���=�T^����.J�?ƥ�"�xn���|�s�v<�`�:Tu�;��Jl�#9� �N�
��Z��ǘ�w����	�n^e�� 
}�=ڭ;���̕��`E����xlC�=�u�G� t��|�A58���A�
��~aq2\.4�d�?�i�9Y�uvY"���u�8Nߘ�F���i��ըڻcjʖ�|�p k�}�Ρ��q���_����aa8�ͪ��{�ސ.�}d, ܫ#���E!�h�MV�������ftke�k,Ë���e\�F��C�tF[5#��==�s��5^'"?_JڞoD�M
�º(�\�+~���Y���u1��ȷ���j���	u�qM�ȡ��a�ȟ"(A�j�-D�G�����߻�q�h�+�J��sbds��䮅����	�nd$G�76+�[=X���`�u8^��ė����犲�W�ZAd�[a��0��p�0�� ���L��+5��1��<�RĹ@�bq���QA9��摴\��n�=.�q@?�WP]h\�
N��9���eG
.�����	�U@�s��9����f�'�`������dv�i�Z�N���2�C���2iY-:m�a�,牒I�(Ag���?̢u'���Y�I?��EA�_��TԔ��0���.`���	C�!h��A�8�ۘ�t'EԠbT2��X��^;"1\Y��.��ĭ��u�vv�sP�$��K8�>LØi���G����~�j]�DG�%���;vN蠉!�ǝhr�O�\����6�;���������!Ȥ�ŃN����t�٤i8�X"�;J�(�jul4č�+l�%�;���>@i$�ے���fq%R�0�X���A��!��8�D=��K�ޑǅ�����O؈?���:�Ъ؄$'���o�];`l���έ��u�1&��P67N����үOR���'7�� Dz�[��%v&*�'�%����1�6[�ѽ�A�u�f3Ƹ���d��)���L���Z<%��yN��)6�+Q�UN��U��x�u�V��_����P�S�0�>�h�Sx2v�X,'�kg��OS��]0�b���@���%�j��I�'��J� �+
i͙s�1�s�	�X�+���š S���u>�\^|+�R�PET-P�iH ��|9��[�*�fZ�9������	�!�j�X0��l`s�!r�����s��B�lY�W�t�x\���9�c�&��/�?�ࢧpi�3.��?<1ϫ�H�5r��
���)40��1��$�U�"�8`�>|�	�7]tE�q�;%bLb���@	��:�갺A��*�0vn���_��?�	�J(M����zk���k�O��{� &�)���4���$+P�W=o��K�e��\����Jd@�։+
8`8�	H^z�DԍR�U
Q9�~���7�M^��s�)~kٺ�;�*BO`�@�E�����
�$�ȌR�����RGV{ �b���P�0UL�(<��W'�>��2Y�T�����a`�T��E] F������Ѭ�T@���n���=��٥$R��Z�Y�0K���A;�Hم��Ѭ�%3�D}��DYW�Z6�B��U�j~%��4W��!�#�v���D�q"�P)�Lw��'���#�O,n-���jC=��V1M�Ѐ�x�h.sv�=�(�/�}���y��d�'�2o;'Ƨa�3���!��I�P�3�;T��48����r��cю��5iZ�֓hk�ij�� i#�^A�l}��}�Y>,6FG�|�m���	J�艢�����`�����t�Z�2!��_ �ĩ(\-j<;ٞ��H�^�e<4 �����u�0���T��&�v�1z@I�0H6O�Ӛ���u� 1�/��f<ƾHqgpZ��3fn7}X�k�@��@Z��ގx�k*Dzc���%�Ym���39�J��G]�U#>�+&��d!-�1Pyd��=ɡ�Zy�n��G��ɚE���ٖHvd��~��ċZ�ݼ�Me�J�����Zz�dC	�i��`��A������?��z�V��ݹk���z'bjXy�D?�1�ҟ>�&\\� �"��/ >a=����D��$g@RnU��1�Ǯ�m���\���B�g��b�*�4�$X��X%�h6Z
�@4����Ԛ�
�l���E��͆*�֥�zø=�ru֮;�c�Ak	[���j�y0)�~�� ��S4+��^�ݑ����$��@眑����(����(3�KB���+ܴ@�,�f�������QJ�N[�FV�w�^&�p)N�(di�s�Ϲ�"r/�ά.@a��I�
���\�%�[���/�s�0����H�䉝�r�������M�$�U�e1O��ne��NFn2K��"(�"?�\��6��B������gL�mjĜf�pi� *��q1�8����Ka��D�?�ئ ��ǉl$�i�A��+��/Ųk����MxK L���(Fت<;�dP����1�b�8,�̜�[��%gl�>����t"�3���9�5�����f~E��S�Z�sh��#~��*���H.�<+:ݨBs��¶F_Pr��v[�ӻ�M��2���sʹ��U� �-a/��%3j��B#,q��S�e�S�g�6S �`���V6��_��F~���zeೝ�Ϟ�vGǸf\u�:7�c��&�My�i�maCH��pl������R֥l񋹢e��J%[3	qӦPj�+Vk���D���{�ζ��TGڭl-@c��y��*�X^.PJ�^��
:��J]
�I���tۦ3%�V%Ģ�����aozӲNTP#���'|Ў!6��͒}��1�R�$}ȭ7���i��� , k^\Y�K�J��(��ҥ'GST{����k�8x�O�� K�� ��x�ףz�|�*Ŏ$SF䢕やJI���k��D��� �=�uɗN�[^'i�k�J�[~̢��#w#F�T�2��>�Sxc����\V�m���XLeR8�H ?K�	c�}{�~J����.�X*���l<������`�[����w�Y�L5'kۉ�PW��q�������Oh~Q�P�F"3o(�tI��A��Q�[t���uܙ�p�YQ��'B]�y0v�¥D#���Ⱦ���t$"��9j�,�ѡ�K+��k9�,�)|At�7����U�6���`��C���W��V�OrVZD[0A�ˋ���kY�@�PI�	�|~`̿:�p�H�թב���?��⇔���$R�^}����IТ��0�����+�O#1?d9,xp�X�jK���x�'5�b���v��/'_ۃ}p�Dd^7���n�$�� o�n�y͓Us�>�CQ�M�Z�	�C5�_T�������E��UQ�=
~fΛ�6�J�跌+;��t釙�'b8�#�����"�'��Y�,{�����9s��������'������Pu�"���Ut�?#�tr����Ш��,�%v���Y�mX:t!/[�P�h��
�������zub�A\�g�{h4���#�Z��o�3�.������mV����,k��8=�(&��Z刎%��4q��������㉁��9�L�9zC��N��.q�l��3.z�R��Sz��`4_�k��$�n�"�,TXLV�"R7�c�r��ȓ��C�k � �VķXH�(*X�	"�+����qbP�U�`H+|An�O���*1����5&p���U	���55C�"<�M�SN)=��2��9��rd��`@��Z�v����$	&{�\B��Ȫ��R@����u=$7(�0���	u��#�b�]�����uI�q��8k���}^�*�j���Z�B
"�5*i˜\���0�c1�9�(6c����lV�ў �OBKDrO����%�#��\'Z'V�?>p���������&�B��O۫������ӗ36B����$�-��+�}��/�`";U��mҟ�t���E�BS	E`��]�D����|}D������a� ������Hr��^8SE��(عx�o�B�����R���7��k/�H���(+,6�:ܱ�L��X��` ��;����$�/�L��B*��?�5������.��
3ω	ċK7���K���ץ��M`��1�"�M���Dd�D�e�Eb��ZA"Db�t��V[m��� H7�8�O��;��_��<��%�ύ@{J�D5�w�a��u�]�un�/ɾ�գc:AY��~шG@���f6�3� je�E%If�����q}C���|�y؇pޟ��qY�4��ah��[��%����#F�Ph5��:�;�#��hp[�������ak'��
A��8ï��!e~q.F�;��MA�@���frq�K�Sw��|�g
|5�;��t�0�F�J:����Q:���E��!U�{�b6���5ܑu-e֜z�v���K}o��>��d�$�S���&�+��(��9�$�?-s|ygTX��!6  �[�Mb�N	�K^��	,���x+�[�c��apt\¼�4������%ә��A[�����g�T��_Ha���B��St��\O�8�>��'f�S9���i���(׷����M�;�G��M#����q�Z���z莛��l��3��HkT�s��G���|��{|�hQo�r�?�#^d��:�j%�7�uǖ�ٴ�̰��=X!�t:j$�1��4>�)y�Fx6����F1YJ�Q�ܷur�� 
&i�(����<��Hu� ؔr��]F����;��^���GǞ���B���:���B⧡F���:-���K�W7�~��I:w�v���Nk_��9�U����}�l�_u��`� (�"N7q<�Wq��޿Hc=�7�4zo�Q�k`%��\��D� P��^iR�s}�x�[os,��k��O��A�⁽�z�|F�j��]�r��~��X��yY�f^�kgcpc&+t]��@�z�l+�����S�I8�w2, X��>�������z쁺ۃnJ���"��V?-�9�~��Qa�]���:�t]G]L�'����OhEH�*�qjKv���ں�Bx"+����0�Ml���p�)fg����汾����׎K̥l�s%+&Q�M�"d�:�ޣ,%�����O���>*�|)���U':�^�1dEnΆ2~f��_G<�eu��y%���I�H�g���E�,>��8Fr̞24���3�˵Rx� ���8���l�Ea��>¹��vfb{�bNq�|����3��fXn v�QQ��Iq���;�0m��lV]�m�zL�&B�P�[e~S���`���t�t�{�N<=�j*w[7��qDt�e��U�������%���<�r����4��L�Ξ�]@ž�����L_pl�3��c�Щ�a� â����$���O�]|X�#�J$�iƋ���,͕��� nh�����4�D"h�1w<��
O
�P������Ӽ	_	�j�qʭqk޶G?��5S���q:���?�[9QWъD��Y{��q�.}ޅȶ�D��ɠ@\��(d�2���T- �&;t�r9�{�Js�6�O��8Z���u��͙�	�Lo=맄�HRu�B�N��iS��yF��l�����j����}�bu��EC��W�ϏU��t�FV J����"�;Zx��P��KwśB�y�`�����e(����龪b��w�u%0Q�<�m�A%t�?���^���ݻ�]VJ3�E
WՄ����^/�	H -n�p.��ri�Fl�9%�E���ZɍPvt�%&�����11C���Nt�����ѹww�"�Uj�)<��*����Dͤ�>+���||ڃ�a�spt��>�#�X ���*nچ�.r��|�������[E-V���;-NO�s �s(�.��W��.�v�<�&��s��J��hѺ[�a�p�C��\�\�. N���u�^��7Xt�J���k==�LI�
��+�m�]lɩ�RE�5�/5v�5e�E���6B�+���:�r%�4�ބ�����q���k���g�F���5�9�gxZK��~�J�Ŕ"O���H��ǽ0v{e�C�&c�P4���A��.���w����I��m���?��9�m�޻+�@�'H��`�K��7���O��L ��ؑ�� ��]ա��``J[�Ol��v�c��G�S�R�Gkio�G�Rw��)<#,/�F�(D8ag�&g�9'R��B�O�(����4�r��$P@�:5���Jv�'������ Q��ґ�h�;�x�|�'"�'*f:k�m���-7H���l���~���E�U�Zs�G�����ݘ�>���u6=��+Ev���N8�8�;P�&L�<�+Z���0�$�Yq��X�>��._Tc��;:���Nx��Oą/��!���Ф�7��Tl|�{��/ǬO͕��2�)>{g���n�=^o���q�#۶�'�x�\���E�v�"0�3
w�z�Z]�,}����#/�iQ�/ 4�;#�L��O�|�h�X��Q�V��F~T�����$�k=��(9Ri5���|�L�X	���e�eٯ�e�a(s��F�^�)1��-��E�<��@�pX�a�V����ᠧ�RN�ǘ*H�F#���{hvG:1ٜ�1�<d�!D1א�'S��:� �~��%b���<�u��(�9ej\Ё�oy8q#�;Ht�*�C,���w��ܾx�7Ke'��}w#�m2F���&i!�,����3�4�r�,�/�x�ĥ�O7�*�cuX��#�6���^���ad8s]���1?�.�I{�������V��n��a�o�T�9�+�0�,`ٸ<�av�"II�" A ֽ�0'��#��<���CJ��JA�,ZX���;yK���E����?V$-��f&�G�7L� ��D�����;�5���mL�m�(�9v��b��֪��;+����;+Hd�z�,��#�="�����W�{��P�l�ÍF�=�n3�!�Z�@+��J�w"ؾD�_��ܷFD3�
qU��I4�� [�vaZfX�
�=GH�e�/^܋��$U6Ri���|D:��<�Ǻ��zR'��zSVP������ӈ
SS�yk�L�lq"D*�圐1�T���ʖr��sz����?*�9���MN��x��;�{����.��B��/�� ��2�v�t�*	���~v�����_ٍ������,x;4]$�}�B�����!I�;�����a���,؀��d�PXE"�k�l�L�{�g���r���T�j}����W`�O���$M[f�Fi��c��T)y�I_�+N÷;:�^�TvB���Kn�ΉV�����`���x|h
�䞮1��;t��x��o+�G5�qA���S���n\��&D��\O�׃�8��8ܟ�l5&��x(M��ˣ���K�B>�HZaLxH�o^m���S��x�� �S�Xͷk`�=7����u:ڝcdd�T8c��^�ya~��P��s���ݧ+�G��iH��0�z�2�0p22��z?|p�n�s�O�F֛ұ��B
�42��|M��h��۽-袛'v�{!C�X\)@��ذ�a����}f�PH���v�~g�b��t���{�9�Nd蛢m���!P���LԐ���<~Z�~s#�.�7 ��C�U<�Cޫ�c�ޘ�/@��[X >��~�����?M�lN�㝽HMgK��D�	T
,�S�����9� ��m=.1�}F0��\�ulC����ŏeJ%��\΅�"6�=���v��*?*��Y����7Q�P��&�����,E��0�F=w#;���w0��G��]�G!섮]�ЮX"$OT�t�;`~���6�Y��3���I-v`�{s7��,���ч����0w`n!�b����^���/ <��B���7��J������$��̛���*������DH���[O�kl�~Y���'�$P�d�Y3��?"�]5g���1��BG�\_gJP�1�<9��u);y�YG���8߮���/���ý1p�`�9�hp%�lHHt�Ah��=�L5K�#�g���/�[�ۼ�p�7a6]__�(����PDGu�+����;��c�z%y�1�yJ�\������5�A���>^��W��U�%�_5�d�aM��`d u�Cgx(�j�M������K����C�ˁ��i���e�z�[�h��r�/zn~�i��Y�b_[_n&��J�t���3�9����O������u8�
5���P��L�!<s��^���a)2*�4�vex�4�Q�afz��s��nU!r)�� ��Fnr�li���ߺ��K��͋���-�U�p34N�@�A4q��(����8-����6�����T��ZH�Q�N���������X� 7"�_���֣G�����ۤu��	c��	�v�����{^���۵"I`Dy�ymYV%�o� D�����f��)��I�	z����'��	;Q�$հ�4��[OJ��<_�څ&���{�FL�|mPB�dy��b*C�m U[�S�Z���n���D��8{M��]�:!�y���(�"��-z���Zu��?�����B�<Z�i�:σ������`��[�Y�6t.�K��SQ^�V͝���8�>ȥA��[ĉ�2�B�lQ8҆����lM赆�t�#h��/�c8��R(DJ���,�l�4������9~(�Q#'n��h��}-G��*2����g{DXv���^ŉ\�8>H�w�K�~7��D1u
o}� j'���������ዦ}�̧dK�N���BKh�9e��k�/NO2!��P`g���6�ݐ��]a�����#�v�?����/N뤕�O�,���&�2/C�����'L�'{�>g�j��N���;^~�Kc�՝���Jw�w��ĩÍ�����h�G_���~����c����R4*���ץ��ê��;K%�<@8���U� xT]�=����7���;$h:*	sgo2�e�$Z�s`�%���(�W^�&�)ROLO�Ja+�2 ���-�\��/���E�7�1b�������H��o	/`g[�$�} �l�?��e��&GH+�8���{�g��MN�.��q@7���I��t����o���9���3�����y���Ԁ��Q������2�P%-Q��Ş]�/�0�rP������M"$���TE�5�z۰����<�����^;ĝ����Ga�y7N�׸Q#8tΡ�����b4�M��j��Y�����޷_k�:	���p�)Q<o��l��������)\1���}3h(�b>E�F��ITg����-s���n!&��*td�{��Lǧ�S���=�+*6K�$���tM8�غ�����>d�?�f��	i؄}CS��������,�JI%8ظw�rqڠ��j����Y��p���w�Y���K�X��OrG&iB&�(_yd?0�D�l�J_����o�n=3F�u;�+P��o(R�{�(��q+��W���e�UKmj���X�4Ì�p�n���6�#��m
7h�� 4�Ci/�4nvҴ��c��n����aT5S���_��CK�|���"r��4^����?ک^0S���B�3OA�Im:��@� &aʪ;�������e	��imy�QF="��9ʋiS�IZ���|��L�%�~BQ��p�&��:�$츆�����'�5 �)Ε@���Dz>�C�#��ןx�z7}�{(��L4�_�Č[P�Kǖ�R��V]�k�=Xd��}v^~~��-FnQh�u���g8��\-��ߑȜ>�)�����C,�|Q�OD�~����6v�w��X�.bYɇs�	r&>�0��������K��p{�]�F����@*������C�D7$�:�へ���:�ד��g�c���T�#�G�Y�y��]�-V�`Ӛ���)H-�2I��~U���cXY-� ��
kJ���d���.�Ƚ�U��%�aUc
�z$)���J�:���� 9"�v�H yŸm����=X5Tf���V60�c��Q�g��ZGV$-���j���~��4��a)�e�cG���Ɣ�^A8��(?�����\�I��:륫�����:c��`3��<��ʼ�\�8EX!�s"�eܳ�c�e̊p�E��&x�"d��_�.z��kŕls�X盀�����ވ�%�v!RjeACP.>��oOS�����xT#.�j�^C`W�l=M^��H' ��a��.h����+~��DLb�q`/���G)�l:9	��ԥ�ECs��bs��ŶE`b���x)�j�8��f~R|	uf�Ep9"z#Fx���V��6�Vmf�L�-|o�V滩v?tvzƭrsuX���C�;/��Il����6"�u����ld̚�w�G�	<��e{���&��;�h�R���k;�6��y�Sw �]�;j%��u�.4
�L�_uِ�l$�j�9�8`�xr�	t�3s�W7뿩/w��j��'B�ؗc��սUq�xKe/_�OSt�W`iU8���%��x��m���FV ����ty��,J��Tpي��Z�O�� ��~�/$�qچҏ	E�[����~�*ے�������[�-?F���l�f�R:��6�$W�գh8���K�[N^�k�.���@Y�K9[�E�'1V���p@K�A��2�j�?"P;C�9��|9��x���oj�x�?�|�� R�п$U�f�DAf�.n����rF�����}��È:���Dw]�l�)IMSs2������ְ�E^�t�@)2"����8�]�)Gy�USar�79*��e���Q�y��� .�_�]E�4��=xJ���6�
FdQZ-���� ��lq�tk��GD%2�Y�D=�
�l}D}g�m�WK���q
aե���n� �E\�q��\�<� m�T������#�6)�9y7��r������8���}�s;�%�g�8j�]`���n�A�mA� B%��{��
[S�F/��[@��ũ?T���� �KRY���L��Ҍ-�Wo��N�("'ɨ ��f�pO
Ju3+}��'SZd��ᰱxW�{�r�\L��g�Ϊ���8\=D�B4Q�}�3�<�q��vƤ��T���|txn�l�y��S�<@��-'V��Ӏ���<��̳*��x�:p�!v t�)���������{�v#�|~����M��uhD��3��\i�ke�Bvc�bV�*		=�ޫ�U�|�&��}��[A���&���0 �H��u!�9����	����~�|`+@�Z������2MO\����cޡ����D��	�z�z�#�
�_��9+%g������n��\��Mjڰ����*�?��4͇�OH�hX²��>�Q�)f�>l�E(��1�)�����ڌ!2 �lZۧ2�0Da"����>�
t�儭	�A
�H�յ/t>���6'��>;o�|ɝ��-T�I	�N�Y�-�w�{��_L�[��r�uQ��|�L_V�ْF�'zJ����������YM�k��6\8���S��
YaO��v�?�@��`�yԐ<}-��i
�M�K�#&+���и���R��>���G�aؘS�Wa����X�5��yg���P�ۢ�E�Č���}D���nd�a�txDFgI�^W_�}�u��>�oj�q��=DI�B�^wJb	w(�Q �AF�!�
Bw��1�g\�wE����U����;�u�sc�����/�J	���c�3Ĭ�H�+�󖗼��@��~헁`dm�>G��� �D�X�_������Q� �-q�9������::a���b(6��U��a�T�Ϧ���6qq��;Rڿ1���1�<lj�����|F�N�a�^���7���<*;F��&���ar1F�tuOzR�k|��Z_#���cHH(��+�I{��.u��Kr=��,����H��x�!�j5�(Ƨ'����;�Ji�l+�Ȱ��ӅO�c�:��Okd�'��p�&����w�!^�[ !=�����/_N}��I��<����pa�yX���giEp��*rQ\�	V�Fq����[]5p��1�r;�{ �>a
���|S�ʅQ_���^��iAA�D1v6%	�/�x�d?0��|a^}%�8� ?P
�8ku����tÂ�����w�1Q4��X�ӆn>V��*��"�%3������˛8���A�����z�5��pZR�dJ�w"�$l��?����/��W�r�rtI�!|��V�#f�g����Йa�g/�g�c�/���>)oWc��`h�\�wB�ZE�Kj��{�l�?����~I�p���~h'�W�a�
�F�=����F����	Z��,Iw-�ӄ�4]��&��ZĤ��N�1>���U������i��f(x#U��tt�IY��|W��3�R��ؒ����4��"����PS]?+ğ�K�����n�(F]�-wu�t����5�G�d�7K:q�q������(a1Q��Ԯ�R/� F�$3��^'Ά����N�$�=3XϾI�{�~(�a�3U.�,F�d)��]�'���g�_B�G��Ũ��&�������w�=�0���Ng��ʇgϔS��#��aUv��(-�I[�u�y.����J#��������#���}��q 8s����;#vz���{v�Ү�"R"������ʎdl��:���<b�׬U��>u�?�󡆑cJ@��}�q�ap��6i|�&��� 2���C��6y�l��#��sɉw��=sEJHv�;���s�K�������$o�$��澻��.H�������ڣfv:_SS-)m�W��ٔYl���r����%v_ �����{�~��/�)',ʓ��LX��NL^r���h!��)�f���{цi�5��@��8!��D��x�!�F�A���uz�'p�OQ�و!��T�Ԕ�.��L+��Қ��|�}(���e���\��$�!g9��6����L ���7��.y8�V3 b�E�y̑�{�:�+g�0���R�����X&w'6��nso�t�.R�$Nr�*�%����1�rK�]*'�[ЛE�ˮ����D!b��2Fu}P}�5\7��i�}���$�-@��x�p95r�.ٲ	��<��Ԙ�,��[a���-����,S��{F'�->g ���Z��:����.J!q���������t�da0������g��+���⡓��/k��F�ܜ)]�*}�ˎ
suyݴ���^g؈�;��A�;�9F縫��I�Cu>�ym�G�'�CW>gEn��Dd��?����f��/��`R��:�K��oq���,�/�R%���n���[o�a�V,���qI�T������� ���j������o�Ko�k�V��	���U7�0�I�ʲ����gO���;>�ƉD��;z��J��6���7��3��k��e	)��*�y��D}`��T1��IZy%x���$���q��uܩ�d�ݼf{�w��Z��eN�����s��<��4����{u�`��r(kv�%f��Z�G#	�O����?��pq�LԩqY�Y��I/�/��]�#�6�\QbB<ڀ_� ���ڦ�>��,�����"x�!>�za�RŁ����,�Oj��T�N�S5�VbI��U�\��ñ�A�(<?J��I��+4�gX�I����7 � ���&���*5�U/�|�,�mvsڞ�S��{a|`���>дH+�� ��ڶs��zV�-�z�W���w�O���+��Z��S�NI$3��j-�����o�3+�t������(���y5 �xo�v�婝���M������|�����n�"��3x���K�p{��8.gzVm��>��%i�t?f_IHM'�6��qu��S,��g����XyI�y%}{c����~]9���rX� @6�%�iޟx��8h�C�<_�ITQ�mt����[h�K�E~>��"&�ׅ�x�E^19s�{��8�8J+�L�s������-Y��ѐ�.�(M�Q(qb�x9�X��%����|?&W�0~��G������p�nM,߳C^+Qɱ�"v"�6]?����V8����P�ms\�ۍԴ� ����� ���e�.����y��MV�x}��|�٭H��F�
��>:�����K�Ć޲0�����ʄ�Ә��!�H2m�J�ƻƴ|�m��IJ�����uȗ_D�G��<��!08�+�7�r
��^�!h!�06��>z�Bh\{��^�xE�r�bd8K�c�,���~*�T�"dXՁ�,� �P!8g��eBE�Zf_4&G��1��0�u�w�
$G>��δPU�Ӝ�|]c�#��\��e4)$�M
/�+�d�ȸ��_���B�#�a��Gd����˪�_�h����Y�N󤑔���u@B��:��{����η�D��(�Wf�+�-V��s��f=��`�K��v��[�sQ\bG���. G�aC�1�k�g��'��~��&ݨ��$��6$9jf8K�Gu[[�->��{(a�4�_�1	�m �|�Bb�EwDt8��M���W����PS�mK<�BW�1ǹ� ��J�}E�G��g=� ��S�X�H�y��C�&F���dB!�E��k� ��JL����5����,F%D�)���\�Nj��h�=��?~q&ͤ����g��\��::ry(9O7D q~:�F�ET�2۫?�(�aA:-��PL���	�^�/(��+,{.'�ĕ�h;�wg��Bb��>;�}:�����ȳ��r�[M�T��l��X�˛l����Y/����y��=�%
����"birJ0��U�AJ-+��}��HR���5�}5�ho�A�V/����ɠT�βS��$�얚2�3���'.h���D�*N7���
Qf�߱���bGm�Ƿ�v�`^J]��Uv�w� l�U�,�xU���%�[t�#h� Ʌ��@{�m[ߤW�֔��Dز� �"���x^��?�	Y>C��9�i�F�8��u�����4���,���R�f�.J�0�h0��Zw:\R�:��{-�=��oNⶍ�[5o4��c���9�S�q����e���M�����[�8Y���������<e�Jn��AFz���ow�P6������xBhD'�{Y+S
4O��o��V
�(�I�1?�kAQ�rk��K���1�9U�?J&:�?š��$����q��������.���K���K�/j`�(nK����,uJu�v�m�{>2s���k�ަ6����>�ݛ�+�)��\�ͧ*�c�F6���Ā�?��ۭ��ny>��4�6~��F9�P^�?�z�u�G�it�ޟWLa;Lnb���/Z�w#X�x�4��}�)e@_7��G���b��j=�t��]~$cf����/��0�ʫw��y��`�ܥz��:剙�8;��J�}=���=-�<ˏ����L���`+�|� +g��VK>ɵ�ڋ�����4W���Jw���E�,�Iv)�V�6Ԗ3~��Ɠ�h�V����� 0��V	�h�=Ip���g���>���s�P}��v���3�׉�AE;���*2�o��E��4�j/"�� �!PJ8(#=���7C����6!!{Б������I�������m�����vU�l�ӷA�F��$`�o<0j����mh��;�U|�Sc��дD�tݷ�>ǒ^�/+��;!d(�M�N�0y
�R���"V/�K� ��K�3A�81J���.��U�Z
�R�A���K��>L��a�Y+~4JD�Ee�����՞�RiWE�L��_:6%�y���:��P�U>�HTI�v߲�R`��c��/ڮh���~4�����F��[�������E��˯_5�f�^�$�ѵ
RzN��@�k��@X����l�if�[�ާ��[h_��/5J'^y�X�$���!��jVi`F6�����y�#� ؎p���&"���ԩ��שܓ�|��g�`�r������-��ǀ�� }ҖP���?�yǗ
���w�o����F).��զ�p�	x�խY����rd�+h���(����Y���o�:��f�{�\�K��B �;�Ή��y�ߗdz�Ԛ�{��7��.y�}�����	��27��|p��Z^SWN�c:�pv��ŝ���
���F���8�P��z���
;PǢ�e��& l�������W��4��Y������)@�:�1����6�3�����Z�$��r�7�E*�s��;���|�ֶ�2�lkT�o�*������pC99G�]	Z_�f����^!����d�������ɨ�^�,�Ҳ�]/CK4��՞V��w�Zp���J����?�B7�`���Bɑ<����,�vz�a�R���N�}]p����Re��Q
$}q�t��B%Uf6_��Ѥ��Ƈ��ڈLR�HX�hY�Cވh#���
.�����#�������!!�����u��i�r��$"'L���~�!�Nx��ކz�M~�H�=�	�CK��<���]!���G��g�ct�u�V��V���4�⦳��uh��_ Y,���ى��2K=�Hb�-�,N�o�OF��,g_%e�.�3�]2V�1 83M0SU��tbe
��V2!�jY"^���x�9
�ħ�˷P.b��5�q1���3`�S�:��K( >ד��֔&ֿm���&����pxP��o�z���q4��#Zt��>|��2��xc��HI���M����'���i	��>�%�A��(Pg\�сRO�o���� ��n�5�C��17H)�����fgu�T�#�X�]��������\+{�9�˒ {��HC޻��nS&�#�W-�@U�1���/`��f��`D�=#nk��C��D�b��kbT��~|�@PB�h�4ll���Bj���,�@� ������o�`�����<u&�6B�Q��R�_���p�{#��l�X���&�;��_�A����]� �I�\h'������,�b��j��{�ap��|����uy�`5�t��FõRq3��Wq��l_`K\���Y�H٦]�-S����=����pO�����"g�RsѺE;O2�̠[+;qQ�{���n�����m��җP�du��Lx��Hc��1Z�xA(���j�h�q��uZc�cIE�����6��ͺH��9��Edp,ut
��j;BV,u�`Q��y��`.B��<������Q�I%�v���`��q�$3Uݾ`hsQ�Ǟq�w=RwNP�`I��+�$�r������d}XJ��Z�&1�ɹ���]���f���v�^^>�oҤf��g��8=�E�w�t�W���;S�8nPt"�jr|�PK����P��ŮS�^-� o�c�*�_��&t/��I�@#>��@vx�wA�V\g�F���wTt\����b�൚@3��m@� lu���MptRs��
ڛ	.�4K��V҂��X���"%�����+Ϗ��uvQ\��7QHmd��xK;������G����:S�H7���,bD2`��PQC���9�!��0���TˁB�,�P�&�D/y�}��tMZ	�D08�ë�[Y���̽��������B������g3�~���<<g�s�0���r00���3}ua1�����?3��Q/DHp��t�U£�WT�¸��q5]V��?��_jF9��0;��n"~��=�?��!�GR���"C�����b��alCv(�kh�U+��lxL	���mvɴ  ���8�N��\`;��AA�S��nw�XFxA0Z�&�'��e�J\��{��a�[�v<@�뉛��ؠK}�:�X�{�5$T�-����HȬR�B�6�8rp]�A	�.��FE�G2U��$9~�=Q�xGqʋ�lqF!�apj��=�s}���r�eP���G�o������\���g���i�����:g^��0S �N��?��*�"�����IAr�)-���x�݆�C#2�+�,_9�ʥBZѓ���%i��Ha�n� jf�0��Ԅf��5z�T}m|���op�+,���V��N�N�0�@�R鲆!i�1aֆX͑�c�����SN��4���c!�h,5Fی��c[���H^�Q|�<�Г��,:q� 	4�8~>sy�Q�p#�$ْP�	[��ö�T�̒\��2+c|�����/��}u��;�Ҽ��,,�q���	U�cB���8nX����P)Wd���π�H5x�}P0G��D�G�z]���!-.Sp�Yý�i?��Y���0h�k�	嘮v�=�S4�C�IV,T��/�ލs��os����_�e�������'��T<�r`N�iF�ܖ0�?��ۍk��� ��E�h��fA�� �\�u0�����=)�u��
�_5�s��2|̱�5,B��m4�G`m8ɥ��Ś#!S�1cDz�'����C9�:�ݣ]Zx�T�����K��%нC�����1�z�K1�~�#jwT��m�@D;�!s����:i���,!@5	[�(U3S +dAm�Z���@x��IqmG �})��ʟ�łC?��LOӿ��,9=> �=L�H�Z��@R<����W_�N�XQF�3˻��o����`�������A��;ٞW�C[��zLXʲ/9���N���}�xo�l��o�رr�֝aofU�'CCZjC/.��� ^���b�P�{��ٱ%� e����D���)=|��������e^Nvz(���J�P� @{[tx��U���wr4tl�v��+8l־L%k�Y\*���]~�o�v����0l���O�T����Wo/fy�x�H��ƣr@��jET��,=��Ҥ�`��Q��O:Wŷ�6�dֶQ�(Z�YeNG�hv���qw�����t�m�0`�[�M�K��
l��
-+�W{v��QM0���8vR�A�x��|�I����x���o�6v���ܴJ�>9�[����Ҍ-<N��E�����1�O�3(�͟Y�A�(�by����8�T��(��R�sf�͓kSR� �5�˵ ������D�T��Qc�����w��z@�8�Մ6h�t��y����Q2S����ȵ΄ć��+�/OOnzr�2����*��,��oW�I�\�����3aϘ�z05!�v���;�S�=��S$?���Ij�l�'
-q���BN���jxck�/���Rm�Q��A�� i71F��Z=FJ�p���o�3�BC#�=��P�"�u&�×�Ƃx5��Qɿ��n��F1M�G���>xU�"�����w��P���@�/������_�%G��[#a�,60�a9����X�VC��ζ́��\�˙���d�-3Q"��rs��*�QJװ'��$y��P&��I*m�P�荌!+>�4�n��V�ydsr�}9�� �R�O�Ƀ/�w�βV�2iS3�&�ּ%�"?�	���Â�4�F5����h�F�)���nT-�v�爄�$b���������Գ3XnX�}Yn��cZ,6��k�u�[\� ��� dP��������l���1��d���j^s~�+>�P[,�OeCK�܅bPM[��#CfBf��80
�����]�mc �3�B�a��G�
p{��AU�~Q�������1����Ѧ�@`�hFu��@�\�~��	(��a�)q���r��Ͽ=�u�e�V�t�Rŭ�����4V�vbn�Te5��j�pk���Fx�5�~��G
��]�u#��:2������@ؾ�ԯ��Gc����XB�//2э�6>���L�B�TR�7h�C��G��<��l^Md�s���v�����O�7����A�0��������7�w>ze��G�-��²eںa�m�Y����3�09�� ���z� ��Aɽ��+�� &܍5(����l���q֒a��
Iy�*ci6h�!9����C9�ٙ��� �{��7nTS��K��w��;6#A�S���5hG�b�9�|����,�R��(�59f[x*"�~!�nI��>h�@��͈������+7.9�܍��2_�~��+�0�K��	H�kgcv�91Kn����]��[]�Ћ)�e6:��1n���P�e����U���d��+6�@�imj^w0y�n-6�} P����y�B�jM�%���ъ�j���Y���D&$Ջ���~B�T$�Jf�j:脜��K��?F}���t�F�se$����o7kMr������ir���n�F�pV��')#��]��j�|ׯ�uf�K�3���io�����)P�A��~�c0>��bk@���'������j_=�v۬��m�Q�][#+���U�Kn'�F���9�!k�Ӵ���U��W�����`��Kƽ�vT˾���Ha*���Mj�.�f/)��<^L��*���<��a�׮�[�RY������+~��ޙF�osۤ�A$�_���"\Y�z/ݮ�=��k
����4�^,���Reh6��K\^�Ѻ?�jF~hB�������]\�YעN�[=���X�R��QG	��l�Q Y�0���H�e�/��g����8j����xj�O|��s�|�.��"��]GV�c|�&y�UH��߈����?8=J���K�d��)u�m=�`�y����ȩh��P���[�`�b��{k3���S�AE��������z��*7��.wr�Zʑ�!���/�˳	��X�)D��L�?��Q_ˬd�#����v�}�qRY]�Y&i 嵟�D��||��#ʆ5�E c������Q�7���&�K{X
�0�r �C<������Ub�L�掮�����/V�<��K}]��� ��r6s|)GpF]�z�����'z$��ゎd� 1ςB�����Bqd���ꇠؼ��jsn��=PX2�^�����%�C��oO�;������R��'��^��7F��G?�7<�6L�H�_z�,����8����z9�]iuƁ�7�+�� 3d�3��c`�K�ܭr���)S���Rm+�E~�į��N  �&�V8�����T�%�Ȇӽ������x7��:�!�����%���|�d�gC�����і�_��@�&�O(���,Xi����?%Y��>=�k+,�WSr��$֠oe/W(�=�N9L�w�"��qjG���\�����vٝp�سж{ x�㓵gƇ��[`]k�h�"���<ļso�m����}{1���|c�دG�(��x�y�A���5^�4��*%��c��n,*���_�@���7����x���Յ�k����K'-�>,�ui�Y6�u���j�f�UHi�&1��>f����Ҿq�z���\��Ͷ��B��L�c�u�m���8���1�)'�cG^�l�2�I�`O��bl3uH�?��
 ��������sFo�@_.j����|:�XK= ���1�
��*���كDYD�]8K^!�:����unȗ���H�����e�6.Qb}e��ŘL�؃��)k�8���t4��H��n���i*(���n�t&��_5��o���Hu"3%��&G�Cuc�%ڱ�}!�1*�	�� lވ^'/)�)Z(-P~.A���7_/z@��3��d1q��W�Mu��k�GN�8*��X�L`+8��Lo͖���5)	���osv�[�����&��誚����E[�q����+�j�ܖ=��rstu�V �'8:��4�6�KI#���k���
�ͪ)�y�C�y��瑾;��m�\�$>©�.�wgV�!d�����d����Zy��1�s�:H�	�kl~o6L�yѕ���V��v���C�;�m�%�>����0� ��4{�H��
�� �3�L·�a�S>�����4��+��n��KS�� ��gu��6���a⮻kx�l�4]��/�@s���mc!t���ę"���m���6�E���H�X�AH�F�yFッaL��0�sٹN�0�Ja��ʮv��\FA9��#kŮ�^��@���l1��ר��>
R����)w�� ?��\8��7�iI,o�+�\��7.��܏"���~���wA埰Ƭg��4�ŏ3��=��3�i�gaA�����,ӽK;�H7��D�,N��y��4�Ҩ���y��v]$n2��|E��W�gX�WPS.��At��<�N�Q&8�ݫ/����j���"�;eI��)�i���f����;}��y������ϟ����.X)�?�K�C� [�^QQA��0px�g����l8��GP�����0���K�������L��&
W,�\��I�q�rDJ�|��z)�4H�0�����D�� ߏ�7��F�,W���ݨ��©�I�3'+����-������z���U�����5��`~M(3�p����ύE�����,PGt�(Vd�;U����5��*f����$���`Z�Frt��Uȫ͝�����B��dxt�I_Ԑ��]
,�F���y^l�q}G*���>��U�V:(���ǊGt�w0�����r��ai������4`��@r����&>��{P�� �+���5��P��㢥(����	Ǒ
�"�d���΋�~�G��H��Xd�Oj��2�y�:B���{3�\���y��[\�G �3dБ7��Q2��A��sNg���B>�	�4���@���x�\���zD�f����N�bdDޓpc�(�ZQ��O�:�,�\VC��&�J~�,{�׿^>�z,6m��j��x=�Nߏ���#�(=��hx8Z�e��i�*7�H���	ଌx*��]�ΩU�z��	�Ib�*2c� ��Ω  �	4�&zš8��{Z:Yar���2�Z��{������S���)��z�%C��5����U���)<ءj��@A'^�?��t�?�&�QKNc�c
��w���14K�]�ԚM�R���/��s���n]DUE��q<٨W�.�eKUGa���D��P���
��~�Z/��Tw��!Dj��=�2����7��A��	wm՟�Z��'�0W��Kp�H+~�/��G���#$�M><�3\7�d.IFGS�#e�t�"������ܫ�m�F�t�y�2#g�7@V�T��#hwuS���^ �Z�Z����"z�U��<M�jT�ЫGE�;���H\|B��>@筈ƿ���S�s�w�������	�I���l��5�����b��
��W}��.�__��u���Q��p�}�N����k���
s�Џ��c=�����𗷰�6�i^lX_����L�dh��y^��	l[1.�f`%�Ȩ����&Ls�4�#�`��>ա�P&Xz[�Xm����':��-j�M�!�=z�� a���^��R��������(���h�U�_�����̫���.���z����	�Jg>�B]�rwR����>��^�f|��B��_�ӗ-����5k˪t�m�)^�i���@������a��y��T�
�{��14'��5��)G�c�S:�y��7@����g*M�ꌌ���z�k���, .�$�Sox`K2;2K� �6b^��������(�z(�>Pܭ��ٕܔPw��� �L�� 6��=nj�i�/<�QWg*��o��(�n��*� i�6�.�^���L
���qND�lӡ���g��QԒBaKc��j���9HL���F��9Ngy�X�~@$A09|�o��T�|�"EISGo�np*�(�i�j��Tym����[�:'LO�g�I5�CABRp�c�HZs�nEk��g�KLZ����>���y�p�FT���jS˫���W-��F�c,�,�?^����9��@�x��'��L]E���FI�Fk�MN!|�y�DJ�x���kC��]��e�3�l6�a^߃80q���^�?i�jYX������!�c�:����d@�͕rSe��*��}�����ea������nܟ�%���׊�X�1�%��}!�{��&C�i
�%�inß��c1�P���U�U�r�ֻ
��c�ΗI>nC2�ޝ �~jߌ�<�N���PM���iJ���>�>��Qb���YE��m<�$���-�u;�l�O7���g�d���I��*O��;rHO0H!��ҵ4mPK��.�U�N�vV_�&}05��������+ñ%�D�%5]��V7GY��N[�m.�ؒ�5�N�D�K��b@�b�. pv1PR��CM�SH��>2�� <�Ԥ��B{�O����,�� C��M�)�w��.���^pޠB��Ѣ<�->��l�숔��j��YX��3��9�kN�T�����R��w�tA�����hs\g2k�7�-[�����ji8mƞ[�1#]6Jd�X�
��wc�@����'&�BX9�-���0]�+0t��"5�˙�q郍���K�g�\{<bGx)�1�&⠬�!�;|h�!���V���%��3�[��ɣ���-O��c.E��8���-��9ѼuR�\����pߋW���X��ŒEY���bM'H�S�#� �^�2Ѱq@�XiƵ<��%��?.!\\SEx�~g�i����CL�W��,^f.\*�0[���Ƿ���6^�f��MbҌ�Y9�N`�tA*��Hѕ�Q*�)t1�n��W\��PjH�*�\�Fd�&(��e�IoE
��w��ŉ=l�더Y�����N6�QG]�ۭyQ��?O����Ī4ڞ��*
����XQ�b�J:6w2p�t
�k,	^!j0��^���T�RһȑuR��s����Ó&��| �^�8��(���[�ӳ��҈�����k:!^����t���v�B�jn11�S+�"s�
=���[�Y7t��;p�o;�rQ{�����M��KMo��"a>�83�� �~��'Y�$і?�9u���g�/�:�<.�Ry�N_����,���;ZIlO@`6#?[��.�:������+���
���c�M�YX�N%��УNh��i�r��j�&M��d����=���;h��*j
�j�% o=�C�¹�������D�-��)4����e��� �sU�8�U�����vG��Cʹ$��=ia�I��G�X����M;`d $5/�%��a\*�꒿6��Gv�^9ma�R�����n�yn�,���As�o��(��hOep=�c;g��7_ïm��*��izGK-B���2�:�q����j��R/p��x�1=��g��:� �ڷ��5bBƪ��hm���As��%a��(t a7@�S[�����&j^�d�M��1�̏�4���Ef�6dFN��p�W�BX���Җ� �'�X��-\�鞔��#j�"тh����*UcM�rB�u�s<Tǵ�������XkZs|�f���|$҇�W��}��� mh�(��v�b�_0
pNAq Q�b��-.�do���hcH�I]6��D����]*�
�e?��׺��_~�s%+;�6E��D�r;�LY#^	z�Q6�G��!�â��ϥ��l�/��V�j6|�]	�%�M�S"G��*����FlUH���`5ev}�_�5�W���k�Hy �����v>6�3��b0��1��@��h��4�;����!�~���̺1�������$G��J
<<yfEH�f�H��=�:Jة#(�K��u;^j�q����$����éWz�{]�=p���b�ց؊DD���0�%�
��k'T�%\��<�ަ�,�����@���R�w���Ф��i�Fn����frm|��=�<��큆{��A)��΄%�<��o�_�.W .�������h�S��/E�2w8��=�̍����H}X�����AHZ[\����]���7�(���L���cb 2�R@R���9�s��,tF_,���w���Y%���w2�7��t�V�YAY0�m�����%<D>�=z�B[9J5�x�U�>i�3�pV�+C`hL���W��RA����mZ�v���)le.l������x��Sw�ћ��j��`H�1�Z$X��� �L>[���N�8�/�Oֻ���!j�U�=��)^.T�>6NEL`��z���"W}�ӯ	ݍ� #��r�ߧ���f�k�ߟ�=hq�����u�dՂ�%��<D!� Σ�!���=}�A�}>�MV̝�;�K攵2X8CUߖq������l�#�d�!`��j�-�њ��1w<7A���Y?�b�n��Jg�s0�گ��B�i�O��z��n.f�H�T�2�}5�]�C~*9���dJa��+�91c��6��-N�3L`j���ח��8���Qr r���Y�yCж���+�uFS�ׁM/5AE����l-/Rw�
b��':���F�<4���BOTb)f)�&N�"_�]ߡ_�Z��$�U���j�d�[r�t�
�.6Y��d��*H����~%�F�c�dβ&�y4��	Ch�V��F��%oA�����YFx��Eü�	O�|���NI?L�h"���-U�F�
�k�J��)z��;��q� �c~������"Jw�<*�fϳ�he�I�����{�o[�J��u���)�1�?XH��QB��r�+y��0DI7<�,�n�u����4Ͼ���2F�L�v@�&8ݵ!���\9��g��5�Dr���4"	�;�S������)H�"�K���� [�����d�*N�x�t����a�D򰞆-F��N���;�(�i��BA�'�҇Q@G�q�������]�G�
�3Oe��}	�Yg�v�"s��O��l���I� ^ǺeF�O@��M�I��Ȇ׍Q�7�K�g@��,%���\CZ�U�w&��J�E�aą5x*��:8Թ���d�6�in}�H����!�+x��M�����QQ��ԉ2Lz��ys+<�1�y�u�]K�ɤ'_�lc�:xs]�hr���0߭qs�v�����8�sG��Rw5Ge��F!�]�(c�՚MD��z7�c�4�u)<h��!��~��s���e�Ca3�9�P%��}�M�*�SE��B�=�i/Vg����W\����GeՕ+�ްhhQ����{�@�#Ӟ��G�Ԁ k�9��uJ�\�N�y��Tf�Rp���/b�['��v��$'��Z�c��TR�t6�J���Ч��C�J@��5��*{���W_7�V,_�LL�A9�k?�}q\徜���91�z�ձ*ޟ�|��*"}�ˉ�m��L�:�|�y�4|8���=<��� ��`&î���=r����Sz\)���
V����qB��N��Ti�P�MT`���pۯ�/�(��'�l�5�T��y-o�K��,���,s�i��R��������5��3Fv�\0�ָo�0Y�
i���.��"�ڛ�3>;Ϣ�_7Q0�޸������\������0g�s�!�"�0bD^K�)��
4�������!�u_���p���'@.�v ��#A��H�z_L�8.�8I,G-S˴�4�W�7�!��%Z{��=�;!32�E2�� $TZ�i�*g\a}�u+����Ӌ.�����W�^ �@ܝ~: �[�#� �Y8������9�qU�����&!���jF�+=��8'>.����\j�)hY�����mP���\�۔d�T�<l�j�hP�����ui#,Ο��V-@Izm#�
�e�5;�"=��nౡ�ut����Fa��y���ɝ���*4��xe�P���3��U^�^����kj(��,��ڥ������հJe{��ll����]bD�=ic�׽&`�^򵫨�fl�IAւ����o&S�xZ-�"���Wz^����p�{�d2�-��Lg$eS�Pp�NKPP�f�H8do�X�g4"��w��~k��&�!,t��7t=�S�p:�c9�,�#�,��'#�r2U0�G�AB�jB1ۣ�)� M���+6X�i��� ��g�ý�T�
�S��c۹!���;kG�f�$w�Y_o仂b�5BD� x�YܚՄ����;P,�o���+]#`RO�|-H���d���������>C� ��d�b���!5�����l�͇0�sL��°�G��?
�lǟ��B�ԟM�w{pv��MEƯ�^���s�X)�g��W-&3���8b$�	�{�m+��j�op�8CcL�
��{ �mԫ�c���<�z��$��TI3��i<1�����iG�հ��#���i�a)���-Vl4<kl����$��<F��t������� �O�>�Ǿ+<�8˽��^gX����1x@�9��Ep޹��N�ʵ��KNV3�A.����'x�g�?���حS����
����Η�� ��'��h(��Ƅ��Ff�Y�siQHz��=��[E���h ��<w��-��m������k��.�)��5�~{-g�����t��R�4G9���i���M���cd(kզ6��K��O9^{���)�gy��`�[}n�%"�@��Ǔ�J �~�=\P�y2�fz�/b��>���	Y
۶+{����f�Tts�'U5ʍ^J�@����-����!K�!y�QF�ǘ��s��Ij�Tc�N����suWO������o��_���	�(X�rE���q��X���Od��d
�&�?��|���ײT�e���Z���ɉ_��$i,.����y�r�1u�Xa��U0��*��t͹����4	X;��!2F]�a�i�����$�y���iQu���I���'^��i�%xt��%	'4y��c~���*�b.�ص��mf��*��qB%�nOQ��������H���䠎�O���L\�r#�,���52u���k�uXH�-�D|�W���𪏬���ӦO�"�������"��"a'>����@pA��� ��I<qfs�^�M�;�d���&b3�6��Ga�;�{���%�K��;Hf��|���_�sH
��	 ({O��1X]
�▹ �x|�X䳆�|g��KJC��o� Ys;�!��u��㰠LM1ͼ�
��] 