��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u��	>e3gB�8��![�����1I~"�
7�@�@��;�/Z.	��u�w� R��b窫ٰh���%G(������:ul��&I���|��DZ�#z�Y�^Fk�@$)`!1��.t���^���*_�'3.�'�I�ߋ��Y�����������*Ȣ�.��ea]Z��%���H]�o�"��z��KϾXs^��U5b����Ӆ�-3`��:�J4IK��4 �i�Oё��j>^�!�������J��<}D�c3[v��O�.\��T݀�����u#R5 �v/���o�~.�����ē;�;gg�-�U~J1�az�{�>ʠɡ��DTDC{��:�t�l�A��ׄf�m��,�vh���*��U��0&�}�*mAI�KB���_ϗ��a� �BT�=�;.H� 2�����j����y��z�F�O_��B.�B-�a�!�ng	ZO�p狘��9[\6&gqxl��!�/��}ȉ���,�#�/,}�G�E>�JT&P���$r��L��094�ٖ�����֞�(@�ם@~-z�}��䁈��|}�D�����c Ɲ���>�0ºy<h/���(a@s!ʮ)��3������ZF��f�;g����@��#����}8	�fA�ў2Ѽ,����/d�謘׺��K�:痰��h���,8� �z�>����Q c�$~���(��[�Z�-��^
s\���nï�&��/ z j^�������1Re�vnr?]����ICN\k�%��ɩ�W�D��Z��O�͠�+�'��p�ns��	RZ}ū�K	n����E!i&Ҧ�
s�S,��v�0�X�g�)���:���t:�P���oU�I�_��d-��p{�"l�PY�u	� ԭ�4ہ�H�h�_�F�ᳮ��Q�"��!�4�� =-D
g�?�g���	2P�w�=�}r~މ����,H&i�/V2�N�.Ry���Ě�>�!���m��^�Ӈ��jvz�x��?�n;��hH�8�E��OG�K7�O�?j�\����+uFm� �	�ڡ�#bw/s�,�E܈�9���3Q;�{ܹDc�}D\s^I>�G xl����32�߆�ٝS"�7qT �Y���'�>+w�D�C�a��Z�D�t	�kͩ��^(6�in�������!�\V�4;�����;�?)��[uQl��z�NN�)=d�z��Ƣp�����1AS��Rp��1s${R:��i����Io���#��#K�S1���e���}�ZrM�agߋ�Ņ#䲾�C)q���詬lj�f���� �ie�	ɒy�.����pv�X��n*�@��	��/�h���}���1��6��z��6%y+��"�\$�Ml�����`|Bf�ѽ y��d����o�� ��&��䞚H�!jh��]�)~#��)eybG�5xO1�3,e�!+�-�l�7�I_$"�Zf>�m�a4|��%���m�cp�{S 5NN'A�����6 ���zF�mfLM�;�Px'��Nh�FZ=�Վស>?���;l�	8���+���]k�j�ng��������H���r�*��P��B�",���u����t��w�n��>��6��N���&�Y�.��Ͷ&*��3���� ns���z��e�$��h�� :p
ԓ���P�E��@2V�pk�_Q�Te�ړ<˿ ��pw��"G��hHU�ؖf��쯎)V�w�������P�����iy��~�W�-Y#�H���*Ʃ�3}��X�l0u�si���
s'���L;}�EC������� ����M�!���4y$�(�q?�O�	7H���@�ݳ����HNy�r�<6�땽������s�����N��n�a�Pj�xv2It��K*U� XDY~�v�o{^i��|�*��.!��mU����[�e��ܷ�3���y�?S�h�>%&�h�,C��lx#�6-AA�U�G�Jݟ6����8�gL<zK��mH#FY<���1�Э1.�9��za�5�t��.P"��"���rcyw���t��������r7��Y�@�:eپ�m*9,�NT���YmBn�R�K*�|�1�.(��͘Q�x��E�-�����p-�K�b��)x��n?�4�Q���_3i������8��lQz��Q7�4��>��]��Y�a��2d���e��L����P��v��2|�<5��{���.�~���U\9�O�P�q�m�����1����N����d1���J��bc	0��b��񎎢]�r�Zl�i$k�t0�����;zk�� �	d���4�?x:��|�"h��=ZF#��`Is'����sU��dE���@�+N¹��G5]�!��K��d�)�aOr�v;P��"1�7�T��a`��)ݤ3�'A|�G���J�xNv��f�_5�^�ߐ�z�u����C�o����Jk��%1{�m:�b����@�a�(ye�8K���A�f��������-�zL���+����?���f�5�1�g�O�4v?�jc�u�R5�3�
�����IQ۬�c�앿�m������[�I*aaa�c��a����r8e�o�7<��H���qnw���ޯ/~:E�(��$�,��2h�Џo��4���*9�����s����%ݡ�٬��O>�<�T��������t�����W0�AM$y�=֚��l��1:c6r`SꝠz��^1#	�J51�.R�'3�����x��c��?�a�x�S@b
j�����n�iv��~أA���o��2��E�7�1��Feʦ�>�%3]��MC7��b��$��dx�� �gx��R�'(��N�8S�/奜�W�=�Xʧ���l,���HMW�J���(�UE�s�a�!�_윗��R$�{�)h� ��Ө�%�%�X0"*��}'��W����p�c��B��H6/܀c�>�t3V��"�rGUwr�m��k;����e�s�P���G��z˯{���hw��w�'�Z|6�:�ƌX2�B�nB%
��)�qrt�2D�R��F��jM/��T���p`U�@�J��e�.��"��F���0��wΫ=���Ǭ�-RBQ�.X}.��B�;7�4�'�Gi�kB��I(�d������-F�c���tU[�8��2��f23�z�o��é�T
�����T�F�1h=8%�aD9Z�C,G�μfjr*�
����Z{�J�� 
��Yדf��ۄ�ނ70XXrY`��UUJ5�dX�ˣ���CF������$���-��»6� �{,��\I��I-�h����g`	뮞����4;�ހ����h��bu� ���AF�����h�z�?穈T�ġ������1}��ʃ�