��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~��o��p�t�zsC�r��� 7�˰X>�S��4@��TI<�⳶T2���T��y�/p��	�����v���Z�V
�k%c:���^Е/a�w��k3���9�C[����yXE�J��cHїKt�۴�$�����3c��n��K�e�]�H��� ږ�t(�x���+���96㵚ǈ��
��!�~�iEfqR}c��ةpȔj���Z��]N��FmC9�� 6��:�&������$��P{�:?����i�3N����|d<�Q��?�ظ���j�g�@�/��6IW{��v>�זm!��t��dBKr�&&9���}κ���uSK�`��I�#�i������:��/h6��1�=�֖S���%��ϣ2����"���.�Y4������ժ��k�v|�9B�Ȧe��fv�{Rۄn����aE$��ל:�P!p�D�P�˶{�e����o�s�
=+�H�6>��9iR��3���dD��rF���wZwǐ�,q*��}�ܙ���I�zb}���B�;�f��C dj�[Ǯ% ��h��'��YH����{@�+��|hݷ�P���Y9bV��X�`����F�;��!l��;�Wu�8��]c�c�����y=q�z�J�(N�w���N�	��h>�6P�[�u��� ��\���@��[�g��=|�X Y�E7��$�k�)�!K�!n$�e�	����~h⌬��¹(��J�o��F)��W��F�F��%/`��?���T��W�gD�.�w^ü7C������1	-~3ߍI�+S��C>�%tO:�$Zg�%a�R���Qտ>i���:{+rM��-�e�����0�y7n�����VMؘ�-�kA��:�d�'�@�׆F��$�1�� ��
X��z�)$"�jv=�)q��M���Q�&�":5Q���5�X�i�e��
k��t��Up->�t��Y_U�CIGj�k�9[�o�%jzid�Ց�fnP��V�|����Š��S�ý,o�Mj�ߎ�Z�`� YH��j�9��,�1^��e��Ƈ�0Q�����~}/n���&.1jݤ�OƬ���ښ�Lh (���~�I���L �0b�Nn�����^����	|L��h��Dufed�^�8�L��z��,�:�υy�r�VN4^�����>����ǖAH�a:��V}5�<�h�*�[����N���x�72ZD��}��?���˸�xj���u��o�8�S�d�6ΩJ�F9V���=���W�S}�}�jCy��ϘWtE�y��*�t��|^��ς,�y��`���>]�K&����&�V��Z
�«+V�Q��᠟Oh�K��]��ˏ��n��-���f/�����š�P��	�=p������7~�R�9��t�����m���*#F!4����$=�r��?0�-gI���J�P�s؁b�+�FuPv��;� )R�`�����|���7����;,-z�>�"��	z�����6��)m^X��ly,Z��]�s� �V;�_\a�G&�����a�)G�M�Ŕ?�2o�I���>%Ϯ��F�SB�j��'@�E�M{S�sFiu�{~wS�	y-�>gV�E@�h�_J�`��OW�+\ih����t��Nf�\�Yv�]?�d� ��=s���B�%���E?-E-����m��Dd��H�y1s]�q�`�'RxړG��z��7��̟�����Ƙ{�ܱY�^��/�A��dƷ�c1Z��j1�0��^"�9$Gg��NN�����c���譫��72Q� ����F���փ����KH�����xv+���y3-خ��usI)�@��¡�*�DM���=��]����c�B���}W/�ٷ7�Z����🫨~�),�.��Ie�����^(DpF������3'͊��%�L��M�c��6��J�n~���g����� �Ot���(�Q{le4>������7�<,�*/�`Kp��
��&Ŧ���[K�yp��!��g�4��'#��=_z�\��&(��2c��/X��a�E�:��@B-��>0�_6��5��[6_��-��6X&So��-�r�b�K����+k�05���*�wH��xO���򹢗�H��PA��	��\GT�b��=Ԯ5Z��;pߍ��.o�lq�]|��f=�75��\�T����� �����S��ź�F�Gd�j��4un�+��*��f�G�<�нx2����"��FBK��I�v�1"&]aE1�M���[�����t���vH�3�O�~<�X�x=���5����zy���&n^�Y���	�nv��r��H�ӣ1����=m�&W��A*}ϴ��/��
U�#�Qqp�?�;>fJ�an{�xߙђ�;b��q]��^o=:�w�V�C��q���أM�`f�&٦;W���/�����9ּQ���"D^���~Pb���ne&Ȋf���_;�J![�GS؟��1Ϻ�wr�|�*�ffJ�ϣ��{���g�4�xsR~t�A��؈��fUa߱ J�H]��h�:���9���2��t���}���� ;���E��b]�pV�UU�%� �F"��He[8�[G'�In�Vv�Er."�^D:��En:1:�-��uwc��Å!m�x�伒���`��c^" L�\Z@:R�����m9R�0�B�L �B���=���Xe������0o�p>i��%�$=��}��S5�15�������2QSјG�>���×��Z򞵽�!��z��6��c��1�%$�6��t��:@��՗ܛ��"[��K���!��chS�኶�iE�H�W��$��~,�����M�RGo;������r4��h�S�+!�=��[�G|�w�K��s�V����Q�q�����T��7��>��)���,'S.O��T�@��U�tQ�����i ��h�����4E�<҉��VV��z~��[�Z+B���˨t-��J�gK������ǿ�E��CF����|��v6�.4�L������x���p���1�J�ܕT�}�i#i�c��g����\��A]}o��jq�K��]�GW��i�*kb ��ٍ�/,,/Z���Z�5�ڦ��N��͡X�<��3�e�e��E�Sf������� �O1���#�A#�<hŨpҫ��S�x����/PI ްgQ��UZ�ݗ�ƹ+|�����9�F%.�q�ʁ��oc�80x��C+^�&	�Ci��鯻���`�%���3�ixk8dU5b���z��D�.pVt��u	m_w{2|iK�~L`�D�(���>OIZ����ڡh��ߔ���������%e'�]k�Ǳ2t;,�լ�Ӎ8%R�;��zNh8Ν*f���L�Z�ԊX�	T%�s}�ڵ"1�'�NI��<��2�Z=�έ^����|=��5�k4%s}�b���C�����3��;�t2�j]�kF���ǛR�|u�Gx�|i�7'f��L\�sʾ���j\N�>�.^QT� Θڝ��.�vO2���\�)�ںi~��	:(M��g x������"J7^�+��ts��T���i�^�F��x�7��q���!0��l�"\#^7jZ�n�qg�
�LāƓϱ�H�e9���(TM_{|U�pm?v\ �����M�_��<�As���������Z\�A���ZZ��+�%�+�#�1u�%��jT����+1P$�Ȱvo��(2j|�]�
�{d�{��d�LS
��W���������^$��S#>�gX��@������Q�u�Z'��dX������&��y��KU�x�<�.&w���P�µ�+O����:�z�_�/��~F�5F���[0�jn%[�n�\]�ZI�i�T��hu!UY�ʥ�bb�c�y��_ǗKn�.�Pq�n������)&��ʇcSi�M�9`�C+�ZG^�8�F�-��� jj��9F�� ��B�H�EQ�M���&�Y�|t`����i�g��
��st��f�Vpw�҈�؉�����H�f�w �5�[t� �Q0ѝc?���kf��� ���y��eT]���+�Ь5a����ɦ��'�s�d�n@3�{�;-��Ɩȉ��T���D�2�SB�b��g�1a�N�#�@'�_������"���U���1�eH���+��#����Q �|�m��,ὍNP1��]>ױ�Y[�-�75L�W�� ?�)~f��Z������!�u8�>�M.��$M������!q�c`����XXN޲E��F�����Q�@@�|G!^����-p ��$�T1��iR��s]MKй���<�$v�������r�)L��s�o�]�9�t�r�ڤ��`:�J]ҕ�?��2�v�M��6=Z�LKis�Ӿ����1ȉ.�m�|wd�0z��~��r��IBэ2X�I�ay��\H�>�^�:�j�}����S	�:eP�ْ('�I�U�_�����:�~	�L��S~��NǙ�y�-C���((��6�R����?�p𔳖���\���ޒkRz't=|��jjUP<7Հ�6��>��ݔ;�˾�md��.����h�>���m:D��׀j�N2*1���rۺl<�T���"(�[�F!�}#^.�_�c����}�{�;r낵�o����佚��\�~}��=�6�C���ʒ�N��@�V�D��>��DF���0hΥ�r3��۾�G���}è�~v�ԹR�F[�n:(
$J�H�)�Z+� ���Y���
g�"q9���f�
�9%�}�G�/d��"��Nٯ� ~ǅN����_�����E��󐝡���ZD���<V^I)��_�f�����Z��=l\{����FF��e~��aZ
3��%ܛ�fd��3B=OTzp̗X���5�v8�2����mO�,Y�j��&R�=8����P�X~O�����������f��z!��m2���B�S���śԕ(�%�pp��c�r2�c�lM۝�x/ο=;~�$(��cBr2\���h�⻽�tz;ϥ)A�6�<&��//ʴ�_|���P�vv�1f�欭Wl8YL�pAU8Ku�+�?��濻������H%�?�����g�)9�N���Y:���_2�G^9�u���(�':��a����H� ��;��M�gZ�HA�*1+VR�8����z�����)�V{%�J#���S�C�X�t��j�wF�Y��wU �1��v�m�h��G�/��)�&&ъ��� ���[)��ߠ��Y"������b�S�=�N��(PΊ±f�� ��<��e�^1��z�L���aA�S�/��N���aR�?��pD{��Ȟ�����!�6ٗ�#B��g!mTx���2���<���+t+����B��r��dK �Tzo��[&�L4®G����j��R����A�r�xD��=瞯m�/�F`S!�E7\{mU~]����٧K�|}7����DX��{I���q;u���֨�6<w!��疕�WQ�<�<��`����뙈n�F!�G�T��'3;S���i6(㹋6N�A���F�U���c@��4�S�3Ց������ �z�x@���2��g�iC-|��F �:l<m�H��[���|�n$�v=�(��k��Ue�,E�����f��{�,�������=B1�}[-��>�#nh
y�b<5�aEO����>���YK��f���mE c�o�4a�����魘u�����Z6=�����ld��7:|���,g rg3�~_"|z�ᶓ��8Y���f٢�N�o�a�E��ZG��RdE�k��HϕFG��9��I��O��v�'%�����^T=��x]�-s{1�����v����5E��mMg�c�����㱸�7(.R���0�^�N[�L�;7�FQ1 �s F���wcp�,��f��D�P_��QV��ݧ��i�Y���+��-70��v��AI�!���R��[���K�H�̀H�6�|���g�rۭ�+���rE��N�߀�������M��8%�gHh���UM8�q��$��gh���-��b�kV�}�%61�9��M�0r<�N�+���ie����D��d������R���%y)�F��3��A*m�wؐ�g�p��KS����i-���jZR�$�v�n�ꌞ��#��~�b�N�"�ZB���cm![�3U"����Sx��TI��!�/��@$ڈ;�q�13�F��4��Y������r ���29'�]s:��(6K�U�99�֍ ��پ�=/䝼�f�  �<d�B�=n�E�j��s�Xx��e^~��.�h�?���T��͚~��h��8S���o��k� ��qZ�<��3�����i/�e�
��QӋ�HG}�#��X�zԀ�5gc���5��� h�����#%h�Eu��l�׏2j�q7;F"Nlo~��T�6�����a~�Y �����Y��՟�F�ٻ���J���\�<�����[贱uz�l�x�tq��"����I��撠�R�|G�6X�g���x�m_K�9I����m��Eu��.��f�l��'V��髭q��u���A)48���rM�L)����9!�V^����#P,��M6�r`U�j�"�ۨ�1S0���B����{r݁5#�q��,�'�;3%��,{8cj���\��:�({���:�Ҽ�!Ȥ�!k)��'C �- �nԟ_�(��^+�F��RoS�-���({`gN�3N����+��#�.�'(�e���8�����Oѯa�Ꮂ��K��G�B�-�$,�ٯ炓|��S�Q�Lh_��}�:g�
�^-3yT&��p�ѿ�2~M�BC�! �Y����#�K�ǵ�t�/[d\>J�G�E%�C�_�WxB�"@&W�P/��\;	�c�E�!� KJ,�,>��-��B��C������������E7���M���fI�;G�%��!��z�nJe3����Z��6��OFɖ��:&i��̋�=� ��<8�x�T�!��k1�3r{U�f��+jd.Ps���i�����v���ʌT�&&��1	m*EӨ%�hG��b6V�Q������ ��}�bg�쩟��\F�^ZOY����=!3fߓ���+��m'P45 !���9�'��"z�_��$�״�ʚ�iQ�I�*�czO�=A�_��?1٘]u���/� �rrC�4>pCdP���`TS���X5e��fi��}C��ap?d����l�^�t>x��|��Bsr��hO3u��~V�N���PY̩��%��m>j��^"wĎ��y��ҟmW�'�g#�+p���b@G��TV���lɿz���%�浽%6�5ͻ}ѪO���������Q����D �����3`�������hR�l���n�k�N�7K�8Yƨ3�����̽�y?G��>�0X��4x�,�V<5��l:;���9��[�% <��>3:/Cy��9���;����I�	� #�ލy��i���)�NxO�#vJ-ukA].�2lGj����w��cM�O���t8����zf�:�;���<���$y����T�2I+�����8�6�[ +�T�&���9�6ȏH>�bf߻�[�b�� �9������dW[�1^^X���g'�V�+$�J�/ݐ�	 �����̮GŁ��D�t`�<��D�V����s��~mf�5y�6q̭��t��'J��Η3U���7��&}Yש 迏ۢܵ�d�8P�wy����b��3���c��6��Vm�8�鲙Ġ�r�[�3�
�6��
�.<<�Vkܾ�!�J.�9�;!����]>_+86������D�K�/1�s9�Wt�>'�L,�� c�%�0c�t��.����V[�WSH.֯r`�_�A��2�`:��:��_��tQ025��C�����&Em�f�T��>]�ӽ#��Y�Ix�?zސV'T�&�DUm� k�r�SkC�y����@ܦw�̌64�?���8�ߘU��zv�O�<�ڼ��!wN�>	�\��8{�8�6���S�|�����I"6e��t�h��o���H�����8�R�����:�V��ض����I���ο�}���4�v���w<���nˌL�6Lҙp��U]P���(�M�����U[s��ʚߎH���Oz�˷�0U��Xz���������-�i���DB5��''60�x��$�J̅4�wb�3��P�l�];�d�}]IC�W#4Ԙ�װq�+5
���7d��up�<Z# O�4�>��-�N���x"�kL߂N)�$�U8�\��r�Pc泃�ܩKfN�L�u���7ǔ�+���6�;y�Ԕ����V��׽���.6C�l�-Q�F�;��}��,VJ@A��聏�����T�̨-c��-`���@�E��;�J�D#�f�&OFjj�B0 �^V�ӊ*��omq������{��u<���1yWP���l�>e,���L�9����\�@�Mc:�o�8�������֊����h�(v���J��f@�w�p85��K�^�U�*��n����m�;����11y*��)&5}-�=�r��.J��Vr���-��������Z��_��N�(xM���j��|x�Fo�Pu���Y3�=Lm�:���łA,KN@"�0z��du{� �;������,sd�'h	2z|S3����َ�c�� {�cavRe8���]�\U��ޛ�wJ�Db�AQ9�n)�J�6�φ�f��=�biU��-=����x3V[)�Ƨ��f�q cN�qٱ���I(�Ae��$o��ENn�z�Iґ��$�P88in����,d�����_�S�������.G��G���|̍U��� ���B�ˊOힵBI:�x9��8�yȐ�n��XC��S�\�/�;K�� &H�F��(�B�P�E�# f����S�{����1x.wl�-�P�����}�@�\�8Sf{V�����Y{���̥y�>A>����ȡQ)I��?˽���zGQ�/w�$��~�^�7��ʍu���	�hg��Z]��1@q��Le
�G���#����{KN�K�L�h���6Q;�-�lh�-�<� R����ݡ(g6�q�½��\2���E�fm�dfP[���:��`�a{��[B~]��5N\�_��v�aߩ�~�s��qFx{waG=�����2:B\3Q-�Գ��w�29���v�l������k���l&�&m�Y��w{�:��� e�.8EH���u@��n��;Sx�� �@>���X��\[c��@tN�����4��A���;��� h4����ϯ���3�2eo՝P^&F�:��d���iP�g9�/���4Z��6�T�m�� ��A׷��,�0�!�tZ|޵���S-چ�g������E��vdk���8��(5T�2_�~t|�MÆ���xdpkOoq�Jv[ɮrx�Ҕ�I�Y�H?�C}�x��H��V���2�w)� ����Ǉ)��9�OP��A�c	�F�1>� ���r���2[�Wשu�)�A�\�� ��U�w��%�vlȰt�dB�fT}�ro�1
��تuZKr;]��=VK<�cls׊�K*3�Iġ% �8l�C��vK[���3�����bDIo%�=���Xl
N���ܷ-�5�C�i��z�X}��*�hA@�U#[v�t�6&A;�ز�|:�%pGd�{M-�&���S	C3��hX�ָ���X�Sqe~�W3��0A<5��XS�@���R�d7�j挴��n�?�f����2H
�R�"��ƼlV;D�^z+�l&�nӮ\Y�;,���c�Q�'���O���C�ɞ.?��d�c�(�Wpe<謙�WJJwK�p�Ï�ul^�2l��k�r��{,B�&�35�=�n1�O��Q.J������b.�0�/����E%v-��/�i�8�����]����3�N�o	�rg����xĨ֪�� �HtEV�>X�knn����C`����c�̯��m����P)5nI:N�֯]����{���A��'ۗ-�q��h�R}��W��ڬV���*M�,�G��L91��1�H��T�콙������Aͫ�������
P��������QH�ME!���Ͳn��r�
���:h�s���@D$�fE�/cQ��@S\�ݏ��?"�������_%{%#�ֽ)۟q ��|�j� ��e�<9�D��W����<]��_�E�,���ǿh	�B �����ɪ�	�F�S�y�X�AqH��|W���o��+))��b�{#����W'㸿�G�$*n\��W�=mEpK���g ����h����S���.�DrW��Oֹ�RPƕ��*,��5U PdA�̯�?i��໮�}��׌��HdF�=��y���� ����j�}4BM��q"�:����*��Ae��W�p(ֲ�x�a1q�3��?�NT�r��G�����J$�w���vM w�����NCiOs�ح��	����>�\���?RC���-�U�T�n�#��|`|����b����i�}�M�7'�,wk-��Ҭ�f^�7�H/R�c^Ο
[t��x�m0-6
���	�Ϊ�)�Ѣ�\kG�QpB�N-,S 0/����C��y��ة�e��)��J��v�]�@�E���Ӆ�W����ʯ���[��3�j�U%��-�f*	%ҋ����no�c{�v�LA��Da�M��J�iռ�d�n����p������E��@ȹt�?ݒb��JG0g ���SS#������j�驩���Ω3�06���#p��>Y�\�1;� Sg�A��u%&�q�!�B#Ę�t���J3�Bb6���i!�^�@K�N��k�QL���-���tJY&��w�U��ym����ֱ�/��3��=�X��J�)��������ܾU�\�@�|%U��Ξ��V?[���c\�tf t��5�+�2��.]�(l��%��U�Ga��ǫ�Y�p1�(z7 �p���d?���j��͓�T�J������Xdo�љ�>W��G�V�`�֛Ns)��v�n5� `�;I��H�!'�s� I4F�����l��^$Gq׊E�x���a_h $ �D�i��c��BJ��bw��r��b�v��u���E���{�����0�	ih<���!�z�.�cq3��G��c�{i���r������'�Q�4(��
s��=	�=4L����{��pU��ub%>��O�d��UO_�e	~�<����V	Q��6�Ye9�|A�
��N�v�7�Ce-�{�a��S���[���F��+����7]rȜ��v{�M1�2���ء��q�H(�K���3u=כ����z�
73�K��p컑Ҭ�+������ă�ޫ�����ѳ���P�2��l4?����
��PM&m�TnU$M5��gP�|�4ڂ8�( *QV��|�G�����+S��d�r��\S߮��E�i,�{ғi`�ز\�����_�O�P~;%|�d��k�'qǹ1�9c��ꐥ�g������JE�� ����:����	�`���JL�A�m�B,��O(�)����WD��=sȵ8����u.�=���y@su��ۭ�!�ɛ��߈��H2aB�����M��b(���;`>����߸4�kTIC�$bZ�rfy�[�O�si��u��1��8:d��A��;�^��rB�}vx���>b�¡�$7��o��Vf�Z|��ã����]�����%oS�Im�i�I��BA��_`�	�.����C�},x3z�M����L�������k)� ���ggDcBwq���b<}�̬�?��I\O�ƶG哊����u�I��2����,_ݝ{����j��@*&�L~Kw|��#�޻��M��X���۶R�q����!9Ш|գ�@�4�����6�f�;)�U��;�[y��0"\���ܦ}��<xW�1f�>��~7��0��}��N�c�~g�(���sO�T]�ܷ*-���UU;���"��n)v�)�W�BTǎ��Bo�*��h�i,�	��6훬OrÞcpҫ����y�� H2f������O/p��Iq*C�ɜ1M��p�h���H�/S�Ϊ�?f�gH��Q*��8��7�H��6/ĭ����3��V]�S�C:!��IG�ٍzv���/�DNO����tw���We��V�bY]X�;��'�9�C�ɶi!`���4a�>��U{��0lt_ѿm�6� ��U���ܭ�m_](�b��A��cp��~���]�cDzk$kv�W����j�ӧ�מ��a[��Y���]��-�v(�)�Eq�}�(�]y �m�F��@�E�M��� �{s�4P���v���/�d��w6�H��RS8�=Q��@f�ݐ����	H�<'���Ni(�> A��BhZ>����	lU� {4Q�^(��\PW��ʡ'����#����`J;����������iV|>��?M��E���� ��j�ߤ����O�{a!���i��;g4s(�~!V/�j��0*��X�Q.goEy_L�^�cw]N����S�_N)�`2ԵS�X��&�ꊋ+`�����_��g�MHU��{7��8"q�fY6i��4S���<�&u9�5U���c�>��vuՌ��v��옝oa,���[��
F�!���' ��m1�0��떠4�� `�m����Vi��}Ǧ�ai��Z~�֤e�=�@��2���9�qSH,��Z��٭�&C���QE�N�/��aeX�ZyB�"��Vu�VC��E�k��-����[spÀ�/SO	1YI�@�ՙ��A�TWl�A���P����q��l���8��!i0�
�04ҜJ<j�rb)d��nC��(��v��C�r>	��.�#ܢ�/�x�$�XC��.��,�K���EWh/��z�����E�s�뗨���J (� �Z]h�|6����t���f�Ǆ\3ێyc�.h@%�`rr?+�G��p�%���-qY�θ��/v�|Vyu�j­�f~���01��9����u;(a"k@Z�Jͷ�}+�h�W��w�w՟�P�*ظc��=p	�E�$��U����*ִ ����MD�n��?�b�m�*^�}��+�٭b���h�n�^����ƹ��d�1����XI�3����q��>XS�>� {ޮ�
��x�F�%^8�w�N�}�T[����$ �eg�%��q
r�>MdɻMQ	�������0��l��`pۘ���ڮM���>��^tB)3*�Eyu;���g$"!�'?�Q���"��8@WY.PGE�lqH`�ߙ�p�0H�no;��ô|���*�h:����e�&H>��8�@p#�a���8H���7F����Ni����5[�����]���'y䦛�����Y��٧�J�mE�db|v�ޯ�"��~��x��>���m�<�쟥NF_�,0T��pǌ�r��+�w�L�ZO8����U$t�l�kd�VE���E3bC�靆����[m��X��3S��Q��i2�yꦾ�R�8�\`F�P+�>�?�D�@���$�����o%EI:��\+;�#�w(�B�014���ǁ�_�Zi�ܼ�ܞ�0Mͳ����X�ɉ���}�����pc��'�l
���e���N���!2jWBs�Q��^R�쪀͝5�sYW����?0�=A#I�▶E��BEC%�=�J��Pgf`�R9D�e!������|������������U��m�`�Z ���d������x ]���<��	�k�괓"�vz���J�h���;L�r���r�Y��=�;`-�sAS�)Q2$k_�1��<�?%f��z�"�]��b/��\���eMR���Q�]�y���|u[L>��&�v@���L�<i{i3Sd+�4F����Đ
��j������@s������A����ۂ��%�K���e	�������ȋ9����D�_���֠��eIZ #=r)�ܢ���:�֊��V$�)��N��U��0�����$��س���$�!�^�n�G��n�3Q����wZ!�w�.�<�߯���UM5x�$Llf�t�s@�śd��Ɖ9�O�G����|���`�������kS�V�&��e�\��!�W�QOK�hKF���f�	w΂Ǽe�����e\^g3P�+� ��/�����.����t}K�Dl� !��`i-����tھ!F�S�:x�`Ia)`�*ͳ���p_��ЛK��[^$�v<>�Z�(��ꡌ5�vZ��@�1Ѭ�X���i�T�hR���156��9K[w�q�f=��Ӱ%Ϛ��6����[���Z�������K���5��⻡��C�_���w���8zx�q����W��$9m�U��1ZVį�'+E�ӈ�׽㔟�	Q��W t�tu��CޓQ���V[�#6���ea�����X�a�;�lJQ@�qf��r���3�Տ�Z]��Z(����]�<p��̅&��Ix�\�X"u�-�	;}y����C�GV�<����rCݵ#��8B�d}� Q������`@�u���?�aR���PD�� C��U�X!������0�<(vE	A�	��ϞC��q�h2��j�=���w��w��������`��@M��>���M�j(��|���T�����Av�s]9���P�2��!N`�U6Hz��x��J	��+1'a�c��k�kG�OI������������h$�O�z��k�=0�t�#�6P�+������72��tXn��E���ex�ק��4����o���	Ѭ?&�d�f�@�
��H�?���"��L�"�z��q{pO�*�
��G\�ό��F�yW٢ZZ1o��%��+TG�E��ej�;��ٓt�����Y<����q�F�%ќe�fc;�Z_TI]��'JwS�o�8aA�2OK��J�I�o���r�D�v�݉�:�Hx�Fa�x��M��)mv�)wj�K%��4w��.m	�!�8E���|���*S�� G���=��(.�;e���� 9�b�X��	��6�S�_�Vj��E!"������[�N��n�\�����([�?B�w����ٲC��Z	��q;?/��t!WPer��G[�m�:[qD��K��]s��%�Fj=���Mc��|{?��}�!ؙ�F��D��ݤ�Rw[�:PQ�wz���(��- Ʋ�9�((��"���Y�a�b¹���q�$�+ծT��2mƑ���󒃯BG�K���D�:���m��{q����!�2˙�>���}%��DUdg�)FDL�;{)�*��֥�ҫaU-�:gE�m�^�HpVy͋Ǡ����4��Wv�V��)�M�O5� r��/�qB0"z�"	<�J>�;���Q,�7��n�KW>ܮSP	U�4?�F���<����dr�}�3�GEQ�)oP�'A��3Ŝg��gUț�HL%0����jݞ#9���yr�iL���� ��[��h�7�Tf�Xw��Ф�Y��)�Y�5���YX�mϲ�bV#������:����u����X�<�,~,����ѐ�Ds����p<)���q�pM�5��w���g�ɜz?�i̵���(���J�ETt������G��o�˶���a咷h~1�e��������7���,υ����v�Yjz�~�AD��G	�kP|��$���' �T��s8�q��WUwIL�"d����鴐i�4%iP��߹1d��IS�'̯^:�W$�⇱y�R�~sL��&�	��l�)|��D
¨�W�a��CTn�X(9��3�����O�����I���vR&����H�̹��I>泹� p�.a5��}t.|�ܞe�����D��|���R����T���׶��h�t�ϔ���)����X��6ݳaI��?_K�0pTv��T%�TL�^t�������܊� �|f\O�(��T�ۣ�.��ɠ�%��WkX�
�و{����V+iM��	\�g56m�hDY7��ow1
l�{��&0��sН���cH�i����?
��� $�����Ŕ��%v4��<�~��C>
I.j�Ԣ&p	���J[���;� ��t�"��(Y�
+�I/��E�ݾ�4��p�1zD�W7�H��0�"e��n'��f3s�r�z4�
Px F.+��v22�IG-�^�\�S5[��/��sԹʹD} �kqo�Qi���<ԭ�X��m+�Y�)���ֵE+e�?��Ʋ&��������J+^�-<U�RR��5�T6�t��b��
:��sz]:Ȥ�+'��/�"��9*gM�Hc�x�H&���L�'���A�;7�"���Z~�D�I��x2����;]�|��<zO�޻7��$�!�¾E�.e�N����<G�L��gŉ�w���������h��Ц��:�S�:N��/~����
d����چ�0�(��o����v+���i@P��}�"�N;�2�w��H+?����f�D-MK�N�,-u��c۶qK�jtm�:'$rd�y^�s�#d���ߐ�4i,�F���ݘ�%���V�5s-�xG���9C��@��^�=Z�3��^l'�z����_����Dfc+��!HH��ܺyPx�����n��/������&�U�i^��J�3���$OC����7~ʈx^�h���{��O��T��ܒ��p�_����Xv�c�á��)˖�<�p��<��8W:��q�����-�ҋ�ee������>��JR#���N�y:��Tn]j�^W��>�2��cD���N��݂�ݬ��"c�ǿ��/r��v�^ls�c�P�<�S�ސ+\��/Q�s_�D�'�#�(�Js���|��q�>3��I��F�{'y3v�Cޖ��ú�̳� �:��b*��E��SMɧmU�b W2�!��eMጀD�f��vw��Θ��l͇��Jr���w9���0휂����K�2v&�%5�j>�D�� �*uF�I�!�h�j���`��Q�ݨ%�ަ/�17�_� O����R�&W���r���X�<�w<��ʦքu�����H(�^�qЙB��^_O�h߾e�*�`�V���!ME���y��c3I@����0����P���b�Gqq�R��塐"I��P�u�Q���;�c��u�`=���Vb��@ �u��<-�[/��u��'��f�z�爄`����֝��TL�%ﯩ��V�H�1'L\R#����qw$2l�W`I��)��p�Y�˚.��ׂ����`��\4����'o�b2��|aCH�Xzs���li �_��医;���M���c�|#8۸� 3=>R��W�3�����$ӓbj�)�Z��n˦OAd�e2��dc��!�����ފ���z��}6Y�YR�B�lw���D��9� �D"s�	�v.j\�7�S��J�rI�eu�X!�A�ǍT�A$�,X��v:s%��C.�k3pP�JJ��g�*i�@��vы:9M������g�f�?I��|+��EtC�׽�*�B�������"�rQ:
$�;���ua�%���H�N,!��1:��k���rUh�'��K�#¨Rs�k��*z���*f�M��(���s22ma��#�fvb�r�����e��s���`_"�9�������2S�� ���v[�<���4k��43��uE�h�V�vX�ι�\��f:��	o��]q*4(��*d���f�I��<����{<?�cZ\a'2�TX�8�`����=���3Z��qj]�a؂�c���iK�	�ilhͲhG�}'F@\οO71g�-EES��I��RD�و��e�P�Mx]���,�3�a�?�C��Bh�����_�7�Ʌ���Mh�~�����O���󍒳uH������8�fv2J��b��q"ց7b�<{�=3f����|.u���@T�\l���nU��*`��Qbc��S�J+ qm��ˊ�O�_Y��CQ����+�*�}:��T�[�q����
G��	�4�(?|��?4?��`1��:F/���� 0".�8��Q�I���7���0�(&j����*�/��~���.7��͙���QJg+�X�.m�ѓ�R�ީ�a��ROh'�@�e-�P�S��0�Jn�`b�8�t<�@#����S���F����Nz{PH=^ҫ���@��z�9�W�u�x&=���h~͇Cz�h�5̦���]-�u��x�ڝ�j�&좺/����UQ	�K���?�b�BC�0��G��h�A}هw��!�s{q��}�!I*��w ��CD��"����5R�/WnF�xVdw��z��Yڵ;����xF0�HΆu�g��kp&���*ĈLFų���׳�?��2����DER��H��D� 3���\���'�{��h��&T.n��g�8�9YvJ��0\�˶�'���I'�81��/�⚷�D��by4D���c��+C:��whu���t�� ��8[#Q��L�u26�cġ�r��K�V�嵼�B��WHZ�����xC?NJ~�H��`�Ê4�÷1	���#!s��Ů�"�/;+.M����M��ع�{�.wQC N��"�q.�9Vy� �/�ɋZ��Y��~�z�C����q`!Ln���$���AiN_��v̨Ş�ͳ�	�SÂKI��w�(��H9�������G�$��=sY!�4�<�{�@
�`�6�T��@u�j��J�n6����:*b-�6�'��à�/"_���q��ȉ"Br�MQ�e���N5���o0|x8����Y��̹#���t��ҏ�T��䓀pnD�P'��:v�x���o��W~)\���8��A/�Z>2H�_�fe&H^/�oY�1uGq�����6����di���C����p`7}��P���F+4���	����P�:�8������0�>�i�l8��dji��w�o�.�Ŭ��o�^P7%� E}= ��as���B�T���F������Iq�(���NȊT����6�*~��_�ZcSX�[$MK�kc]7Ѷ{^ؿ
"�f�� ��Ss`���H�\���G!18�W��1��:���O���Z�U��'�xUpX�iW�x��ӿY���y��6:!��B{(���ќa���+���*���0;)�h.+��?��i]ן~=���_K��ev�zt�'+T� )�~�nf>6A�Hh��G8mgzt�ĳq�}x?�ʬ�;커�Nz�X`Ҝ4C��'��`d��aL`"��З�� �B]�+�|8�{<��c�����3DT$]��H�[�w�C��ۊ�6?�؛ �!����	 �B ������v�%��mz�@��r��� ����ʘ̪$qȰA��kXH���z/��	q��O�CR���T�V��% ��{�4����3`��-�R��:VTa�¸VY�ۙyҨ��G�}������2!P0��ᴫw�I"�%�%/�>�5�=GĢ��l���w����$����#Ylȏ�[�T%p�K�^�Jé{ETܺ�6��6���ࡷ#M2�˓��ZFuQ;���~?4�; J�G!B����-,e1fY�1Vj�Pp�G��v�WG�����ap ����~��&
�Թ ����0�]�����	/�T6�WXx��7WK�Z}����8��֐qG��%�����)�w�( �Z��(����d��DV��h��
�>Uv|x��#�a����m��W#ֳ����O���N G�+��(�dB��k�!jז���j�?Z�-�ΏH����	���P�~��B�w8���P߮9��AW���w��V��q��Ւҗ,V�F*��2=�[13P�����z��BӱJ6!�#�0��
{�q(��V�+���t����r׳�nv�~1��
s�}�`�+8>�y���	6{f6Vm���8Y��7��_EH~ZޡQSJ+&��G���*��'k_�qm���Q����:ꑱ�ɝ�oP�Åk�!���8~���ex�Ӊ�zx�?0S���lf�.�[4���z���sU%�p���Md5U�b�#�"�#��� �)�,�)���:+A�ʓXQyH��۬���E#c�7�*�y�'R�̞��5�ߎm����Z�����@����u�z�&j��t��_<+Z��-��酸9K�����:�I�����Cr)U'~�������H� /�0<0�&* *xA|��C��H�a�~�ܹ��JS3�N��8�.҅�*g�xp)�1\N'�t�fqø�"��Y�r!������
� #��Vė�q�m8�im�TB�'���eJz��@���Y=��%�����g�H�1��C��R*�1�O�}�R��gמ�����g�۠#3r�f��K�k�J>����KS�Be��bp�"V���2e�T)1�~�sò�ps�'���p?������.I�&�g��Z��+FCB���oCK��dp�K�SO6��b�Ѩ��LS�$�\��խ`��"WBx+85���R)�~��7yc���m�4����	'������0�E�	I��-P��P���躱6IV��s&c?������U���2� Ӕ�z�H��wrS٬����Z�����&���\騩�q	��L3�l6��'�2r�In2�� ���l�}6������k����&@\��V��ތ}a�~E�~�$����|r�y�@��7�]�lx�U�g�!㽋��rKJ�V�Ho�Q�p6���������߰%c�lE]�!�IE3��ǳG���D$wˢG��T1�#O;s��#窄����C���xnʥz[��W���<+�T�A�n3e�[V�4�-LyA��t�ڗt�-�I6���D��1���#~���ޒ��5������:E+���Q�4C?�%01մcPa���Rd��j�I��� ��#����_�5AL���h39n'�m'���̅hU�r��Q�J���]�^5]ҫ�ӵy�ܷ�>Y��A�I�\���Z=�tl����S��"�����1V���	��Ur�/'�8T8�ox�O�Uo�B��V�g�0Ot�v�Fz�O�N-��yg}o1~���=0� ?�h�F~/.V[�=�.i`�k;�U��!X�kGǵ��-�����c')5�캥$-tK� ���$��PS��Vq����=¢�x����OC�$8���(�Թ��`��/�i}��u���"�+�+��S�!�Qøz�8���`��H( �����c8���V��R?w|��l���,c��}����S9c�T��ɢ4u���������[�t�v���9�=\ee�jd{�z~W�B'�!�Jv�������m�t(�j����R<F�;��D�	$zO	�!������w�E{݀��9QƁM/qnKNPp�2+_��~i�猿�H�ix��Q�吞^�bg�_��N*�	 ���f׬j6�tge��iu�v�r�S��T��<���`���DN5�t�n�N��x����:���U�e�wG#ƹ�����u[�Ec����T����达_?1f�y7WF �,�����2|��/d����S���@L�z0)<sGgϨ�a76���ÐQ�R�?_�oRs�z�J7a�D��%�	��M�^5�����ݏI����w��H�q�ª�O[��>$��i���Q�j���JXp�P�LH��_��v�|��{W�04����������ûg� D�1%�Ȟ��%�R-�|�ۯZ��$t���66���_0MtRg�����$9������g]�Q���*���e���6�̷c�+�x��ɋ4���m=g[ro�TXܪ~].���쌴�B����*�Ny�{��P-���_�Y�0	� \�G$!�ED��2�b��X��?�II�0��&�Z���p��!�)k�+G��y2�h�u��f��S�P������dSX�~�SE.d����K��7��r����Gn0؍`�캖K�*�te���݀��ؤi���)B�,D��W������}GH�a�������%$/��X�4	��-�����\t�Mc�C >r�>M_B����'2�vKX�P�3V���3�=t!�$���N��S���>���A�z&�X2ɳ0���e=>v�X����^�'��]�'�i�w!�)����	7��3
Ѭ9�0����WxnWΪ�֩8�..ҽ���V����'.�B��XYZ�65��J���GYϐ�`:.�}��!We<g�t���0?KdЍw�̩��6�G�MX��S�];�j,"F}�n����~��QV%U'a�	�E�p3�M��7�;9�����Z����:;�)O��"]n��j�Q��'+(�q�4��S!no�p��Ķ���
��ݺ�k�͡x������>s��������!�Kp&jb��:��L��K�P�C�'�pk$h �F����F:�$�rr8t�I�~!�u�	��J��8v�LO��Hή�.�h�,�K��dH���<����g�9�Z*d�]++խW��.�O�s�;��bqd�����{"�g�nc�����ԫG�~�w����W@��m���k�j�y#�aL��;�