��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�__I����Zw�
��Z6?pN��)gN0�dTrঽ,��0qqTi�m�s���W�g���m��?��ْb������1M����~������C����������r ��/�ݏ6�ƪ����_��T����V��"W��n
i��L��HG�<k�5Y2h0�/��쫅0K3�Tm +bC���|2��q@��9��_#�+��K�Td=O�ӎ<�[Bߛ�QK���� ]���tKn,�v����͜�jq�n+�O���V,uYA�X\��!��SZ�NhH�{�/A����?�u'�k�/�!+e7�ÖAI�|����
��:�I�����`=#sV�H-3N���(ʶY\G��;"iT�A���v�q��L��
�CEӊ.�B�=�l��(x������{�b�[1hFW�~$��3����쨰¾L>yG��ߝ�|W�(���Aq���=��Fe���^��3.�@��Z)�۫��ާ pggz1s&�B%��~E,��<Y��d1�`/���WF܋�{
�Y$�Ҁe���(f���RKɵ�e�3x�.b���~�ġu(�S�2]w�xo��z�jn�"�S�.�Yj(1'��[�� �ool����7����܂=�� +:�La�Il{]�S�7f ' ��h���;5�H�yy�tj_W���Ox �\�5����żL�gD�K��yM� ���5�\����!�
�����p�ʴ���MrD@�	��I�@��IP�C)�E���-l���p����	Lǵ���~����Ceģ���#��?�E�7��/�!r)2$�!��a{�m���g�=�=9m�#�$�od�®�ʕ�T�}&���Hv�@a��rb*H�~�Ѽ��L�lyTc�ĥ�Ï��i\w�a�!(*h�d�Z�7�e�V����l�>]]�����\>����'���p�&�ho{<g@����9�y����2_�A$̋4D������2�HL���:���1f�":7;B�Ӗ��w��k���<�c�� �M�1�V@�&���{7�#ﻕ�������e6gM�#��Vy��I
c�/߻����²޻ �N!JV>�'�v�R0ٿyá�e<b�����*[C	v��r'�*,�7�K�m?=��T��a~��hK�Ve����A�Y�|���؄�U)�Z[�vc����l#��G�r���]kKJ���+��'&<^~k������������l�����ꭳ��mP�s�I="t_�]8�紌�����;��#�}4~!ZԀ�l&^(�9�qTi��ʂ*��Tx�}�$����a�����̏OL�B��]�����u��A�z�]3T��xm�*�0�Qd�r{��ݕU-�����p�{�^ǀ����Pj��vv�\W[(n)��n)Б%G�XaaIY���KS�05}�/n�~�4�tn1���x����u�QT�vY�����Z�4�K��>��
�ͺѣ���uuٻI���ϓ}a&)�A&���=5����i�d�ZaL�ѽnӪ��:vK7O!<�����1-)4;9��7�T�E��>��Y�r���#�0"�Fp�g1?����?�R�ƥ�;�D�W+�#&i��!��N�P�Y��$\�����4}��쇇ZIA)F�A1Z�(eQ�œ�4>������8lD�t3��ۖf�Ѱg�����C�#@�R��Xw@��	�W�w����F���Y�$3F���j�����!bL�ڕx]ɖ����4l�U��F�y%��{��}�l���Z6��̞P��4k�q�P�q�r aIz�/y��qL�#��C��Dw��-8�#����'�]�(iB'�ܵ��B}��"f\%<7�3ځ*�P|ʁ�b2���F��.ZI;\l���^��Io��*4���;.Z��o��)�	�� .�c,�F�lߣ�h����u��d�^8M�2K�%~��{�yh�n�Rw�Mׯ2͆J	:�6n=�������D0���\AYOŹ��@Q�����K��k�:M#�\-��y:�u�JD�ȂB�E	�A��-�@�?h ���%|G\r�'���"�Jo�����a��d*|�Y �W���=��!+��0Ơ�!U�t�x��لvL��GZ�<�+&�N��"
���4�.�w������v|o/'V������t�m-�Y54`����Э�V�:N
�Q��q��eh��� u,�it�	���(����tP���է�suU�	��!���{�Q'���Yay�Ê�F D㣸l������Ɉ�3�O��n���sL)b�K,���iJ{���ȜrW�G�I��ԋ�>ۢ��}�����A�[8�	��F@!�7B)�ʱ���v��Vn�e��àj�H�nF�yh�}	�=�����B�*�޻أ(��j��ȓh.�����R����F��	D�ڦ Q�InV�N��-N����A>>�^b�Nz������u��!�1ϝ�ML�*��wg��Y��'�(������mS���]S�qu��U��i&�����Ybw#�@�U�}���w�>�J�xl�N�n���o�f�O�Yk�Ŗ�;3b���Q���y<�9^e�{h��ڵ�;�Dd�i��B���k ��ɍd_������ !��j�ch�-%=��xO��&��n���:��Rk\t�K�>O����y��pp���:Q��Xp��\�D�li��&�^����k{��!g�l���t�>��V�62�e ����KS����$��nW,@=~�ŵ/[���t��1�s�P��(_��Ŧ)|k����R���s|�H�������-u�t�M��d$Qg�� X�_�%�M���'l��,<�҅[�}�`���&8��c]qU�����Ta�vp��CC�1�Z|����@������R�9��=�2��K���1i���4?*�'�3	o��'�t�b�M�4�u%�A]T���Kv�q|l����aK_^�R�Fw�QB�J�)<[�x?�v#}/�#�X^�Z�Y+�SJO�c�ق?l���A:y�ǘ5���4����p�mJ�un�%��*���B/0�&մDɽ�}�
s~��b��0�W��2l�w�KL��x��gة(�)��3G�Y�Q9���vY�w���3�s+�s,/���(j��9�8?}$�'b�r���У�H�i��P�I����o�D ~lF�y�v5��C��l0�ac=��mʍ�
o�%�(D�lf�!fĢ&U�=sb;9�$l�
�����?�k�L��++x{���4�����Q��ܾ3��裊���ך���Xqn��ip��>#�!��yh�� ��%�iz�6"���/�C��/$]}����_ȸ��@ =�SƁ�BY�'�(��֎�/f3YAE�DCտ?�4�I��񎉭6������S	Y��n���,���+ 7Z͋�����.�-��n���i�4Q�6D���C���w��X�RKyM�BCH���G�X7b.�s��2^?�������gl��������[��L�t�� Nd�;���0 ��J-҈ѼR�=o �o�Í��`vz�2|p��q��K�n�G�f��m9_��c2���
�N�yKId�:���:���Y���Xu�O�m�xm�o���=]z�:] �����b�T�F�s��"א?�)1������.Y�C��:bs�R���� �9ʱD_/i��*���1��b'��۳�ˬ> ����αߖ�'-,�dXӟoo�OD%ۏ=g��{"�'S����*'�}��r���V	�b�w_�/%v��)Y;�.�U�	A��Ko��-�gp�Y�r&v�p�q�&�A�H�E�<�����a��f��Js��c�q6DO-<�9����.e���t�����W�,�X��XRj�q��lS�:;��-�рs�a�������J6 ���Ӱ�v�E�`�����۔�(m���O���{0��(:� �����2v�hq/V��#/Mt��'�"�
XN8��4:���y)�Œ��fr4��t�ݽ6B�t�r$e>0��.-(���#N/yP��s��c��4L2e�בp���3g�٘綾E����.e'I(�WIIbӕn�dS���"�}�#��Y���n;f}/ӥҩ7�l�k�|!7����e�6�Xǎ�o�Ш\fԡ�$��;��c^ʲ��S/�&����
���H�b?���䭤�F�dh�i��&2ZS�g/E)��=F*J�D�,K�����f9��X{�M/�NlZ֊������� ��S6��V��i� �&F�c�m��2�q5ӵ�ϱkCø�z�;���k�������\��?��7�Cd��U\<�
2i�����4�0Fƞ˺b�6�D�s����_��ݺ�����d�UTQ�:j�E�G&v"%���Q�ePEy�d������Zo���;� &r�@�F�K���:KB�aT��f�>�7%$��s�~�\`Y�{�̀�f�+c�o�MN*O�d R�2��TC� �U��.[k�{B� q���s�B%���d�]jSV�b���f9�����z�O��J�P[j^
[�̝c�WР�I���]x_O�����O/r$���-^�M��}Y� �|	��l��-c��_W	�R�K.oBdz`JK<\��9�h�O����"`����ևx��-EHU�J#z]ױ���nb����j��s4�4��9�ܘ�}C�Ftu�b�`L��4�6V&)��n"�;>����w�Kπ�a�f�Q�}��T�p���S�E�J���$���R8"O8�4�9PJX^&s�������6k�$Lj�L2q�. ��M�4�A�|�)^V;}�!%#����������d������2XSPW����.z4GnJK�	�fc�Ɨ�v���D1���ߎc����<��� j1�v|IY��I��w���䖉[jw/��dء(�s�	�&^��C���+�G�q0\��Wu���[�L�P�4˪!z�mU��KC�LJAǠ}�EO��sk���	*�"� ��x�䥳�ݦ�5�����/�_��`0ZN�5T�����s�W��
��;y��q�����fG����M��y�V�~Rq�j��Q��?�<��Q�J�|_�Y��	�NU��R����g����toב��N��_�:ဪ�N����?`ǚ+�<�����һ���rݓ�u�����x���6���V��0V�:�(�h@�]��AEU�i��F+�z:Ov��g�EX_1%"Z�����~X6b����z<���b�nX�w���Ī2�)aC���yg'�<�G{�
���M)�FJ(]qibp�P�S�Sm61+e�v*��׮�ekg������
2Ydұ�Ќr=���׌�&GjG�zC���.Ű��	}��� ���I�(�>y�u�V�Pß�h�����Q��d���l�E�'�K3�T�2�%5ų��Ԍ�<L�{���u����K�,��]�ej����[�aU�eϏ�&���n�oHx�d!g!������[CG��B/@��5(��,�J�?�|w�9ŻT�#`Xqӝa����H�<��f�����HQ�KC��JA� �&��t��6�d��ä��!�3�䲺�@)�-st�)��*tHܕ�|*n�'!}(��Pa�1�[u����7U�s��O�9r
���"@���5)��.,�luE괫�X1ps�a��M���K._ʽЀB��M�33d� m��m�2��������#ʝ݋��(HjM!�����.�}�	㻔�|pe��y	m�j+0z:=ѯij$�&J��ۂ��Yˑ�P���g�b�b(� /���`URNl��bSSD~��%�h�'Ɛ�� 3*��|�qv�̢9�}�M"Hj��ϖ��)Z\��s���(w9	�85��h�PB��1���N:����!��4p,�X\8c�y	��ޮ�Մ�V��/�L($a���y;���d�_Ui�!1�ۿ�=���b��h�b����T����H�M�a���z2Q��g�$��ʅm������p��Xf/�f%RƆ܈4��V$�0����\ ��>f�~ߨ��Y��_�o�|�a�e�p�@�6�z <�,*aA�X��}w��gd��a�s�:!�YZ����� �8��!d��dK儶��rB�z"��T��b�����7<�%���U3����R�Z�kO�T����d�.eJ������x�pI�w�j����r��pk`ѱ�_iu��\���W0�_�<h�Hx=	N�xf�dH���=ךH`+�{pQU��J��4��K0�^�6}��@�44�:���QZ��ٚ���8ʭ޹�2"�Rl�2N��x��:W� ����L�vDV���&Oם������ʊʖ��)���d�����ά��cT#P��������X7�_�]�.�Sv�j�ע���L��C�����cx$ݦ>���Y;�Lk8�pa#(w�H�󸻟�Tߧ��zYi7�cё-�$V���T�z����LnS�·E��i�ɷ@e�0ݵN�t>)f�]"�'�šZMxS$ٝ'��M��0����h�|�D�ȸ�v[d�W����{��8�,���W�8«�U�� �+G�P �^h}r�J�6��gmFf��:6�-�'�y��D� �)ͮ�D������e�3��Rۻ4�oW����VÃt���}��sb���� ��NJn��2)���u�)TʖB�*��մ<)�﮻���u{�JR�����s�Ӎb�.,�Y�j�\Н:����a��OWW�t�Ĕ�����~"G(t��k��vb�z�n�6�q�=,�C�]��&L�	�~��{{:`Hd�-d�_C����D�9�!�4���0�C
���h������umȡ�7���Gg�&��D48�:3#O�vQ[���Nw��!��O��gY�9�q��u��
�1������}SQ5��Uk�b����jK&�Q�� r� p�D�
�F�_0�@���$U�����_��k�X��HJ�WVF98�<����޳E�~��?���L�}��J�=�]'��^m`��J�o��(����R2Ɔ�IѡPe.��	��0�Dc��왮�R[���N+o�8"n�!Oaq���>�ݼY��p�u�<�욼��kLC�C������H~q�
="n,��5�������@�o�Yy��]l���};����w4k�j/xC_�T�����y�m?CmUGE�J��g��8�4(�Iei�R:��;?l��b�A��:�}fLAa*f��.�Dcgu�\~m"���Mo��sZ��=حդ��s���L�?�$�빭�%#���m��C��[~�z����xji�	�қF�0��e��z}C�m㻳7���z�!*���{(�4��PIeMqt�+�����D%���놱��{�%Q1� ��A��#������neB9�P|3Ց�X��������ro��~������9s���+H�E���WEln�	���P{d�;%5>��1 ��d��Y���1꒛���5�<T^��M�	�M�e�/�\x�n���^�D?�ҧw�D�\<H_�X��+}c�/ ���e�ŕ��ˎ��^�
X~��'��������W�XE{HG�cH���ڧ�`{ȷ/���j6Ǒ�����IMkM"�s�3����!E�Ҥ5d��T��V�[ź��v��I"v���)s�m�6�4�oSVA.C>�K�=�n���69��~�v���Oa�| Z�h��i����c���f�{`{��;�3���'z�9z���xڥ>��_X��v�U����9�өzh{��@&^��3�f�ɆH%���&nϧ���ے�zw�P�&�r#d��c�%(��e�I�>r�d�|'���<\�4�?��j��={mL�ϷO��lZMji��)iL�Kt�5W��c���v9�o^ĦL�fE�4�~�<�C�%���*�F��ѕJ�#����8�5sp<����w��`��Ug�y�K�/0���ϕS����ٯ���"��5A�ݓ������au&��I��((�g�s��!�<�,)����B��������'ߦ#C	KףHÃ���)��i+�W�j^�x�#$�@×������j�D��D_���wZ'��� ����DK|�=˕���*���[7n�U���o��E�)�%$oleYWdH�*�hҞ�]X���K^�������|�7�*��ʾ9�>p �a�36��߂T�>%�`��d� _Y�x����j��Ĵ{f�(���7tM��ܥ��aW�B�5�}�w9��@$�s�d�Z�ø��Q�]ĕ�}�`�v���W�y!��+��cŔo�$l�yꦾ��1��,s�Eh��Vf	� jV;�h��bn}�J��b�ڎ����v�b��N���]�TO�Ї�p�Q$Yx��x�+z�����I�4�!(��
�Ab��b2S��L#�}�\������-�P��dB�7ʞ��ƓY
��V��#��}b�W��G�)N��]kS�A�Ԋ�*n�.��<z�,NYG���)�J�[o���W<��+Ĳ闔m��>��l*U�I�x��Z�}G�c��{�����Q=1�u�5�USs�a���&��cॷ_3��8��H�$zY*�K-�&����0;Km��ƈ{*;*S��ۥ���th�T܏o\�	uR�l��R�_LSD�]�x%��
�k�-@#t�^�T߿�Lڃ�����Y��xfT�wX�s:�V�*����L���K���L*F��X���킚 �%$aGշ8f\���l>�~�P+��]R^>5�|,p�YL(|b�0n`?ޘ^*�ce����0P��<|h�W*�����^5�l}gK8�`M�V��1`(��c�; Z{%	�#7�+�&vYa�9f3�����.^
e� ec٪�^T?K4�P�	�S?DX�9��'ݪ��l+V��[hOL蠙M��ɣ$���=X�ɪ�P�rwzf�S�v�=�:v��c.E�%PB�����S��V�A+����,]`�%�ն���y(KG+mq3>��vE��B
�����{i�-샵�U��w \ԉ����#n�m͐�t�{(ͼ`1/�ռ�G7�A�kP�)YI�zh�s�׷1l��B>�1���Tߗ-�K5:0�`�����҆{�V_l�r�t��Y�Vy�H M�1�`2%џ>Q�$r����bd��}o#���C� B׫ȧ��m��Um��u͢66�X�\8]����DM ��O ���H��м*�an��8�r���s�]�[4�2!^�C���ƅ�]�ݴ����
���--����7{>�]�@>�p�d��i�&J�x>{�|���|�[$kq��jFۥ/��.*��j���3�$����J��J���7�o��+�$+**��ܲֈ����J5���,j;�����t��˪H�_|@q}�}=_Xn�m%���"+�$�w����P־��C�4d������P��l�X��iu�S,}���2gm_��IU�̴����4
+5�Qh�8��W7��?���m�_ƅ�A�!�K9A�u(M�o�!�����T�c��
wP'���HD�C���v�1�nSo{:s�2�"��eV}kD�_j���h����&1	�I<�ݒO��K�v4���9*�ʼ�Ƴ2�T�0�Ek�N�2,���|�u�9|�Ȯ�jZ��d�bqO����]R����Cѡ�t�ga{˯�% �&ע�K�8n�]��G��f*	�HU��F�ؑ�w�rZ�=5?t�5�^6�%�n$��Yb(;KI�E4�@�͑��Bn@���m8���!ƣf�+�0�p�y{��ڒ#v7qJR�E��z����]�i���O�fՇ6>k��oR����L�³��q�wT��2iCx�L�ݫ��~߄��e��ʐ�J!�&�a��s^Ġ��D]�X�.·y$\�eBE>��<�5�hx���Ucʛ?Q�lZ|��Y�`��43V<��ZP��_X`��&��H�a��R3e�jҵPc=M�'v���K��݄�e[��7�5��F�����cګ���: rFlާ�7�v���{^���3��H����1��Zȟ�՜o�Ss�����o�bVK�V�S�^��7g����+*! �P:p�"a��vjY=m����M���p�)��#�2��=�^��EN�t�H�.���i��e��֠��i��t����
G�oc�DqtZ�e�tE��\�`�5|m��V%G�E�w,4u�P>ǭ���t�
ݞ�uk�}�k-�Y�Q���,eub����T��~9���am�̈́���`\7��pav�O�{���r��q�����6!h�hT��:1�h���E��"��f�~qX�m-��~�O�O�_���w��v����V>��W*nz�R�&�#G]�8�e6�z�I停==9�iN�ts�=�#r�ǽiы�ւM0E��8��b�K>h<e���h1IP��Y�y]O�J�����OX�aB�S"������Z0��W��Yt,�ʌ�QD�e9�?7ỼM&���M_5�Q�'Mi��nbM1���J`�>��ʙ�G��ӕ��D�?����Kɹ����_Sb��,���m�.8hD�R�}���[�U>�k�F� �5�|?�y�\:����,􊇩9�gǭUq���Ja�HN@c,11�,Q=�bsM���� �A��记n%��@���Ֆ�12<�Or�T��T��!�WAH%P����QKe<��33�B����!�u}�
����ܖlف�"괽�Nx��a�o�#�߯�ip$sEb�aӨ��mv�H���	�D�S��F�C��y����\ t���>M����$�{���{�_�?c�(�^�O ��2�噜��X��a�J��O�P����2�c��!��͐$��f>��®�b%vn�pG�{���0���`j�����@�e6E�B��o�rt�#�^ ���`#�Qj<���W�>�.m�i��ܨ���w�z m�O��ǖ�����r��X�	���c��K�P�����͟%Џ:3���0}a]��Ke�+p���r].�A�ϭ�Vd�PcPW���C�QD��.\�9D�+y:$n��rŰ\�s�a9QK5*�t�����m=����:� @�>��l��&Z�����Ma�#H��n��X��h�%��T8'��9�+������-�������_���!�{TRs�}��5}q�a��0YP������tn��%�2�KKK�=������A���ZA��y�={σ�U���D��sC\|��g�+[����L�29��f���6|V�`�t�Ъ�E�v���dϸ#��[F�B�3�}5(�SJ���?���FM��ZV!r�{m��h��4��$�ڗ]��N�sx��<,f-�涝��z[����t߶�m�5s׻�����4/]M��~����hP����BU/[[�b�A�����@��-���p�r�1���Aȼ��ٽu�CR�<�y��ߛ�ָM.`�pR�0�v+��u�2)q���@��e��<����W������:��J�s��-�	aY�4�p`L��Ҷ�2��b9 ��XUKiƧ(D���L�7I�z@#]^�	�N� ��~ +9��a0�0����xn�
������B>�k�|�0��6��kQMx&�H�
�N�f�q�����1��|�I�V�xU��`Sɡ����u�w"�7C�ŧ�,�Շ$�^�в��M�Ia;X�{'���fv���B�(Lw_���b���X��y�u�P�w��ZM��-�R�Y���bL��o��z?S$|8p�+��(O�Ū��*�A�K1�I�����^{H�YXep>W��yXUI����ar��UUQ�����\�^D��!�_����f]ë�MΑ
ΉU�!�|��tĞR��� ���v2�0#���[(�{�XWe��+Q�~C�h�KゖEV���N����2�FW��K+`��Ss���t#���ofm�o�;c&O��E)9�a��ՕL�r���%m���Ѧ�I��_��s@7����X\Gj��*sٝ0tJ�ʏM��Љ��{4.�w1�YM�^���h-�0�71sF�"A<��R�v�&����rjQ<�� n����b(�X߬�f<�w��?F�-�pnY^/�o}����'S̵�b&h*l��"<�_��Q)�_(�K��zCm���i��0����z=3 �d(��
��'��e�i�W5�)�=77�
f`��3x�&
���F��J��gC!UHV�F����ڜf��{���8��*��
9F�l����piK��y#.fgy](\r�r�TLQ�+WPhg� �0�� Yɚ`R��''`p)VL�uMӝ+�e�y�Z�Y�[ka�3�+Z�8̎�ZK���n�������J�<s�Y�o�j��0�k@����8n���rD��|&���y�u�q��O-D՚�S�٫.�5�wF^|1Ķ�Ȯ]7d�  �������������=-�S���zb�#���IU4�n�W,e�x�N�g�Zݓ�f�P��ǘE�ɣ�� P%�P�?�� ����ı��2!n�����x�<��谦���}�,��{l��^�$�¾G�ri��G��D-��7��N��V�	6��w
Z��H�
K�H0E�)W�Hk4v0��������)��	��>�ئ �:�Ar�T�W��r=�cVm�!w�ڱ�dQ0eK`R6`d�\���d�E�ϒ_����5��`[�坯qb�z0�j��w�.Z(�5��2fkk�Ī���t�bҊ�� D�e���r�Ni�0��x�2%����JaE*���D�,�D��QǲSx�%'Ho$��Vkw�!�y���C��4��{*�%�����~\���VZ|收�"�(4���h����N�[#M�|�ҽz�%�w8�1a�p�U���>��TL�x�Z�)Xb��/�F��l�do�/��}�B��a.6�#�*�T*��E���I�9��
'AN��:w<G�ږ�d�P��T*&J�K$x�0�o��!������x���z ��T�[�Z���2W�BX�&��6C���K7���\hEI4����Gb�w,��̢��ή����?���޻T�јQ��O��n��M�:�T Y留L��>D"��6B��z��"�7���,y��	�R����Ɖ+_����pW�f��ˏ��J�E�"�Q�w�$*��X�2�Q�i4L)*�x�8	BO�[tP��]�a��-�Di�+Uo�N`5����h*�P�^@ɏ�jRMC����$���l�������V�a�W*�`�O�󑶐=�9ʔEp���Ojq =��oO�0�* 7�ڸ u����c���"�w�iʤ:#���csC}�b3l�0�����\Vg���g��t�O�����y?��P�Q�Az��