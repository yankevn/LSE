��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖw����$�OkA����.�⍁�cWg�J���>�eI
/��%��G�~�g&ØtW����t⿞.��� ˙!�q���Ch;�IF�N.��.I�u9*����㱽�q����6�c(*;q^XՉ�n@F�FM�Y9Ȩ�����JS}��� ���X�u󞍄���7hw{M��_�{��Eʛ�R�L}%����O./!G�ǯ>!�X�7��O�����A�9d��î�a�_���X��Y�-h"�����۳�¼���2�_�i0$(\��B%gX��jѻ��=��.xz'��:@�@"G�@�M��)�wQ(�"�q�$���f|�}�?"j��cN�{�n�T߽���K�n���ӟ��)���::�I�B��@�)qɩ�z�c�����>ح �Ug��L���������x�g� q��@@��Y�|�ZHQʼr�Q��t9�w^7�-�)5� ŭP���!��8 �Æ�?o��֧����#;ȧ�:���4�s�9>�[$�N������}�<v��ksu~�x�,T�P�1��L!��ߩ�
\���/�'�����q���^S��q�<��N�,�b�̂�-B<�	*������K�f���aD��{��o��e�s�!I���Oό�(����F�D2��R0r��Ce텘���`�{�W�B��E�《�%U����\�'}	�+�A<|����!�omU�4��!\���⣿�K%�$�F��[�7�j�T��S��+\�������#�Fŭ'��%����8�;��J��g�Ӡ�u���t�*.{�����SBIjA���
Ls���0�h���n����k�l�6}�n�?Gh�0Wq9��65�o|
�����7�:�!rΕ�w/��.��U�C�����⢯��ys��=ա��0��MCZL�`_gU���Ƒk�J���C%jf�u�٠�H�#�2�{�!#��_q��
���ѭ-�h�2���ﻥ@������P�M�ܻ�Jr[�#�z���y,F@�V'��EI�������l�p��P�n�D#e�`��B�|������2�G
I��>O��K�A����v�f����������$�k��C�V���)���BE� S)�.�O�J.� Yx㡈$+@o�^�'�[�ϝ|Y疺y�o�x�R��~�86�thy��:���_��6��2�L�2C�TھB����8��o�e�d=6{�|�5fߖb�'l��J��ٕ�:�j=,)~����?8�o��U�lՖ�Hv��p����mv��8��)�)��f�_^�W���|�������5فP]H#���4P1l�!~���G=�Ȕ�����hM���7��[N8-I�E�iw�I�Qo1�ɇN�K�	:�e��>3�
Z��W���"���q$?_恿��Fw���@"��Ed�LS��,���%�>X����]}?�jj�td�5A�#s`>�o�����$��NB���a%��{uf~ѓ�ɫ�W!e<�/�N?�oH�V��?��$�cޑY���f�Sj[�.�a�JNK�y�gR�T�W�C�F(I븄��2�Qxhj0I�5���D�J��=��-�Y7`�����k�(�T_�j���	�h@� ���>5�s?-n#�YE����{�3���\���w��-��T�ݤ5�t)k�I�ɫeb�gϤ�"��vtE�6h.8�l��+���`ʃ'�A���� ��.����+�Y��>���C����|)��/�LT㌺�2��)���']f�obu�$�tJ|��jc }!!ɢA���é"��x�4S��u �πex�0C��r��v�J���e'�gV�N՞9˩"K�?�\iA��z�t<��Ǫ�u:�̆.ݴ1d�Rx�������i��}@
�%[H�<��!��?f�����}EW��W]�fB��>>sl��sK��ќy7�Ϡ��'�
h2� 0cLU_��ljG�"��+�6:�0���8���'{��%���������z�(�%/�Y� �#!4ԉR7TZ�����׾�sh���
��I�_������w�l4���h�$����Ǉ"jU�;_T!,�y'��@w��׳��)��Z�FUZ�.�=���*oXG���<Ǩ�5��ұ�Ӌ!:	�^��b�|��(d@�?+W`��R�V����ês֡Ҧ%Kk$��_����fA��_�V:u(	H=e�;�����}T�h#>PO�O�`��9y��[���tF���s�
�׻ݵ'36'fWZnR�#>4�1�+T 8��=$���纛qhD#����B�$�c����!�̛���QR҄�BS�6�����Y�F/�KJ�<��8��lѹ��YvT�|aq}N��ݱ��}�hx�8.����� �����f&h�Ӯ����B�g
D�^�S�b����t�,N~Olյ�yIve���
�h���l�L�(ށ�Pw��Ktjq�C�S25~[���_�(��,�3�D��]�����=����{Y�nB���Snx�Cx
6��Bb���G.Y�np?���R�*9��}�8ټ�yRǺ$�Gq��L���_M8�����	LD�16'k*�߻�RI.�a��1=�*�f�b��%< ~1O�/Rv�ŞG�)�I�4=�8�1!dB��DLu�����8���"�MW�F<'bJŔw��� �=�C���,�bGM%��hX�P(� 1gf�n�c���S���?��,&6�$�_�u���(>u�v퉨������ŗ�|��8���ʾa��>o�����ڈr0�C��c+���e'��\�%�82���p�O=�J�sKfd��Z�_:﹫��!s���2�ȴ_e��Vt��Sq�­ǲ���S� ��2A E�H*�\���[ھ֐W��k"Y�-�~��&;?�>���߅����3u��t߶XK�d�Ƽ�e
O�`�	$���Ѩ6�X{(�U{���9F�9�F�8T5(TQ}=�Ri(��T�e��2HȻ��hW�E�ӉK��蓃"
y9���D\���M�+���g_gn��UKÉ�!�!n����|�%�]�9AN�dځ��X���eU�B�.R���,��:�I4I52������}&�"o��SoD�lЈ��,����g��/��g�OrsQ_� ���
�f;���1���͸A�^����$/��9��y�#ެp�C��^���b�8Þ�����Pq�-�לJS�c5ì�E��1���į��A`<t�.颲i�m7�66��92ת%��ֻ�^v���7B�v��C����C9s�P�kQ�<d^t��� HE�z�!'�زg�6y',b���9���ھ]��I6F�f�R��8�|�d,h��Dry`&�y.5��jI��H�l-���}�4M��ǫ��F}�'64���&aZtem_���GY�s�=�u�����pK�%3���frE���m����X��>nQ.��P��f�P�ip��]���!9Y�ȱ�veዉ\�����{/��ğ��&�[3d��u�h�y�iR�fZ �G~C��	��Y?4��{�w�/}�Et�J�6�����x^�%rK�3|9V%���3q��H:�'Cn�_�N��t�7O�-T��	j��%�u<��s�e[����z>�n���1�5X�Pu���/r�Z\+Z�/U�V�d|�����.�E�ȬH�U��7�G��P��9��b�R
Po=���1wH>��li&�Z�X�Q$��l�