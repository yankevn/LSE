��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�\|�m�2X��L�JTz� W�o�8Fb�Q�5ʙw׮�7��o-Arc�P�k'�T�F�?��}&������9�1Kf�i:�$�Ϝ���/x��.������@Sk�e��bM�п2�v�%��^W��1�o��R�{T��Е�22��f8����~=�h3�������$���^�Cmg�r��A�8���]�Xw�IK��Dl�0�v�֭�4/;��h�����4
�;M2�X��~�Sk�d�ϵ>e��^pV󷉈0�mg-S�n��<��m�4�z��0�]�����"�������]ٺ�D��e�W�����v4@��F��B�U��fw��c�jmb*�ߖ*���U���W;*$>H��w���]��y�3��aI�8��0�k|���M��D)��GK��z��~�8��B����t����T�x�uQ-�d!�2�Gd{d�z�#IFzx�5����A6����Z�x�����I��ׄ˞1���������K��M&Ԯ\�=��c��6��p^�t�
��C՝�s�O�@�@�謅�"{.m�_�r!��/ע�L�6��o"s��BP�6"(W��AP!������r�y���@��5��5GV�� �p��e��䕩
�r!�'��m�O~�f��AG�-����a��!9W�%��\�2��N�ǝPZ�߅��8�[���`��[�P��dC	��#�ޙ�����������N\F�t�3d���Le=�yU0[;r��9�	S��J������p@�w._\"t|�.NG�C���`�' '�%9d,�9"�X�ifQ=v���$du�Y�)�r����MtG�jA?�K�yP�F"��͈��C�XЏ�\qA��Mvi�W��~ �">�����/�3�2,q\����	�����C�nw�����y�w7���*o��ku7�a�)`9X֦��(�НL�o���LI{���o�����vc�5�5����!��AK�ӛ���>���?ԪT�)�e��[q�=}���<�Y�oٯ�2��iK^n����r��4��U�WTκ&�Q6�����AcCr��I�����P�����d�u~���%�'E�`�[ � ��9*y���K��_g^�=w�FSa�7Z����bK^�)�3�@�#��w�X�6�@+�.��=�N7�k-�l�������X�u�m܊�����&��a�Mzx������~0hʵ��aIuV���獑`���  ��2]�K��{U�������Zz�;Y�E�d߷�HB���է�@"���e(\I��soK�埵S���t��V{6Ȣ�_u�6u�G~��j���#u���l�I��Oa_�A���u#]ܮ.���hc�`b��8mT����6�U��hb�H�v����̡��54���N Tt97u�Z2\*q��QQ%��r̼v(ݡ�޾'0X��:[9�r�������5�?�0�+s6e�uý��st�s���;$�D�U��9��C%�7��43����Y�����r�Z�2
 ���η����|���?j�Z�;[���a0�(�_������Φ'I5�a|�l�b�v!<��%�������n��-�s��ܝ�'�ٽ��d�C���M��e>��%���)�P6*��I����Q˴'IB)Wt�6U�;ap��?��N�VJ ���1lo��
�(]V���Zԗ�0̰,�
TV`B!9䣽�OZkF�ސ�\D$�(�m*����v��.�FL���Ã���e�0�p�E��J�lY�n%f0j�<�P�_E���{��lt�+�f��Ļ2�X_����&0�g6b�)�lLK|ɻ_H��V褯���+�x; �|�"r�"-�)�r��2�%B�)��/����8Wɏ���7/�-�E�������)�t�����!���me��L��1�����&����P��S��ۻ�����ZI}�I��wt�5�����싻�l��$��Fz�	�����щ��_��s���H���%rN&j�~gm������6@��IO$��:�۪.����6��'X�kF��ꥫN2�o�ȃ3�:|�I*n�#S�U ����6=��'�;����0�N$?��A���A�^�0�w�n�qu���s(�Ը�H���u YH>�	=䁣~����dF��u*�����m�uH���XC&� �Th"VD��I�\��(��f�n��8�)��?ǥb*i�������0�>��Z�����u��&��ҫ���쉻&a<��9�G��mL� � �\0�d�UҌ"���BmR��Es'�v�o�u��A��3*a�X��7�{��O� >9��Y��������n[�s-Kt��񹜜SX�/�q�߰g;�n�X>�����(hl���Tl��ږ?�+2�TǍ��a�nԃt<�2bu�6_��grvx�}��=����,�w��5;�T����#�.�x�o��|>ɷEf��	h�Y�*���&�*�#�,�#�%͠-*F<3�O��Jbs܉M��Dj�=B�sS�u"�/��h����v��'9�5�[|��Qܙ>�-S�����o)�x����5\�A��nIwn�����X>������"�`g����9Ѧ�q���3�L�:x" �,�i��g)�7@U"�&h$����j�ic�`Ly�w��u1]��QHL8���I9�ĳ.r�KM�SF�Z���As/\�Qt'�Φ~S��`s\)��L����Zggҟ�T�pTO�cD���H�c�@e��4�g11�W�vG�����X����C["ذ���k_m�ˊ���(��^��Sѹ��)���T�NC���.6H�㐱XO���O��\��Rp�<oXf6�2ی���O3V��������Ƶ�N.7wt`�^��s1� ��X���'�j���`����2�=��FA��FNJ��q�%c\�t�`8���^��J�N[�UJ[�����<X�Yy������{���_�+�������%��<<?{]���6Nwa��m��_őW��|�VK��AY�ݷ���R�,~��ٌ��UY{���-_�g�ě|���<�%,�с��>�5���ۭO�ݲ�����J�}װ�9`���1so)˼J��s~Ɩ1���-�:�F�d�$���"e=�!xQ�Z���8<����d`2��ME9�1}�w�ȭ�H�
�m�Ð���m\ӈ�Y���o�Uu5Z�wւ��=� :}�g��tu�P��Բ�{�ʹO�<L��N`���"m�ԣD7%.��q�G�Q~�4�z`�X�5X��+�{(�w�f��� ���C�]���bn���rv��������c�(/a��u���W{�Γ�D��jm���Y�rj����6�Df���gP�4w�t�V�w��H�b��ȼ�-�󸂒�-]ϼ�:� �1��*�q`��ݵ����i�c���������E_��j9�4%b�n$-��0�*>�����F��r��m_y����B��]�·c���>p(:�����}����F�b�Up�����}\y��V	��u���8�="~�<O,��kQH�a B��GQ9�A��kẤ���^[Uf�J�5���T6���'���'���h�V*��PC�Cu�M;�-�� A����M�J �ߤ�	�1!���7��B���1�	+c� Y�����L���}�Rx�'��FB�y�a4
��5{/��ݒN$�����au��z��6�%KM���N���L�۹��=��������p��~�v����F�bܜu�=�~��lX���r�0t�]��������.��;Y�#ze�؜=��M�Ҁ@�-
�3���w�P0`���B�]����O�^!�����ϹR�:ϕK:}�.����c�3��\��[�|�����v2
����Gz�o��"J_��҈��E����Z)Q�'��szA��6|��A+�[���`��:?m&��]��ҩ���}#� �끚�S��I��G��f�s�$>�~@��k���PARo�m��'�?�B�Zm�Q��R��ӎ�Є�Z���{�� �]��RM�i��?}�oO*��&m���^tg=s̾�X��������t���S��	�\w�-���s���??l��2v*�Q;_;�Rγ��gX.PYh�g)�^(���6�%S��\���2ܸ�r�B�$�J�~*>)�hV��[� �z�p)7�&'�������SO����:�����D��ܪ
����$S� �J^��ֆ^7�~��֎8�B���&��%3�"q#R�֯L�O�|\�вb�>P�/;BU���G��?�; �&|
�1�g2�f)�	�G��gh�:~��:��:т��o�%�����bVⷾ�LE�1�4��R�\R�H7���@Q��:�����U)Rx�l��̡2�E�ۛl��h�Z�k��kW􏆲��ہ7��
"]#Z�e�B[v$J0���087����!�a��z' _[�x��yR��6j��z(�VY��-V�i;��}h�RJ�$[UH�:J���$�<�ވ�����2툴��{7���)�2��2�3=�M����ea՝��� �;q��#XͿ˿>j�4����\ʬL��`YF�اJ̑�M����q����A���2v��q$N6o�=`�F��TN�>�~�^YHaQ�^�1ɂ�ulp[	HݖR���]�T�U��==48N��΀�� i��V1�U����CB�?oեokR����za��;ſ�����
��4m#YB
�ڪ�$�����)����ʩ��gr���2���+&��6�1�}Xr�m��{�Z���G;�˚;qO���
\f
O?�o*c�/��o\�!;2��O%�4T����Hr��V���V��q)�F�M�U����L*^>���T�k*�=`bytmoW���1�B��"�f�+�����v-��G,����-�2�@&i�@k�`9���@�˫����v�:���[�
��s�]��I�^�qn��x�8 �yHY6�n�v$g��l��n���3템��I[WXd��DEQ
� #��+�E�?�!8�$��X�lN"&p����xX��u�{N����qr:q������v9�?�&ȷ%����5�Ɛ�!(�7aX�#*�j�#k�5����e����@Q�+!���������\�d��Uc-%��,�+J6�]KN�#�c��ۺ����W�B�(0�l�֮���D�o{	
\��^���=��oSuL�]
��r�)��v4�Í<?��_ ��ZϢ���Iy��Q��z�'��.��

�r�?RMz,K�iEM�Z̟,[��#V�Ut؂���G+Q�F)(�����)E���r0TvU�O��?C&=�i�`[��VĞ���`S4
.����Ҷ�X�?��B�[��\o��@��84�7g�pn�������1���H6tvghֆ��w@}ʉB?��ӕ試��A�/%[;�?'�^�Am.�ʍAH��~����
^�M��5��h�#�b�Kț�>'Pɐ� ␢w�͎�ąDٯbq�#�3��NU�5�<E���s��JV��I켄��o��{x,��ώ���J���-^࿜PՐo,
D�NA�c��E��ĵӐ��l��qc��,[@���=_�H|��<���H؄;v�*�>`��ꨛy�3g+���8/��.�D5��vy-Dꜝ>ҿ9ZX)_C��v�����rl������.���ypAT���_P���7
� .���ȋg�����yK;�����VlgpE�XА������ܢ��U��='ʙ(opŐ�;�n����/B멘{�.Czy�ҍ��hn[��� �W��һ)�Db������C���+Pi'��[�_�f�%��$�H�k"�\��ybW�c��cߨ,Ė�B�ѡ�����x�
mؙ�����M;y��QK���.a�͐W��79 -�������u.��N�ܔ��h �cgG��I�\����