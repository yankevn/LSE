��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv 6�$���m|9�μ��:q����H�r�4�A�����ls�w�"�E~���Z�ޣ��IS��K�l��ĜJp������2Q���{
����qˍ��|���e�����g�R��hG�"	�/��,+�J�=F	�k�@']K��lx`Bp�&c�Ux=����R9nG�r��\W� ɞl�b���~A�R�:�gI���ν:�a�81������E48�ԁy�G�^,u�����\�`DzZ��0��d���$7��,^�cN�w��ʜ���A"�:�r�|j��vz��Q��f����=&!�[��������;k�	��6�U�W^����E�p�D�� �[�@߳����
��yt*���`�u��ʊD�B��m���z��7H���6�[!{��"���@�;Y��IsK��c����X"�Ѱ Wa|)�{iG�==NW��
-�_�^�'���,� L���e|ݛ��lQH0@y|���v�Rf��{�?	�o�bp���K��d�ܑ�OH~��θ�-1��|���d�2GIߡ	[�X��d���G�J�W-��=�D0w�\����d��j8FȖ����@D8-so���t�-��Dά^�V/v�:ɼڼ�t��"a�(�R�f�?f�4��|�A���hU=��l���5`����$r����kH2����``	Gݏ�*�I=F�R��g�%�p!:�`r
������.S$\��E�Qh:>+"D��W����0��Mt"��+�8� �W��L-�U__M@�3� #�ow�L�.��� ���4V��[�d��wA��e��GP��vS��9B��к�`��jGk�OkT�[y����"��@���v\�͎yI�v���,�6�5C�"��#.EYQ�ۜZ�v��?{�"��ՙ�>/�ԁP����X�R��N�}��S�9���6����1$~g��;����s�t6�"���`~D�޸�y�4j�ɾ<̼ש �%�%gnX��f�M�Hۖ���47)l����J,�M!['� S~K���Î�XA�Q�İ�sjVP�������'ӛ���\MV^�RG��#�(9��Ĩ��n	��-4�NL5��@6���H�\�sP�( 5�M:�M<�GD-�L�JR����c\����<�g_�4ũ��`�Wz���4ź���[z2c���ae���_���7�>}���>�=�V��1��e4�FA����+�,!@�Ud)�c�����7�p�΁��@)�f:�ҳu��"1�ul;a+e��0��m��y(�\�����}iȍ���Y��S�P4�:��L���$��j�q�i�W��������>z�/HvQ�Ud!%�����1�zBP��d��0�ئ��oO<�GV��y������,�=������B)92]Z���9���=�@a�@�Rpș��F,|���vP���`���|�X �9�e��RnQrw ��F�	r̯X��<�a��f����)����+h���d
?g��Y�஦���wbΫ�=!��g�{d󾩝�6��'a��s�`������}�RڊF���v?��w��	�$�G���&,���&49�(LO�&�����:��Ny#�+?����$�H��"ǒ>�g�ጿt6����y�W.��_���QCI�8���M�byŔF!��bF�6�tu��Z�Ӡ+P&kY�dѬ(���ӕ�J���9E�r9>�س�M�s�ul���� �.�/�Ԓ�+���vӰ ���	qy�<�};
ʧ��.�_��ǤJ���I�ԋ{��q�vmڳ�8	N]8�c^;{��_C�g.��h������'��K���2�g�j2��q��f'!]�W+�9��>����i�0f3�?�]�]���6$b�0�h"s��ݘK`�'�fX"�릇k�	ةp~�bmʴ��ݙ�N_s��\����{�6a��e�Q��!�@T���zOW�����q�u$0��7��B�O#{�<5��-0��+�&�LR��9h��`+�k?����3n�n	_�#�
UP���w�|�f��֮
T:[5�L�a�Ԗ�
��v����K�?��0ؐ岷�6e#��$�5X"�OrV����M�h�y[-�<�
L�J��u����/�$D���Q�09
�fӋa��}��v�^��RT�,_���*����u�;lh����_tNډ�d*0:9-,EB�0�$��!W����'���Oi �J�>tx�w�}���ah�8��'�1�\n�k]����QI��$�\��3��u���r�N@�������CSF2!�!k� ]7����N�[�gg�4R�[p���ՠm��]�}!d܄��z�s������T����E� ݟ�"f���@}���YFGXG{`k|H��3��J.���q04�ì�O^��m��nκ����ܒ|���)a��%iMT���ބ%)t��!��3u�C�9yӨS��䕞Ɂ��&�5��o�xc�ʟ��d������%�S�4G͍�,���y���pN���M�ĸ�п,d��ºi�'�GH�# }�.�&��E�e�ݣG�A#k�b1c7�iUl���r�Rۇku%�vkz�_Sx�J��ޙ����P�l��C��R�H�h !��9�tϙ��4�/�]�<TmO4Q�y��z����}�p�%��щ*���C��7u>�qH�pR,��`�����[VGƸ����>c�R#�Z����9(��{'���}y2c��{c�Bs��eׯ�{�Va\���E���'\��Q0�o>���>r����}�M.xqo%�B�8��1�k����2�?�N�YP8w�Tz�*ۆ�:����t1���u��Hɣ��m�"�'�>� =�&{&��g����,�w�xG�f3���)v�D�]�`�	���c�?�	��M�*V�� f��e�?HTk�w��(�;2�����3cu1�D��K���3�o봫�+͠��p!�t��]�f���2ӕ���3��ŧv7~��V^J���,�C��~F�[�ƻ5/0{	�"���W��|>o��3�,f�������q�ſ�s�1Q�O�%a�j�N��c��hoyA{��b#�iw��͵�r�9�+;r�3@��46'�Ec�����O#����"�f?<L���m��	�Q�yP'����i�9X� }�J��P���ɯ������Ĩ���1�W1�=�j�o!�+��
m����[{�uF6�! .��]���%���*h-ۜ�ge�
q���W����t�N�0i��j>�,��/z�V"ƃ�� �	h|����2�F]����X����D7�-��r߀^�#e��5��D�8`U�`J%Ҥ��ܩ� ���%�zB۩a���M�6[r�����#]���Z4<���~C�1�p,���s�� �u�<Ј<�잪i�/	�坖Rl���5<7����q�Wa����{\(T��I��� %�%�/�9��5��&Cr�*�m��|͜:�&�	��n����ǧ~�DضC�T�/�Ğ�z�ط����y�E%�LżFpdr�U��(�Z[zT�̈́��EA:k.uxܲ�(^<Us�)����@�ǍmAB�>'a/0����nU*�'`��̒�Q�D� U6h�Ș�	��Y$l҉���[4�� l�D���H�sX-�{����Ŏ��M�[]ղ:b�!��u�zk	�k�\�{�o%<�ρ&*�?��a���ھ(g�(U?EK��cb���#omC��.�&�ݾ��u ��B-�Y�@�v�*&ya�?��b����6K?�	$z{�e��|�a\ +�R���86�f�߁l�>Z��)��}E�7<:��%���l5�� #g��H�ة3����2����Q�D.�!Ƃ�kx
�4~V�dAW��1�X����V��J*���5o{�߁]�vHK�Vgޞ��Û��F��d�Y Yg��t6!q�Ry ��Kzk���I��u��EG��rZ ���w!���k�)��<E�n���-�m���=/�@'{��D8���CT���䯢m�DdrW��z��C �ҿ�z/��˅Erҕ�Ot󎫲#��9�}8�����:�6��V��D�j�U˄��Gq�D��u�����<Q���'}�bM��io/����I��`�+H=b��:-��'Y �W-����
܌����ɹh��rb�]��nfr�nc�@Ӎ��q����xp�Hu�e�kEV]*%n�[���(���{�.a�/�
�~Ȗ�k�hrw������!��8��3G��d�2		%�@Lpy~�g�1�RC���"-��}N�?<��R)����������x����"�y���etx-Ѐ	X� ��@553��5)�N� \��0����ω�lѶ�����y��HΥ1�W�u�X/Ӿ3ָ�=�N	��^O
�B�sQ<����q�ax^qx��:ZB��#�6���%4穄����A��-`-�c�[4kt�碐yx�GىY�!e�s���WP�tX�ݷ�9Ӗ�d�Þ��Y�I�w@����B��p�\��S)��Yb+h�hTQ�z�J���a
a3�&��<�w�P��ێ���dH��(�|�B@>��m��
�;�a��']Һ�B�BCğk�_�J��8�(y�i6� h3���f9���3��`�e����v�^�HSO�?��_�;�E��M9uG3�d'��q��j*�ڵ��a'�u��"O�&%�����(X��Q�W84n��~�%� kJ�Z<1����Sx�P��TN
��OY�5}�L��y�r�JS]�RR����hm�A�	�}���4�T��g����9�m�J�����Oo��\�;���=����4�Y��*=��^�q��N���j/K�ږ�8Ku���AR9���&��VܥC�J�������ڈ��H[���aʨ[��mL=�0�Q��n6��7�#�3`�.PiD5ۃ�]Ŧ_!�c�gm3���.���A�1��J��X�*#��΅t�d�?���]u��a�CQ����{����������5�,�z��8r^7�*b�<�4�8|�%���>����>熪��;��R<�_a�MK	d=C^�d�9�2�����b'3u	S�'{l�S��.�����~�����xbE�r1>��ۻ�\��$�b�{m)M�n>���Ƚ�A��� $��+��@l��Y���P?���֑�P�]T,��r���Օ� 8�,���
s�کܠ#ލ�V��=;^g�b`bc��ǐs(�/����}�Z/�վ��G6Z�Ǭ`�)ʵ��r?��җ��5K;Y	�4y����@�������$&�5=�vJ/�u����HQ�zb5w"{Gc�%��ݺ�"\��]#���?-Z�0�����Z���ٞ���B��1kCf4q]�[oh����70�-��*�h�r���N�ih��n�ɻ�T�v��r�#��5���li��9ʾSa8�"~h�y{��H��@GYi$.a�\��vu"ա�����u������kED�i��YpﻭU���l��uc�h&M�*�9�/Kю������__���K�؄c?��ْ)������Sg<�w���6���/�ؔR�ڮ>�r�swP�K.~�	<��$�j�k��+���gWhEv��m��<Y�Zbv�u��2ev�h��r,%��-#�_�hF���|z�T�Q��{���(�$�Pm�Ru������H�l!y-��p�_���nM��'��C���-�2����?�.d�l�c��ºD�p]�h^S�Y���c�H��U�<�p	ta�l��j��u�ɿ�:�弸���p��|��o�|�*�(%����o+vI��Z$�eq_�*�4:R�{b!@u�ɘ8���9�Z�<p+�ZcƊ�*Ȳh�[`~�*��!�uU�I�5�>F��J�Gqe=�|g��*JZ���*<�󤕂F�é�wt��`TҐCj�|髧N~�mB�3�� �2Ň7M�A���rú��X _q�C���� "n1v�mW�oV���0w��5}�9s܍��\�RzS��LCQ�a���nb���{�.�Ҟ�g�b)�-����Ki��q��?d�5�@\�6��UL~��r���ayo��b^����[�*��
I�q�\�;��*$u�?���jQc'��;®������i:��$�(�p��U14��`@��A
����^)dpc� � V7sE�;�RQ�uV��_�;9�V��4������R���%��:T��W�4e��	\$�}VA�(_��,E�[Έu6&�*!���y���(���1����5J��}=�,���O��T�9O�B9=y=��A�
�|�+��P5}�InK�:+{��4���Y�E��^����ֿ�Q����[b�n�P�# ���F�Y����x�3�/��.��{�آ��N)QD����,�V�M�k�O$�[�26`T0�YY�k���v��C�8�u�������Z������J��Y9Z�E'�["�<�A����e�����Y��~<�ݻ�����^n���3� 9[SZB���c(U\�z�:;�X0BB�
Iu�1�ф�C��3Ħ)����PQ�W�w�]�C�e7o1�`ZZ�B����x�iX���G��"�%��7b��ȅ��?8s��.�*�G�H�CUX��rH��>���K���_}�� \d!�-�J��Q[����_`w�<���r�A�\T�f�X[9��e�����n��D�֞����t����R��j���(VRs㫡�]M36+m����	\u2s������uZZ.���ޮۺ{�0�����[� ����f�#3O�7Ɛl�s���!o��rf��U�M�ZE�g�9DPe�a���kQ�@�2�y_c9�_�nP(Eӿ!Y��>��b��T�;�Ѱ0�ԑ��z}��Kzv��b�Pju�DnVd�S��\���uW�:�-)DL��IR�B��/�5��=���M��F)-' c�UHd���������Iq���y����	�.}�ЪYNN5I�L2e9n�<���N�B8�\U���B/�(z�Yu�˝��ί� �O1�5�$z"��	X)ͧ�n��u��֢����Y`�:`�����8-{��ºگ:nJΞ�Oz$V0�9�@�� U�Fb�L�2x���ÛǏ8����k	ݙU�1	Ɂ��������(7濪�ѠE�",c����H��Bp�"����U	�v�&�z:b= �|�0��:���R��0ŵ|��
c��"��\�qu�Q}�X+_H�7������z��rD�����C���`\Ԕj�6����{#k�����[}��U�D�,�"m�-���d�
]���rF����E:կQ�B�{ofы�٠���⾵�w��+H�
W���<�*68Mܫ�[��.d��eiD?}e{�AC	�`3� 8��! ��|@��1��Gr��^�BI�	?���\$4`˳� d�D!e���iJ��6<
X��x�1b���7� �eR���K�Nט�H�0V����O��#  ECX��'��9�S̉u�G'���/�1rl�L0hp�v�	��Q�N��$��v|	�:s2{ �]�k|</1�X���{���>�2���(�&�5!��/��8��B�`]�^n���,I�^�$���ZE2-I#Xk	�3�qB��]�Q]O++va� �5�x7X}F-�8�DR������������a�7���вp��m��8��H����W�d�Q���$,�\](^^��p� ��x���g�y���y`ր���Sf_���.�#a���@e���0o� V�m�*��r�"]v��b��y���y��r��:�����.�������|de�F�5�俥z�N�R��/��K\t�Di�� ɫ7����-��qY=MǤж;�(s,��Q���:I&Ʌ���aH'S�������ى5뺯��R�i9�n��DrH��(5w��
T�v��A� �_�J|l�r�CP �.�jL��}�L���e�E��_6��;�՚��%�HI�x$�b�!A��$n�:��D�6��ߍ~�4~�Aa��]d�a?��9iyZZ�{�3<Ho��X�aIW�~̌��j�ߑlD���F	K`Ùq>X�o�@�a8����o�s{��I��CSs�݈�kQ�Y4��$�Z�?�zO�8���<��L���?��2e��C���VP6X�*�0�Շ�N��a8� �#�yփ|�̃�e�>n�5�_�M�n�RV7Jjurթ�>Y�5�^^١��s�k�n�!B&bsQ�%�m�Xd���2��5%��m����0.�����H��`���B�13W�1_=���ǜ��~�Q�f�5
d����X��:*ssS��nϜ�Eנ��-I"���D�:�����(� �t^�ڌ����ǯ���]�>�� �F���gH�����0WRc�g�}r�sFuO�Wx�M&H�m�P��<sNhGT����Y`l���VО�~&��=!.�^���jGcƖ���� |�J�����u�����4xϦo��X�:m;�ȗ�T�Q
� оwl�^�Q�^6��S)���ی�����LW>��,�~N<�#� )��@��6gO�@�!9\�ja���ޮ����mL�%�!�B��K�j��Ea�p+��eI�*5��gt!�?��0�j� �DV��-�Z�E�o�B� ��ZJ��9D��,n
h����K���6�R�>h�Ԫ�g@�Pw u�ѻ���nmp��yo��D��(t3^�vy��H�(�ld�N�q+��}�Lk��:��DǾj��=��|�r%�WE#�A�vۅ2k%�g1��-u&�X�%���?��. �}`����`� .�z$G\�g�NsI�7V���� ����/!��k��뮓�t��nꃣ6���	,ax� ��a��8f�ݑ���v,�u�Z=��JEŅ"�#�q�A�n��%�֙�_.������տ�>Բ�����c�.c��g�k�8ꗇM�%0L���w!V�«�9h��(�ҭp��ݞa<�R�86���Q�Gl��ߦ������K���k�w
-�J� (�����%s�0�V��4�0��!&�f۱Q�˰PC�D�Ԝ���Ȏ�dfT���k�ҒҎ���R�c|yA��"c�P��D���(;P��ʻ�~��
i���p8����A'�7z�|�43�����⨚�;|�e�6_�z�M�giG �����ϖt�LHt>4Y�X*�d�CՉ)�/e�bB��@�YM���F��z{��|��U�d�Uqo��5h�v��YLS���u��Yv��j�;��T�K���#a?��UV��l��g��_4��s�:�S�w�҅��ϋ����|���x�Y9��E��ƨ�k�����	�w�Icٸ%-��m ҽ�s��scO���������y��B���_Y��^�b�̞^�{TĜh����&!��8��pZ���E��7�ܨ��؇�}��d+��MN�.֓����7��*�a�]Ʌ��X��"���,��|����7�A����(~K�( ���<\?�.��dW2;fʔ�s��!�-���S�Y� ˨y,�ԝ�+"�U�y#y�!L�	+\��(�����>�ޖݸ����/����i��F�5��T�X�I�
f�4��I3Y�Z�_ܦ���@�8o�.6�8���e�OO�
�XJv��^��n�e�+@G��o*ȡ���H_S���-��6��/��9z�ȭk]�*!�ȼZ�>�����a��1�--�J.u ��@s����������<L����2�~JRMpo��U�bl�DS�IE}�P�1-2�C��+�:�~�@��
��&<>]�B�� X����i/�2Wo���t�k�޾?IA��=x`��� �v�w�w�橵;�aeR����ъ.F;�(i�s����Z�t[1:��F3���2oH��+q
��L���T��q>�a"�{=aYo3y�n�
ɺL�Cܿ��]Ѳ)��XN���� ؃���1��/ ��A?��$^����A���n�%ׇ�&$C��`dIe- ���Cن�X�q�Y7��l�ߵ{�^zƺ��o�X�_��oT�z��v���MX����iv��M^K�����w$��S?�7�ZP!etO�ϖ�i�}m��b͒��z�1���:G%�0C<�8�nY[�%$k�=x��I�_)�=s�e����8o�h��b�F��3s�4��
�Qj��H����o��_���}wX㉙V+���WH��ܻ��O.����-�iU���0o�`��$�:1N� ���^�A9����DJ��iZ���G�Ou�憔9u$��Zs1�6�A�m�?.��OղWČ�$�e�~.�G�W� �G�5�_���"���7���"<l���^P��� [���wo�SM�b!m�����	���dT63$��%˥,�
:��3�TN;�]�EQL"�e>�u�n\h���_�e�>��h%7��!�E�R�|NG�/C�L
{����G��0U�l�4��XSGD��.٣��B�Gw��3��[�:R����Z7���K���!�Յ�q���Tg�>��Z��瞽��>��M6$M�G�~��$%+c��3t�Eә��͹�J��͊�ҩ�%۾�l��c�}���|����pS9�8�9�mLq~	A�Jl���	�ni8�a1�|���[E$鹝��!���y܊���#k��S4v������Q�WW3�yт�O1�>�v�Bl����8����_�����Y� ǅq��QW9�*\��K��O���Y-���UUx�1G�%Β����h���$�;.�7%/���6�hl+e���`�$̬,k�m�����z�����S�E�Xx_�Q�k;�#��0�FnE�$�^# ���LR����*[�!�Ky��gl.���|]\.q X�<�5;y�Tp�j��r�>����G�7j3��ϰ�hӅ�Nє�S6Md��'�X���o���ƱH�A�w��.����\�f�H�r�$]��b�����,�l�4�vFie�M�~�52M��x��8�hpCCKlI&t�*	�(��h�⏧��� �#�mcN%�;����|v�bFc|�f�%;�Fgok���/V�L_;����Ct�"/�In�#:!,�_�v �͜��F�KmP��*@gۼ�_�1:�HU�]�[�S�֒CJ�@)C��1�f����-4�A��p�b��S�cx�Gz���As>KG����x!�m��4[�1��]�B�4��Ds9���<g٢��MXD��EJ� ���ȘM��*,aa����a�<�j�Y)��!�c��o2�o���rM sG���<s�q���YQ�f~|8@�{��i�e~`V��'�e3¹�d,�x�簪�?|۸��윤�^j����]f?nn�d��P��+��,�q8^<P�U�A����sbf�����P�%�@��l�*�ʍ���)�lbF'^��'g��p�)�]7#��x��l��Ѧ0�șxX��Zٞ���K�����-Wj�t�>�+�0ڙ��XIO�r�F�a���p�7�#�	#ѝ7\'�6�x�r�O2�F�oj�s��Ϥ�8-�����C��Į�p�-i�Mjk����n���@��yx"�{�ƍ&�䌖����~g�w`���7D�ʭ���֦Q�S'Ml %�
���Qr��k�B.:
��A c��.k�dm�,��zw����ըYtUd��~��9["9�uS��G�Z�%q���°��]�8A+�k�[�$�]/�9�6:�u��8�Xq4�<���
�yP(�.f��B�}5QNL�yNV<#����_�Sl����
��Gt���֋S-qأ&rCV�x�x�1�l�`�=��o�n����'�8�
������m�@ts��K8��H����������:�i���L�+�6D���3O6�%z}+�Zw6���T5�6�/�B���鈆�!$8�d%�e.�ǋ�!�%�UA)��o�\Z��m�+��O�xoW~\�'gY�0a��|��1ɝ���A�J��ŭ��:`�/�e)N����f�`D3^���y�(Q%��3�AW��i7�c���a>�|tx�0���5��G+Q�ʬ�%&&.��;n�@ڵ�VK7�D�B�,����bR�i\�u�QB�͎e�\d���o��n~#�)*)zҨ�H����������fvcY���u�Ϡ�A���@�*�ySw�o|�6D7�F���K���/f6W����x��P��ͅލwogq`��\|flI&[6��M�u���	<ذ��|ώT�(*�:�@\�j��ZEA������V�h�9
y�^iD_�p�4ᅳ���#���v�0��+���w�wV~�P�����v*����k}gw�Wk���l�*$D�w��x���<�j�g�^r,�'G��@-�
Bj�:WaEY�jp�����2��E�%fav�KΌ&ؗ�[+�"���D�-:~V���i�XT7��W$k�l��D�y#�;��m;r>I5xy�r��0�\a)	���Z��{��1im����G.��;��f��W!��"�Q���>�"{�?�=@�a������X�u�y�]k �.
�	~�kb���d|f!A�5��	�K@�6}�/6r)_�]��z��]E&��{�$�w 즯��M�Ԑ��Wq��$bg�՗BP�ǖ�t�r0�,���B�D$ ���#�@�����a};���ޒQ�����Y�_�o��)N�
9�[�NV�<>(�j�Ԑ���^g X�X��vꠝJ*���v��-���ڄBל��B9�G:Vj��]䅏`Wܧ<$h&k�@��=��;��N�^c'c)Q��om�����"؜`��:���)lӌ\�(�jje��W΅ܲW�6�����_Z�g�&�ؑ,]&P�#w��ںyV�A�P�kBh�����12�/��='+#�vS�5��qۻ�����D���l�r����5ۇ ���������9N��?*gjF#��3�c5��r�m������|�V�gd8��n����7���}�_׿U�띱�EA[=�%����FM�(���t��qW���!�� ґA�2������!$ߵ�kH3�/����֦��݈|Ō����D}�1֫�x�l��v}��l���1):�68���.zҎ�+i}�/���^�д�����h:�����C�a]�(*/AM����,8Q�e4�#��P���&�6.Nq�yƊX.�AԸ�ݶ0��>�qWκgTT�Ԝ(��c^��Rj�|�ֹ�e�'B4h�x*t�ϊ�HFk-8����2A&�讞��
$*�a�!�C�������(�S�(��w�$M�.v��(�~��Y�1�� u8��&9a�8o8�KP�+Ա�b�!š�����Gw#��oma�0��#��f{e;le����§��#��]����j롆[}aP�_�̧�3.��W�.��WɆ�C�	�ϕ #��w�D���(�Mc�����`M�C-��#�n���o9J�rSL�!�J|d�n��v�Ck§nc������{�M�*v^!6T���U5��.,� �|+�?���Լ�D=��n��l���LPe�g�dD Y�a^�|-��0,��
p��8��"ԁ����-��9̸~Z��C�뚐�NM�ᩈ��;U��P�h�#���#���Ú����@ʲd.����
>���nY>-3J����������ljX�`�dO�2��V��\�����A+$��� =��S�X���H�{�� �>^{
x��_r���4Va=��gY,;X���0�I���~0Q��!$T�"��O��G0.��Q[���ښ���}��5��F_�"1P#7d�N�F������;G�uM5�D�DU��
v~Rm�8��Y0s/�MF;z!�b�6E��=�82��vM��B�2��[A$Bzr�9!���G���>� @�m�@�H� 4��r'3/[z�Q%c�HB�n���g�F�z%� m���ەz���V�:_O�ܻ%��3�f<�aK+�����!���>|��� &�C��Il��_�& �E`�u�@��!���/k�/�AB�:�3�g�Ii+���Ks+����B�ԏ��t�c|fS�\�1�$:l
ւf�:i4��2�E(:[wf@,��X�� 39�6�@�.�|��{���M��a�Ǥ�GV�D" �5�
�C?i���h�-��ʿ��fg�m��e�9�mW�Y�%?�E�P�Ơ ��+���%>��ne���huI�;b�;��U0��H����H��+p�|�?�����^�F�èy�d��X�1�}�	�!ү�z'���⨕������%�7�UPM�(D�,T�|�>�Y�Z��"����!+ĥY	�6Y(+E%u$ =lZu��	Ɯ2�`,��?!��j��ė����)��t��"��UE����n��G���
o��w@Vn53~	ݗ���~��-�T�릶q֮_Z�}�.�5�P�t��B��܍n�t�.u���q�P�΢��K�
�I��
�|.QM $��M�¼�7��X��%L����4�C��ό��զ�G��-z�tX�/��%=GTU/B=�':/��C��_�`벬zJ��U��Q/��1'�6�w�8�������K�d�P-�]�D��h��%#��۱,�-�)���Z�2RЄ$�&�M!���(������M�4:^����#ZO�\��H�K��a��xk2(�$l�3-E,��8����~��z���#��=wE^�����-&X�#=�l���(=f�ݧ�M
���5:6��G���rׯf�9.��*{�陣	;FV�av��\�0{U�J����p`�\N�?{�T۔-{�V��~��,�A]��i ���O-6~5��I��wݼ�N��_�.5�i�� ��K��w���}C�oJ�/^[ї�<�Vx_���r��M���}mh̻��QLD����U�%�?l��?���D�&�J�+сWo|���M�z����	�b[���
%�U�7�i�[���	1��ܽJ٦�i&ߒg	�;�l$z`�8ם:�b��p3��f�r�c��[H��F��J�ؘ-����Z~;�;�g��9ב����e*1��Mb�z#M� L�|�=h��S��֌Y�G�|?9&)|"�z��h`8�	 Me+6�|�Z),3�ޕ�W�H13��<�zQ�|�*��IXS�����j5M������,q)��Z�6���Jז+��Y.4c���v�\�n�%0�:�f�8����e�JY�GR'No+5�f�x��U�O����L)uq��Z�K���F���֘E��A�@���֞��>畕y#
q�B�4ޗ�٨�� &_n�E�}`)̃nZ
x�����j��X�=����3AU���&�S�E�WՏ�Y�dhf�\�xK���z�ǝ��h�#�ȥ8j�P1j���W����*�.|��E_mUBB�����]��`�KX7���s��S�=#�V2>!���!��ގJ됟):	)tv��h����+ȓ��u:p4�d��a��r���(x�T+i���4h�!��\0-� ��1��$N�����l%��^}��������,a��w��۞���̈�`��Aa�f^	��>��OpD�k��A#1�j��ū9O�. !3h�)A���e�y)b�joj���l����˵�;¢`k$��rm�~F٠�g�2����̅U�NO4�w���e�Q>�m����R�pu2�܄�މ�,ə�!��C� �������4&��d	[�s�Qy��M���YX�UB넼`b8� �5~�;����h�5�����9�_�� h#x�mu_&+�S���`;c5��J��M��` ~qD[�.k��iV���+}>��NM���z+l���/���A�3I�ϕ�V��� ��t]��H,W���8�ߜ�w��AP^�:d�&[;ʽ��z����"��a%_�(��3U�u�z����_=�<��D�����Ǯ��$���"�T"�+��_kEG�ʉ�}z��fzN��.4���KԌj��])����^�>N��G��A���͋�He��FC�(���^0�o��}�J��\J�#�S�g�!V$�mmm+���|QO�gj���`RZZ��g�KT�P{�!/��%�S	'��62�+0����r	h1K'C�-�^�&)
��I�+؎U������Ϩ(�^_⎆-�b�����o٥���+��/�0\�9މ��<Z1��V���{��q���A�fL�8f��<it���埣�&0�*`E��1�����K�h�]e���'IGiU!}�h##8��t�\ߕ�P�������np���ξb�(���MfV0_ݙ��)`u�:{(�x���hp���;��b���:ͽ������F�-�[~$�;��򖀋{��Pc`�@����߮�&���`�/D�'��r|S��%t� @��)�w��|�T�}�����שq��y���X��p�N�X�@����D�8&��NmE�])��4��N�<�S)��l;�<��f��	 >ቬnϭ�?-�g�-^�&�%������.VyÊ�Q�F�d�Mǔ��~��)��}
46h����=���K����ÏH��"BO��o>	��7H�� ڱ�K�׺�O�g�B����Z�N� ���nq�1g��慎*)���;��O������̤��+	O�� �X1;?��R�[D�U7���C�r{�&%��2{�mԮ�ءÛ���R��a�Eyz������ZA-D�BE[HS��6x���̭��^� >�O�� �E��(T��h�^��(�Z!c�×q��Csxr���L�:��V���'Yr�R'��iGp��ЫFj��0�ɧ���#l��>:�~`v���1�B6����V��` C�O����������N���^?V&��ٺ���Lxd�G������ q����49��˯�������G�Q=�2ރƮ�j/s�B�a�%z�<Y��z�/�U#�؈?ei�� �d��m0W�~��a��%5�\w��$��e���$�jݲ9��>[��.���*�Y��M�=�*Dǃ�ծĈ�����E(���VW�!�O�E^�f�M�t����Y[:4�ܮ�aY��	1fh9�5�eL�{8ˍ�&0���
�Yi�� ���������ȝ7�_����SH�!@2����Rh��2���]�6�ʯ����-w��Mė��V�e@T�6C�h�$ط&F�wM�&���������ш�9 {�s���N�!�V���\��ݿ��!�_`���y��,x��w����A��}��bά އ�O=4.ի��.h=���n�!������X��Z|�˩��\��� g�Y~>��4�t�ȼ�!΃aJ����JRӣ1�f����zGZq��Uk��&���[ ���J�៮Hv%ƛ�xř�XОK:��n�UcCp�ܦͨ���M��Q�rt�W)���U,��Y-ڬ�x;B`�!��׉�c���I����-�ñQ�	
c��:�K��A��Vb�����u���mH؝/��_��ʵcIp����2����4����hxQp�e�J_���t�.�~��)zP�>����̡�����z�Y���-DH�M-�&����� �x����&�/6]��9M:Kk���i8C*bqy��sB���=.���8��Q�wN���+�3W9��{B�:/�aR~A�l�w�*lB�ƃ�^[��"oQ}ȏ�e ��m����k旛6���,�P#"�RK�-t\3Y7�ٓ+7�˨���A'��#��� �{�5��f�'�i:/��g��',I�� ���*�}�p�m���-�x:�d�Y�4��B|o����,��V�)�K��m�)��7W�~�dDb�h�G ��	E�ἂ������	#*�2tO�+,��R$Yh=c���d�V�c谭��=x�G��2x��?�岆eثb���/�U�}
w��M*�b�����db�}(-�V�]lc,=�,�m����)W��/d�W�G�C<��9r�S�v������V�	�8�z���?�z�ؼ��r�E,���J�"X����Ͱ���Q)a-�Ϣ=���&� (ʞi��2�M��H�׌E�!��a�X�!E16G��&uR�L��Ǒ˙�C��SQ�w���yRC8iHn�����3��0r)��0Yw�D�A�8��s3�)[p�����q�`vLsJ�dP���7�$�L:��L�q�3��x(זj��+��g��p��U��eE�TW�趻��O����SMTwp�A7�t?'D`p��`@��nEG���y	i5E7t��/�Ԋ�A�\�>��J�_R�:X���_�d��4+?M 4�k��O�VM,�d���84cg��Y�_�t����j�3?)g	I��`�_L��L��|�|�w� _	MwĘ��~�-F�QEXkB�G?f���U��(��sg毰��h���R�=��2�FR�M���.��W!)�1hQ"d.�'\ ��L�u�Wfp��nkT�q5�~p���:���-¿�cg�5H۫�Hp���s����є��Uv�����z�N,W���{D���arB�a˜
���N��ڶ'K5�8�/�5�������P� A�����cpͭ,�ԁ`�Jj�r�#{��6&��V��I�����M����<D(}����P���	(ˎ�K�f]8�1�@˟���K�.���н@!^Ǥ
��t�(7<�Z��a�:&�*��P7ҹ.�������v�������(	O��w�ЋM��ꢰ1}�!.��?�}OI�;1
���J6H�)��R��0���vg�U���6����V�Q[d�'\���T27��Gj�F�L�Q����7䰛(��(�.�KzR�BN�s��ks����qm�P��][z�I��f]����d'�~�w�tP�%�`=*�y�d�P��jY@�I���E��8�	Lɸ9�����a��!�>��fl~���bi�SCB�6�А��O�7�N\-�nw��8M���/��xȿG ����L�S-��k+��%��
N�ta�@ƔF��)���q�[O��O���iG<A~��Y|-(�TCG�+_i֊�8z�R�Ht�
kR��F�)b�AP�/��s��)�狞�N�'aϭ�"�ܘ��7�٨7�-�Q�>*>$��m�*|�Q*#�W|�M�'�|5:�RD�ٵH�Xu��nɠ���myL���3��'>k/���K��g���c�gkH>Z���i�ט�2t�J�lp��Đ!�m�vC��cm��m��;&Q����*@����:Z"�fJ�H���kn��{v6��T�X�OnV�I��	�����U�އ&�;��М��`z��7
y��[��i��)�F���ի��	�^kv��Z��"�3��ES�
MƃXI�mOq�*S]��<��DM�m[ª8|'����1&����Hk�����>]�S�ګ�{��b�RE���<4�8�=�(���􅜏��ؓZ�Bnb�Uv��ZbNu;AwB�"�z�d���U蹫��3씍Se!�y*�+�U������]�e-�g��E�Β|�P$�.�
���-c,�@�V�e������!�fWE�j�=���¼b��Nt����G)�n���/m.���N;��֙ �)��(M������P=��,0-�\e4������jV�����`�t�RR���M�4�D���^�Њ��&���;L�]���{[��ά��O�N'��,�;�!�h�"J�u���ǁ��Z﹄9Vӏ]:fe<i���+���i�,�^��X4�v-����i�Lc�Lŏ��G�tp��5����f����Ϊ�bq�o��,x�NT$D�eV�1�����:�`��Fi����B�@���ZZ�VZtB5���y��N-�S��\�g Ӻ6e�t��:�����B>~��♳��MxUÛ`�,�i�x ����O��X+�@�
i��@��]�V��x����`��e�Lb��&���$����7:�o�Eh"��f���q	��3o-�5������`m�+��1D���d[&���@jk�Y���D�1�`��,�w� w�d����V&��q��T�_�vT�ꏳh�AB��'=`(�/l#�4I'��5��U�"	0�ֈ��Y4 �����4���	�T(@F��J����-À�6�U���	��|�4C�}��SΡ̳|���ؘ��|������h�ev�B�N^,Q�J$�vy��HX�~vo	�^j���.3����L�Jx=?=iJ����8rj#�����O<�Acms�SމU�s�����p�^C�M�c 9���w2�\+0w�3De~�1�����8�d�~#��i�b	u��_'&��Ģ�zv��c��h[E_!�+B:�Ce���Bi�V��z���)���L~�%=����b�3��w�a�Y�w��f1� ��2"(t"$G���Fz�3�E='�^�Rһcn�g��!���8 ��nX�0�2/f�9�{�>'S�*�7�����TʼW���Ijo*GjaEʧ��q��:��VQ��������Mb����Kp���,��<:)0jc#�Ya��1FV�Q0�\{���u�EQU��n[.�W�_��+���c��٘��"8ƔN(��eD�^a$��KR[Hs`��}���v��R�k��'��}�'�9t\s o\��+!f��w�f!��A��*�}R��V�S�܀�L�?��6���5α<S�6;Np>�T�r�R$5k��4,�kvk'�Pc�����Z�����&{ �q�Wv)�P'��4V����ҸQ�;�y�sQN1�S)��b���i_L�!�S����)�w5>6<2�=�W	��a�1_����0�+p��f~d� $i|�f����a~�g�)�g��Q"^TM�=��<�*r���
���*����Q�
��6�?-λIJwf�\��W1F�[����e�����:IEC�-t�y#j�����=�H������9��H��.oY�_5��Tr�W�{�;���&@4U�/��	>��ad� E�5˛�}��J`�%���D��W��xϽ�A�T�@�mk��MT?�Vo<(�m NQ;���D~6����V�;As�tGL<C�����=��K�W ������X��t&�Y���=�K�te��ݞ&4� ���B��N�l��ʁG�%TH�/��f	�@�F9�0���q���6� ���B"�	�%�t��Q��i�\|Ŭ��M�v���)>�l�W�#�M΁���5$�[=|�w30m� ��S@iM��։���� ������-��F�.��bK����r�J̾���b� ����h#��`��UY��ݥ,84��s�Ej�V�ͭL��~;\q���ls��Q����, 	�x���	�or� @�Mqx5 �h�&h_4,Wj�"S{f�Hs �W��
�*\����E�_�@gC��~�*(��QpϾi�-��2wv/SEǿށ�I�M���fVG]�7��i��8_����}T9����Ͼ�֥7jD	2��>�����c쇘nҐa�rm$����,�G�S�&j�L��Y]/ =�G�SF��GNiɮ���FT;����S��~#t�z{�|�2�5	�C�2N����b�d-������{���e@�D�4�Z�0�6G�gηKu��{�~Ŝ�����h��5"��{��q�����3��6N��v.��_	aN���j����,X(���pF�8��)��1W�GC��˔��+�aL��=˕v=i��! �|�`�Q�ʧ);qP��&��#0�)tPs�t���=�m*B�*�����m��5WE�~U����Z�)mgƴ�Q��<o��"���t
��ֻ^�ڛIi?b���'�0�b+�]
FO��e��L�n"`3Fϫ�	�����Q*B4E���?�m ]��-��S�چ.����;���~豙S0��^�ť�:i����R��s��.d@<�e;�u�Y�C��DV�~�}A�#
I1�Vh��lT��k�n'y�	 ��F����d5��IK[������Ӯ��&�\ҘΨ��`P�ٍ��
BTI+`T�����V�Cف0/�r�\��0���)����zV\���K���=���������;���)o$�j���2"��jTd_��E}��� ��.7{y,�u]��gůP�>���7�VM��j婃}5����1i��l��Y�:|���s-[�������je�0p�G�QF=Rڷ�k�_(��