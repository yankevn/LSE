��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���H��?7܅�9!T���.N��i��(<@����+-O�Jf	��al�LQ����'��X�K��(�])����]Ƈ��r�r���z�n-T~�5bY��ӣ�ZÍr肸�~�|h)*��d�̊�j�,Wq�A�c�%J��Z��7ο�����y=�	�@✹R1<�]�H�+�]��y�qi�r-�;���Aԇ7S�� �pe���Ĝr;�[*�Z�@jIKUi�����x�[2<�S?]�H&���iZG/�/C@��q��	k��&e�]bY�L�kþ�o\y`ᝁ1D�!�1|2����j��^���DAv�2Z_�=���
���?H>|z��n8����r_�6���Un�*�XY���
��/��a�z]2��a�X�؉%�������'b�F��f)���Iח��W�L��*	�T�S3�}�[�Z�Џ�r�Q�Ф�./'�#��Q��n#�
���"���rv�EԄTrS�2-�(Y^G�����wҩG�E�	��Ȓ8�ft�. ��t	'p����"b�X{��x���æ��������R��C6\�X5��8�;V����5���(�7}�Ƃ���%�"= c��Q搳�o��t�"�&e�r�N%8���J1��_�b�@Eb4�h�|�S�I��9i��F9 �<��0�Xڻqw��$�Q~n����n��K���	5��%�T�.c0V��O�Up��?d����^L#�4�6is8�N��&����h�S��"RS�\�I�hu�����j����fX���:e�������k���Q�ez{M���l�/���炳�r{�,c�
�N��X<OcSY�������(vH�"\�jxu�l͸�ھ4�ԭ����t{a��M�oyꩌ��w}��P�s��Y�>W@|�T�H�0�T-�/<N��g���3cu������zfX��}��όQ������뀼�1yq.wbuNG���I�itf�G=��Pq�[4}W>Qȁ��x�_P��c�%^��::��D<X�t�{��x��2$'4�shm��àL��3�\ŞY{T|�m�Rҋ~���7n+�I5c	6�˻�M�X��֚P��g�V~*����M|�I.�$G�k26������+8R.^�e�ۆ�4�8���,5�X��a�[�P�7�.�L�X{���.��;�~
��9�4������a��㾮��f]܋��q<�wm��R���)�@��Zi���=�OW��-�%�7ܙ6�V����ʌޛ�n\9��je���J�lU Rb󬹏 j��U豗T}�|�LX���]ueXj�7����1��e)��>��w�8�B�)���Ǿs�0?������n�Ԯx�	�x�x����
[�D��.b��e���u&s�4���n�C���T��å�͢��w2EcGs�Ɓ^��koK7Z��k�z��hT��V:�*�Xd�˂�,.w���Ѵ�l����X*'�cK)���߾vͣ�(踐��8�?���Un���G����-��\�+��#s�,s�~��&��S�7�4S3�c[D��[ �+qv��أ=f�;�4�-�D�0��!�H�� '#靡�	ir��3��?�|� �����e�x��`��u|�rzi�펒����P@s�c<������;j�3y'`)>�V�J�ם�'���Z���N�っ'��7��O�
��E��zIUhB=jN�% �a��D�ܼ��3)fo���"�k�ISO��b񂗇4	��_���+��L���#�
j����[�b���7dΔ2UR���nH�τL� k���6_EO��M=YS�6�]9�!�`���|.3_[i.�
~+RL�Y-g�T��e��W
�3��[w����t�G�,�u�.�#�j� y��/ˏ�i�P��M�N��/'�� ����F9���X��'���@��P!��������m��&�{��m��;��"ƪä�����>:9�a�Ui�}�غ�Ƞc���*�$��_����Ԃ��0}㱠� �/@�AhmE�WgE�%%�!4�deɟ�ō�N����~�-�Ni��Ѣ��^�����b@9 �ݫ!�Ыl�t�X�i�7��L$ɛ����:�L�Mf��"UTo#U2Q����Ua�����[pg�$��$�.����+�%]!�̗���{��1��O�A���;����v��.��.O�r�î#s%����:��vj�q���lqS,�r��T��[S�̵#�v�ϐV�)_�S����ܓ0IS�:dmOx/�	��~ϛ�=�e��J�[�<���.��؛�<M"l�O�� Z�#���dK��ե~"La�~"|BA.I���@��-7�c���,KX�4��/�O����W<�{a�h>���>�)�W�ctWIv����.,\��w;�{��R��*��0gNB<�^]�ݏ�?tz�^m������E�Mcd���[�!�.ģ?У��\���4��i�+��9��"=�&�.T+�� �ˀ69�!&��⩊Z{W�#���O��}7ٯOh��|@�J5T�p��FV���)�B;����r��P�$þ=�s��z\@�hKNn���?�"2�\�W3/�nR�h_�Է�U��Ýz�R<��@ő�����~1��j0|/["T������e�����cql�z� ��`�z�c�"��]3y�`�:߷��gX�m�񷷂��ԭi&��+L�swm��5CuZ���u�}��qZ�]�wZ�j`S���~X�KY2�C�d����T�.��g�|�haq�_g��"	��$cO3鷮�|�=߅�@P����=��(�� ?�Ty0 ����i���~
hɄ�V�ׯ�i,a�v`fU��T{,@SX��d����a"�Ba�7*�~mX��I�1�q�2r���I�E{q& c��.0\�l8F}O��b��۹%�ţ&�WF�&m'�����a��G|&R�������Rȸ�I���!��6�~��Lw �Y�}��<��l���v�H)�'*70)�wdD6��&Z�c��i��X:��%�i�^�5������s������JjCJ�M#rfG#���CcHn�����<Wa9� ��J�X���DX"4Q�t��1���я�Ö���%;x}	ԺdfIaI/�Ð} +�&1�*�J�v�%����e�#�=ЏiR�r��*�Z���ހY��ׂ;����_����(B��3���%�7~����.�2���H�MɦMͤ|�����kf D3��]��Gs }�%�d�'��*�v�M��FZ��InƇG���ɣ��r3����j_�V1"9SHБ�	�ZL�h<.����`˲�5��&8\[?N=ģ�����o_��)}Ѩ1M]���@�9(�\$ū�B���T��/(�� Z�vv��L^�lJ9�K)�� ��6⟼���Q�O���s�g��eՐ-�E:���+�E�mb/�k}�����b�c
����5�^��c�Z��8�'滎�����8��`Z#�"�}"��v8��Ǳ]�S�$��>�l%��L��v8j�/#��cx���~vZn�0YUUA�����ivL�p��52��c�'��nG�se��3��l
I�1b��95m<Qa�ĺ�01�E�M��6��v��$L;������@��I^��H��	���X��OqD�<.[~k�w���C��W��M�ף/\x���
�_[Q��L�?V�Υ̞���n|SҠ�-�[�Cl��=��|���U�dxHG�z�g���e�$J�\XXq��{�`_&.�p/���n�Č�#�$=�h�G͑��Ss��][��.��fy�nK�zM�>p�Հ�n?��l�������P�x�<�.�m}n��������w�Բ�&�$X�3��K�����ֲ.��qE�s��^!�ז���TN�!	y'��y�J+�uV��������p*s���#'��g�dv1�<'+�{v}�����Z��j�Lw�PR}�4��GB��A������U�����q�K�gg���3����<�����;�<����LpH�H+P��sf����_C��;��"̈́��K�W_�͜���0J��FxV�C|��@�L�� `�L����[?��&D��e�m��7��r�7?"�l�0�0�#�C��p�?/��x�t���D�!r�U�����Ʉ�ەh�r	tkb�E��&�j��1Z�=긠8�΀+�X�"�Z�!��&�F���G�#zU�Iv��F]H_/&�|T@[](��4g�b۠與��@���z�g�c2� {���XL��5�=zV�2��PL���NC��~���6�t4���*�����W�:i0���B�*�.u�� ��]O��,4w2$D4]fE��>�ܛ�h�b㝊q�^]��@���=�:L��`#q���=!�B!IL?�xpE��Pp��k�_5D��h�E�R��M[�/�ؔ�}������4��W XT��T�1<�	�j���Ńq@� :e��>��M������<-�V�𔉏�{7_P_5.��OO(e��$ ;
���_%E!�b��T%��"w�
��7�0�r{p�� i�X O�����*a9�0����3�S��F��Bts�0����q+8S�l� �g5�?�$D�Ȩ�jݑ�%d�ܨ�o��L_��'�BX���<Skߍ�F���}��5�m�"3����嫂�*i�y�JY�9	U���hi� "��5s�t1R��c�^�*_V�d:��OG�OP�("r��Q�yX̣?A���⁢�7��(y��|�_��K�f����?r�J��϶Ot�PP�d�z���yJ��������F}T�+�`��:*�N-:@� �ןE�U/��J#�8��Юw���T����}@
ϒ��g�r�ss� �����،tM	ݹ�$m�`7�� .9��1�	.	�4)X���^��i���g�7Ǻ�$��7J1S��}'�zPf��dS�.-��C�2 �¡�)�:�iv���H����_�=�s��p�F�Re$���X���8�Z��J���O�b�(� �4�0����
j�C��	��A�yߊ�/����|?_iݠª8�i�c8��ql��zV������*CW0>d:[�7R]��D�ƴ}��;���K�0RPk;���4���� n�ʈE���,؀���5��d�#<]~MV8UUy��������`�h,��W:������r�Y��̼w��sʮ,�����5�[�cnX��9LS��4��9�,>C�W���g.���-K�� ����ޣ�>�A�|���lQ�ſ�r_�_����F`�a?���b��
�������e� ��S!�� ���o�^ǰ��Lt�ރ�r�=�bM�0dX)�g\6n�O����+(�8���=9����Q�9+���eT��oZ�G��ߜk��p��k�Fz���z��p��i׋����hb���*M�"�z���N�����0��e�j=~3�Y����6�*�@�����=�c���9KUa�%���ܵj��\�m���� >�/kɺY�8��F�2-b��	�d� �$.$��^gYA�ݷH'N�.������e�;~ȺJ���1`�<>�� �dO����z����U�A@�y���^��V��!��
J����ovg?�1�0c�w���p��e�.�2m�ʙqv������2�)��Ţ8C�kԢX>��5I��&~uz� ����k=�q�B}����Ym���+ZjIō�2�:�󊠜e�V-�B��@��*ϓ�X����G���Z���X?ֻ�۴�9s��B�6�N3χht�`]���?�pd=�w���?�s��ި	Mo��k������P��e�ir�6j�˔�����P�N����i�eJ�Ktz�ݣ��N�E}ޟhuy}�<�w��$������%�� � +�ȳC���} "�ё-f.�k ><������$���H��P�\�y��*q�	��Ёi뽻���� [ �N�(ٔ��N���o,�7�}cD ~����$����WGC�d���ys���Z����8�Q� � 	�FR�����ߩA�G�iDѣ�~BՆAmW��:`�+(@U2����M߁�PںD�m��َ��PƗm=1�1vHNŏ�S{WH�^FÂ�A�:+�M�S@���D��A��7�;-^��:[N�9̢A#G��/R,���ꢀ�;rM[Qu�=֑|��Ƚ;b���q�������&Ӱi����v�����)��x�x�8(`C�o3�&L0>�� ��;@���s9�05<�9yj��V��w��XB�Z��ыkOaCɓ����B�UϤY�ջ|�EI�~�ݛ�ﺓ��ԊYϑ��'S~c_oqjW))��2��0"*�A9X��c�X�fO�X��$�t@z�%�����Ν�ޯ�h~�z��6�~�JN��x�lK uM|��Y���b�.��^�h+�]�~�
;dHjk�:G)!.�d��t�3�R�@Ͱ>�ߝ7!�1=&���xB�b�`��H{���H�����&V�&lS�{y���D���Mt'��TAI9N��N]�?H�W�&1P���U��;1u�����j���J:m�6�S̭��`��ĥ|n:lf�e�-׬�CY���Mñ2�,�z#�:l�er;���K� 3o�U�M��Y��c��9����Ȧ��ݐ��a<C��QE�u4�ź�9�Ȅ�������8�ա'^g���T7�m2���_"b%5��<b�%�>g��̵�z��u�E�v�J�2�`��^2�z3B2�	7�+�X1��g�!^9�ψ׻�څ���!w��8�����|r��Q(�'�4��@����q�E��]�9����E���h���̌��<j�d0��K�{	��i|�;kpRK�#!p��j����֟ij:���w0�S�Ñ���������@�v�oT��ii�LC���`]Ғ�$e���Z��	O����K'�� ���ʬE�����	Pĵ�/��G0{��^�����9�� �-ӱu�sm�E�1w���y^4���Bl�/7�WԚ��2tgL��oX>Uڏ����cF3�[�}�� X� �N k| tPk,߳���^S��hE>�=���N/Z] ��2�8?�����wHC�.�Z9W ���t��|2(&��X�q&=�O�������l~�f2���7�?� �T�QZۮ/t��"��L(��,]D��gi��7��R��u���OJ��}ڝi��)6�X5��.�5{�����OaM��g�����u�+L�/)�6�>G��=E����TC���t/��T���q��P�d���k��`�Q*�VIz�6"`:;f�Y<b!�5����x����[�d�6Kr;B�̢Ɔ�b �(k-��wv�#A;�4?�މ�9���n��Z��J N`�z��_����=�fk�j��r�����}��!�@�"<s
�[���^�7|�?C�n`>U���O�h���d�ZE�p͂�F���?�����B�����5	��=p�<��u�/��2�o@�7
m���2.��95o�����'�݄瑑E�z*~|�{L�?*�ƩԶ�><>��Y��&�grO�`M��9��S
����o+�f!i�»�'3��	�<()���y�q�,҆}$��FDň���C��=��~~��j(�󍕚��wla�Vj?�u~��w3-��g�e�U�F��S�'݄�|����<��S#g/�B�7��v:,����|+@J~�@�9�W��P:�Dh������re-T���`J���,�J�����]g1p:x�+�D��~�v�ufL�A�d�`�If>LӜ��:pJ�v4�� K={��L1���4�Ѕ�=*�֥��%$�oO� �'�;q*e�L��,i-Y��o��w��I�A���%.�J��Xj�{ch+�R�ld �m_O��5s�f#M��Ra�"-)eo�I�#��\tR�|�s���z�)�Q�����ʭ�0>�J$�y���k���r���;r�~Q) �'������Gi��0�I3=��`