��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��@�yU�ߢ�Aӿ3"��.}úRJ{%
�	Th��\��hF��� �c6 "�\V@�m<#ޣ�՞��BJ_,q���QFssU� ��4l��w�9�UC�urVo�_��\��>�DӸ�p���C6��� ��O:�>u�o�r����ls
�U����*K���5z���C�S;>�ŵ�#r�tSY��_��˙څ��,-D7����v��%`�];�[ ��wK]�����^A�o
P`f�L�/�XXY��E����6 ��g�����"��0�FN�sS,�y����b�P�eBOB�����|��	���)�4�������������MK�袿�4׬��V��2z�]kbN�5�Q�
��y�<��;T��rc� kD$wV�mD�q���4�B���Ͷ�ȃ>������b�1&���
s c���fL_�ɽd�v��w��6�؟�^Yƒd���Y��F�U�6]������%i�� K�s��ST��8��v���i�WE�
���R��A>�7���C��+J1X�"x8��_���*��xsz-��IC�%�<d���鶊���L�u1V����vf@E��Q���VN:+`��h��-D�㆏e����?��+Wc+��J@
��9�d�,�Jo��v��x\Mv�{y5���	�z'���#�ָ}�K_��/�Mb~��1s�f���2�}̋�!�J\�(�G`��o�xJ3ȅ	_w^�����|Q������bg��c�����v�;fp��z�3��E�o�=3������p&Z~0��X�pk�ľ�G*�)��%�4`6o���ɽJ�� 35����ݗ��ЙɝQ�������L�a��-���g1(���e�аwb��ش����>ےUɒ`����������*��D����N,�����vZ�?�.��J!��%��v������Oh.7o��mV��}�B[^�tx,]�9#��<���M�>���A麂�D��J�O�+~��,?n���߻�n����:+]"����b~��w��1�� �y �ߘϑ��I�WU���S��,<ka��]H�rˋ'�s4��sr;t�E��r�2Ԏ/�׷��S
?��6��Q|�]�uՁ@�h��G��8'��U�E+>���̻J}|���Ծ9�N�2=Wj��鴔|�M�8�3Yp�o.��r�)��\�z�F��)9z��~�jě{����Hd������m�ȥ����B���Gd�\��M�(
T�b獫n��X�L\�E���Z�S����o�&pW�ۉ����n?�1Q^,׽�� �w�S�$L(��}��s2xc�.�0V++ѸS �
��������`�8l2F䭆s���@&�=O���w�Ό���̛+���-i`��H��ڵ+ Zlw�qo�Qs�yq˅�+B����
-��iD8�Q\z~k�m{��-��uͰT��6)���Q"g�-9C��a=�Sb���L��*xe�:ΛAy�r���_���T�O�'V�E'�0g�&�m#*l��d!	�M��_����o�����:��6��yeh�vq����1�D��������z!Ke��$�ͤ�z�L�1� ��%�c)n��o�_q.@�=�O�tg���,�FeC����� �֪N��9,vp鏍��Z�-Lb�K�5���Z����5�i�v�);+&�Tq�56��h���,��^�c�o�4)��=��n����=�clY5�jO��&$�g����;�\^TT��Lap@��$cɵ?J{iT�7(�.Ei/��Cz�lvT�y�����8����g��|
+B,�=	�	�����w�j�Y)��᜞��e��3J ���zi?�?4��2YD��`��� ��L�!a)e�+9��l��W����4;\n�1�bc!.��&��{b;�w㶙�yc�S���A�~���y���,�)��ے���3f��tl���p`�Vf����EXO����j>Ev��� ��Ae0�ؗ���X��<�+��e;}u���V�|� ���t"a0�e��$�Ѱ�U^���U���m�K��NJ}���c���M{��W�K�=�3p��nV��s1)m���N��*�4B�_e-0����d��c��"6���v,8�@���J.K�3���>/�}�M_!�0B}�3
٤���O�����"i��@�=�5}@;�Qo�q���� ��cW�< ��)2�$�d?���;��	����V&�s�ª*6���j�n���B���x�U�}��MA���<0.�^YAv�]87�U�?gZ��m�a�6U\X.����a�@ʇ8�k��Xsf{�A�#�UF�r����P�yچl���K�)���nM�Dn
6?F�#��޷�9��t-g��zI��^=":hz��ټ�Tt���e�l�����C�?��9��"��킍��?��QO�|{�(ɑJ��4q���]��E&e��(kv��z(Uͷ�2�N��B�����q	�p��|�=D��b����CS}��֕O��3�JQ���"�"�B�b�<Q*���l���
n���	�i�)�L���!�dt@��2p����̽�/j26�s�Md�Q�ɦ�D�C�d�}�3������ fv|�bme�E��K�;���װ�Y�mBJ�ڡ�B��-�7����Xhp��R��:]���a��$B��P8�K݅����z�}醈�u���ď��C^+�L�8�Q;���A�F&��M����'��&W�"�m��R$Y�c���z�l�.Ѱ� E���G�%���qVD���G�z�D��Rؚ��/��G�3��:Cs�NRBJ0��k�=��;�%;�V�o&�����H�>Ia��}g��e&м�4E*��̆��*�P�sw��!���~�]���g�"��,�@�_�^r��)��q��qdh6��������E�%�h��X��I�2^�C@#�CH悌�,���!���P8���+�,��=(�A5��7�u�"�I���+����5��J���o��٤�ŷX:�v����i3EP�*��8���tV#_P8Q]�=�sz[�u��VkXY��)|Z��j��j�8�ύ��6!f~N��H����ڤ� ���<�R�&��ƹ�v�wKЕ��ͱ8��hu�=��^��Q���KY��rq=2h��<k�'��Ҳ���/�J��x�t:�E�|;d��C��p.�޵|��Q̐17����	8�_�^�ZR������%ڝ�z��N6H�ͦ��q%��>H��>{�F� ���@#��'�wX���w����iٌ���J�U���1�f����q�����8�={U�>p�,�U�6&)[�{jrd��6w��;=C�T[1�t�.,����앚����K��i����$�.Z�Zڞ{�{�e���3��ӭe��9f��LN��!ԙxn�9�u[��@2v8���`�v��8�DY�g��S�`2T/���B����16֟_8�A� ���$���l���E�tF��i�M}�b��������keSmbz/n���׾0o�#`k��-��'R���M��k�g��V�Qd�	[�U��!Sm�M�=d�>�+�}��DM*��!�2�-�<�pI"+�z�(��}4R�^��~����X�(�b���T'^ #��ַ*1�n+�/U�2L���%�=b+�G�8�) �����Ӡ��!�zs[�I8��:��wV|�:��a~�����zp:	���J3C}� ����
L\=�Cq)�F�EO�U10J�t�։w!�q��8����\floDW�̠���՚O�ct��7���Sj5� 1s/)�%�`&-�Lm��%6�v�?&����+��Z:�Kҽ���`�8F�!�K�駾>as��W�qք5Jc�0b�,�������砿�0z9*�'0K�H���.�Z��n�v�v�[�{tgy 7&�MJ�|��8}M,�I�b	�v��Q?�B�9N;�D���H�G�NC�����~]�$X��L>���Yxe�y��:ֶ�|ݠݫ�M^Ix���,�qT�����`ߊ.�y��Ec�e�@s@2����x��2�\-�o7�c����0x>?O�H�m���M�}5p���O�������c��l�^\��n''�Q+�V<2�%��O�eb��¨�3�5�E�7_1a�T��Z%�!�m<�>+>&��؎��?���� ����JXb1k(c�X�6�v%2�G�kOsiȝ�_v6�h�ٛ�=�,�?�����`'$��h5����P�v@���я�1Q�:���ը����nu�U�V���L�)�a����v#B7e��	�T�'��+��3���{Ҩk�pdއ��_���Wm�H9���W�C��zo9eHM��M�L%MR��d��pg�L�xX��wYO�#c��q B?�l���s�E��(xq��7}n�N�A��\O�V�n1�H_�(�x��N��̓�H2�-�.����[���^�N�������dA�Ѵ\�G��y�aQɲ�9�7ƌ�U��6�������}(�D������5xN���֊�=L�+�:��Ǒ���ա�s�w��ɝ�VY��15�5��\�*@c�-�gTX���%&��b>ZZp�z���1����!Jjv��!)���ʈ�a|�M9n<_+D�K��I�����t��]:"��sM�����{nڭzрrt���cӘ�(m�RA��tb8`b��B�@]��A*
�q]ۄ?|a�ʤ�w��0����{a#�a�aK�w	L �0�c�"���r-V{"���G��Z����QD�g��PE���z7}����!q|�N7�/O��N��X�R��:Vm�u��ړ��-�䫝����щ�i�*��	��d�����C�qR��9ro�8�}�2�_xD�9W/�n9qb��\o��Pc�A�q/ȣ~��u	N� ��L[Д�@P?��#�:<�@-�D�5�8IgOO������EĚ~��[���N���5��ZkJ� Q+�&7I�B��.���YyJx�1���ra��;�7*�%fG�P՛1Z��bN��� �ן�&�+�V�0����0]��y����h�V�5mC�QS�`<�I	��)�yG�;l�'��t�)�p2�<a�~�D�9���!0h$�9�Y����j˾� 0���w"���M	��
���!�Ÿ��3�K�0�C`���p���%��넯���"cݞ���FG���n�Hh�Zn9��)��"jhC�vtF�|��t�=��-����I�D��&�W5 ���0&���݋�f�	���i���Y����ZWN9�;��d�ҿ�Rp<��_����A�>��^�C)�<w��:��n2|���K��+���jŀ������#���}:�FӤ�ZJ��#�P+;�p����Yc��m�mShs^��jz@���-������pB1`��-��c����"���M��ŝQ��2���-)���S�l������ԤT�A?�n�K�o�QtYy���y�C�6�p���V�r���IP�F.�ț�K�,DS����-L�5`�Qͧ/�!�zx0�y���T_Go�¨$�|!��8���;�sH�����X��u�z�%i� �h��s�#3�'�7U1dؕ@�9�-d8��!N=�'w�s�-g),ԇP)������r�א_:FwI���n�:��V��h5�]Dr�ӭ�Od{�p�����|iH1R닱���[�z�2ճ�@�ɐ�����z�r��(�X�4*лz���|��k��g�c�jf2���}�Rw���\�~=��?�7H�$���|��z�VAQ21�VIpMj{D�M����/x��dnO�����zy� �e0�cCϒG��j�ɸ��8��\R�SI��)������!�q*����V�G:e\;"k"�C�)g UDEۖ(7����v�t�Q�L�����ğ�;�0�8��5�6]��Bجc����7/O����#+2�<@Xq����+h��p����~6�<m�=O��2A���6�����o�����-�4���=Z�k�\o�2�ǘ�$�{*��3������{�P��P�w�}g�
�ؼ�x�+w���Э#�9���#�(:�B~]n_�T��N�Z����pm�T��|��T��q�)�9�p|H���S#��l��Z>;��F(��u�r$��&gE�,ff�Rr��ޥY�nx:Zj�H#��m��Qc�_��J�����ys��� 465Oҽ���Im���P�/��}��2{��ӧQSG\9�%��c\�2.�gT2$�_}I�u�A%<�Ya��'��:fJ~q� �>�Js�_&�|��@<���!vjU�A�S�W�M&����h@ ��W��0��]����G[M!�Y��W��+N��d�I�!���m�N4���Tѕ����c0*��|�>6]+!���o � ���s�2<��n	��8L�����7�ҥ��g.W��Z�qM��0�B]H���{��j!S��+ט.`�B��"�vn�Cȫ��+�*��,������8[��3f ����=p>�q�s�|8+�k�_!���ٔ�A�r�ȑN�y��K��Z�3¾�����(���@Rb�l��u(*�U���~L���AX�n���Xn�����i�0����%�fl5r]P
Nb�I��!��1��`v��4_ߨ17������4@��_5%Q9��'�X��S�p���K��O*Z�uD�jt�I�`
�6烛2o+�V�7ˬ���=�)S�-��inǪ�]�܁ ��zz�p�+�1��5��@�(�O���Y�xN/�PO�6$x�5^ė�] �˻�!+Ubf"�˽)-Zw�0x������j{�n����~Y������Y���y��{2m
�A�|*�[U���mu7,���k� 2��Y3X{"*�#�ě��T4\O��7�-u%7u`Q_&q*�pN�aba`%��dP�Y��GN*���;Zf���'�SU���AU��Y�+z�%��p��`�6W"S�udT|�C��TK��ߔLF��R�'E�����
3q�����:���%�vJ�z�Q�3�폣[ ����Wִ��?�㉱�������o��':����{K9�Ok;��0��բ��m0/&
G�����Б�G��W��y8�����[#r���<?_Mg�fؤ:mr:�f6�=i[�̷����ɧ:�],r�׻	kѕ^�h�0=�J�xr<�z�̋�ju�������>3T�Vh����$�eI_�� ���N�ލ���m�e�t,�^�3�Gg%-Q��J�8;j��p�7��t��������RKiM�%��Z����c�P)t�E	y�&N�[���ʲ6�i��������A|�����RCc�����t����'�]�l@6"�ZtR ��D��N��Y�@�>��-��L	����-Yg[�wZ(kE�}��/�N���do^]����(ܬ��D��GD��S�W��ȼ╞�#��H��Mj�{�P+�@�W8]�]돽8#D��"�H��Y-����cE�_*�ݩ��J)�@��:�v$c�V̞���t/K�d�eJi� ��e���|z�=DAs*�.��.f
ŦUc39�*�?�P�r�=��n��%����˜�!��.Q��}����om��~�J>�S�}�uJ!���a
�14L��H����fQP�b�7+�qȂ�6�@�	��Eps/>����́ %0e���|z*�А��{��
@q��M���c}�������zN�s>f�ٻ��0�s&7,YVIG�G�^[H9�L'��띰;`Z�Jl(r�T~��e��
�*�+�G��m�䂾X;�.=���;ն�6K�@�QЂҖ��~����&K�:����j	�b�7�h+�1{�S�ډqn����ۆOSΆ��arQ�!�wK����-�����B���m��!�O���rX��v��$��m.m�>q��L�eR��9>"\�jjm����7(�_0�H�R��F��&��@O��0�sT�Z�n]�i��[���,,+�֔��>�%ݎJ�o�6�g�=�����fFb,�+�_�Gg���<�Єm���F@����RŰ)4��:��S�.��M�rlN!_B��ZF�ܗ�����
��e
���(�/���獂�V"G��c�&�xj(�t��u���U#��m�fP{t#�W���ң'�����pB�L���f���V������i�����s;�gc��A�M0c��,q�Z�ި2��m{A�_Ҕ�3D���b���o�j��ǣ� Ɩ�G3�z�C�"��OX��� H�Z{�)0J4D,0=�&21�i_�Tj#�\��#i��m4�f�#cm@����qTaK�]��N�j*Tn��/���
]EdO��@3H��5�a$�������<Xօ\Ʌn�(��GD5.���F<8-f���՟�k��dD��q=���I�w������'��GD�,.
�i[�Sv	�0�s����	��Y����OՓ��M.�_j<ɀ�|AZ>>�;��^@҇��
�q�������;�V]ҷ�*y��1J;��$���J~���F�����<������j�nп����ͺ��Ko��mG��*���St�$�5|h�`x�%蠦`ǆ�e��]�)��҇,]�F��m�T���j*ٓ�<8��#�(�mZ�]�JF7�������nk󴷕�b��7� ��:t-_�v�eK�����f���~qؘs��!����S����n��/�b�
Ex�Ju�H[�	�af�!�	~d�}1�m�j��ᥚ{������4'��И]c[g�1nC��h�2�q�/�}�ⶆ�C{)N쓜�ߜ\�`�!��#��>IT�@�+��`�VH
_�%��<���/ujb���J2�S`W�W�N
���Ly ���OA��9aZ��%�3��g\�`�j����d(F�hh/��t
�