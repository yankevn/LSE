��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K����;�U�����wh���Ո/G:b;�x�]B� �Uص�u°T�&m����Inx�F��|�uR{u4��GH�xh4��9�%�\x�c_v�O�h���i�p�����
�h�����J�L
��lA�Z|�~����1�=����}�k	��XV�Ŝz�4�)�t����W<�$Bm��(��SBu�����W�E���M�-��j'��db��Zm5NG���2զݟ�u�7��~���f0?�J��=�K��\��`0�ȑ^�\��}�j+B��rh��S6�D�*��b���^T���r��)��zÐ�ᰂ&������٤���دq}����E��#@��0Z�f2��w]�Z"�][b�s��$K@���j�ŉ���舂���P�J]=�9Y�~򰛩C��}�yN�����ƹ?Mk��O���3_1�˰�ʯ�
Y"@�w��Y�@���k�n�Qxpx-p��a���w� �-՛10k��`�
��nu�amB�"�G�Ns�Qt_ ��s }�~N�m�y\|��-i�~���GGү��=^E�n�^�л<o������]�[�x'��h�Lҝjr��vB~5��;��7Ki�2(�����o��q�0
?�7%D�{��~\Z�W`o�7�P*(%:��7���U�]O��l����%�^��d����H���
��$ifȖ���bd�aa����&kBѷl�{)�崛:cF��4��Y�O����-���-�an#�3K��.��,ׄ�8�q�z��������?$��9]�����7���l�oL�����"o��=�j~��ap���J ��b�2r��0���Ç>���t�, 	O-��W{Ɖ�NdY�J��6�A9�PvwZb�n�Q��_+��tJّ5EJ�:��UP�B1$M�ǌ�����=X�i�Ǿ�䝹���N-_�_5�!�0�mxz�U��v�����
���ϕ��-0u���m|f�<�$D"��r�goHr�ak��՜է@�0[
��U���$!ϙʮ�]Lz�����Esز�K�h`I�{?���E'8��^��W^zG,���e��\��a��K>��Н0�?a�D��aҋ��Bj<UU�g��|ess�rd����mh1��rf;y	I7ލ�|�d�Ó['���w=H�"D�:q�^/ו�vI;�������.������,�<��J�M�\x��QT�è'��A#Q�p0KO�0>��|���L�%��K���s+�2�EZ�b�EhK���}��8�����Ј�a}i���wi.� �����4R࿣�&)��o���"� � ��M2ɬU9\��RA�ա���0�.��e8�Y��)P�(���ah-j�v� ���	C���/}�dOU���ҳr�%�f�U�v��f,�y�R�P{,w�t�+[k�T��<~�
�*]��v�i����
�]�Wj��w|�}�$T�����N�­��j��J���G���9�B
Ȓ=�X��y��DL6; �]���V�G�8�֊��wa ;�5�;q_U�vX0i�h��!�v߹�Z�l[}���s�~3Fb�T���l-����n"KK�$J�M�^0*���x;ݜo�g3%Q,���b�l��EM/88���V!.�vd:�ctDз�<�-���	�Y�ǣU ���B�,�Bs���	�z���^� Qod�1�>����IVB�(i�=	�z��͟r�5���s�P^,�XZ;9��|7vGq�A-�x��iΰ�[}��.vУ����s���8�m95����]~�O��iĕXW�0|��f�tI�sE�ޱj2��@���RY.�_�Q	rM��ʔ5l�6��9� ٷ��p<>��]{A���D�j��WhU�*�5{s�`�V|;��+=�i��ܷ��-qHɶ�a�C�;c�͝!��b���c �5�qXb�z�����zߤ���,LC�u:�|\���bsCDk>Ō%}m�Yf��-���A�"5z�}��y9����2��M2�ڈ��	m%rڒHbjH��W�RjV(��@�N�/�IL���`���m�6q���y������V�ʌP�R\��ʑ0J����FX/��͚��"����K#�t1�g��v�{r� #��f,lX���l���no�̺rT���9^bQi/�Ze���O�3'��4�p�$CM�rxc3�<V8�(��P�h/k�f`Λ��D�bJ�7�:c42g�kW��e@�=d	�X��S��!��}lƋX²l�p[������?�L8}�oE����V'������2!�a��X�V^.�!g����nz>Y�_���1�µ�L�]e'
X��u�A��@���g��s�1c��?0
�}����ߛ�=w���!��\ 6�#ME�!>�del�7�����k�w�1�l����T��Uz������L�� aB�D�W��twj�9 �d���R���}pxi�v�����5�E,�E�*O����_No�����;�_ðM	���������J�n����`�*���X*3?��0�Z^GB�sK���>\R�N�T��������ޞh�����vx#+N�ɬ�K~b��]��g�2��ڜ�)w�-�J͵"�H��q��Yg��:D�6ỳjq~��<׾��j���F\�k� OW xT6�8���`�����@�5R���YQ^�1z��9�}gA[ �T{���C2�/<�y�	�A�#sK����CW:�:��8@���^���"���/0ST�C4<`=1GTI;��D͓��W:\T��bwJ��%����f����e��n>�� X�4S�-�33 X��2j�뒃&M��.!��r�І��9��Ov�$c�Fpy���^�2 ��ݫ��ǆk|.�0��:�}�H��M������6�2&�����Bzr�{~�^GH� ��+P���� /�Kle6��kA��op͋��t�&�7hd����3�sO��Wr��f������� ��0�?�]�Y��3�eˍ���)�_d[�¸<)��0�@HZ�1պ��#��%��k]mf��A)Y�+��P�|o��WL�W籊Ii��( �*~M:��	�N�����$:�{���8��� �pML���U}
l��?3񴜚;�eNA��������^Q�t"��n����������O���+8�uU����^`|\C����b�����A��
]R�=|�Y��ݷ��Nʠ ����qT�ZK#	~
]��w=p��O �_��zd�O2^z����(K�
�g�	�=��V�y%�(���x���M`3�j�a"�z���B�]+��߆��o6�u�}w��E�]���_�4>X#=�L�UF��X'�3�