��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��(��ѣԿ���:+��rYV��;��6��!�iG�{#�Rݕ_����JkK�ݽ4\�(��.*�[{��+����3J��� ���J�S��pթ�`�]JX��X(EЊ"����sZ�Бx���
�Bo\Q�t�����vw�ջW����ccσ�*^���%l���N�rd�!����Z�q0G�nRu�4Q� ���������㜕�f{$u�6v���9,(�l�Sj�[V�����&�F��=��{+��T��ca�ZR  �9�%s��E�ME�4�����Տ�ϛ]�䛝'����;��MmFM)څ�+H%��1�r��ۼ�l����<�K���35�I���wp4:c�*�׻��C��
�i84J�:츈Hq�Z��B씩�'�JD��4�K{3�g���?P���C(������� K��8��##M���Y以��5�DU��j�o�K�ِ@[��{d��otТ�q>h�s��i�e�֡��4m�����-�Ҙ��9g�`e��-�^���x�w9;{���QU������2�Y���^#�I� ���G`7�Rx`�k���]ω�o\����}��(��ɰbUޖ$��y�i���XCJe_E}��ƅ��F���Mn�d�]�E6)�^��;���X�Ǒ͖O�?u��+�
�C^~Q3&B�tA����\�ݏ\�By�hL����i��4�x�K<%[!�&�L#vZ/�6��H])k�s`R8NRL��N[��i���/p��n��JF@������o��X��d��;��G��wi"��CbK�/75��(�pĆ�N}�W����u>���k��%�ٸ�Ui6��Wy�!w��g̸��d24s��,�^v7���:�W���m��k0�E����?�'��>��!��o�N6�(��k8����"��A���0�R�Fh�|V�hfG�\U�H+�iȤ�V��~��rQQ��~W.{k���GT�.��zi�h��9J&dAFH��r�P�b
��R��tX�m� &�s8�MP��uP���Vj�/��w���<�ٍ�D�5��M�*�o�>Y�� G)퇘��>�:>��"��ۿQH#Sj?LnlC��b�u��7[��ו<K�T8p[��
����*�!�lnv�:>Â>����3)s]��#��6E1}ŵ���?]^��q�R�s_ۆ��Id���5tE/굛ĸ�w�/����]�A!?j4cJ�����2��aF	�n��dE�4a�����`P����x	z�Q��T.�W3M����G�"��$V��F�քr����M[äth���u���)�n�ϋ��a��q)3���,514r{�\������D
�6�s�>����ٻ������{�T[|��V�/����H���m��Gβ�����N�ժBL�c >"�� >�@�8��Y�z��:`te=O�lFr=�W�첀���%c��8�:�OG9ԟ�!��)er�(��g���\��l/��m�V�L�n-O	�t�]`�U���
�w/�	�,�	F�U܇i��:_��*���WO3����6�~{z�l��}+ ��W!���Lv$kF�y^D!l�ҭ��E6���:<��,r@0�귆��d��Ûڸ�Mi�[�����t�<_�����}�^�n�/�T�b���br0A��a�p�׫�z~��""5�B�\�� jB�m݊�����k�?>k�����H��*9A�tl
^���{�u����U�]������t���^ B�٥�,�N���+«-)����3�WĎA���9�cU~ߎm
L/�B�(9	�m�W'O�����p�>���tԑ��(� 1?1�Uڨ�u?�G��Nͣ�i�K��{�+�s3��w�9t����ۺ�/�ߦN]&"��K�-���ճ �e������LRm(CKK�I�A�\"X{�{Wb�`e.���9�:����ES^S�$��IZ8��P(4���e�K�ʡ���i�
�uy9*k�ph#ڵ�d}yGK��Uxyy1�m����[8�k���雦�c���&v�s�Ῥ[��[�f`��3#A�է,ҽ0��*�Z��7��6��;�r������zK���ʂP7��W��+i'�=ц1�7y�̩�ՑsZ'�N$("{�ؘ|�������S���b��~������;O^A#-�71��iϋ2.9C��c�ioJmsd�����} ����U�������|�Hf�^af^�(����E����"�&�_�2�W�5��ِ�*P���d�Z3|�O�����`R�%�D�z�}.ئ�ӈ�o�����U�"AbH��� �_,�9�^��=BB�;�^�@�en��x{�$Q�_k��`��IF28(�c�4tU)�ڄМ�L�2��x�po�O]�|�B|�:�k�O'�RU�v�Ƃ�Jqq���{\%�E��0�,���dc��ܒ��Nq�I�Z>��&���q!�B��u��4�S��bX���lK�B�����
���`�ܣ=GJ$K,O�Prh`�w`iTwlwai��lB�<��<��[���u�K�Nd,�kBdrHvN)��jh�j�aN��`Y�ы�f�g�Eݛ	|�ng�ߕ�n�i�6���`�_�q�;f�F���T�T��i�w8l�+�4.�:�w�8�v���Ƥ)�6�@����^�h���Cdw��9�T�_�>�븿v��t^���,A�a��m�0?�+���Ӭ"�����c�}҃{�A=r�LM`�&;O���qr���e�xPj{On���Ϗk���)�����i�9�U�_D���u7�kVҦC�:�����ޝ��Pq�;PEŀ��'��W�)��(�ҽ�`ѝ)S ҟ>�|*�
N�$�|�uݱ�M"��0Ӵ����t����٪�:����A���>av��&��v&`������� ���Ì����M��E+�9Y�Y��޼ϪnA�������}���|�w�B־�- cL�a�*4�\� v��L?�式�72Q�;)+}Hߔ�[C��YG�<���I�ZmN��EF$	Lv!}7vt�Ȳb���[�;�EE�����H����lp�1ʤ+֫7]�z[}�C��l�<�aW2]@[�o�Yu���H8U��Xb��h��(��U}��(��H�p�������doW��hvw��!ߝ�r�;)�7��n�B� ���71[{p��֭��i	M��(܏M�Q�@C��Z}�B͸���_ѹ7��#H�6B��H��I@[CPPV��c�\���#q���&�[A�'3�ʫ�nW�ӓ'7ƥF����"N
��Ҧ]c X�<u P2�Y�i�?�K\���ư�.�!���N�_iE0vV���]Ɣ�_�V�OcPK�O�s�a�~jE����Q�΋my\y:��k�`���:�[Ҹ��8��ǔο"�$�)�q�h��!,r�s��������m���,s�P�宜.�)D�Ӱ���$�yVT���T_"u_~�z����=�-'.�=��SUJ_	j����E�zj��7>��q�M>li��e�p��o�� a���R��C�||*��5�.��6~x|�k.��t-���$Pzc�Y�_��ŀI4pF�+,G)k<�v[� m6�Ηq�\ǣ���B2�ܩ+��O���l��(̅��0� T�&�Tݛ����]� �s�yG�K裠��a.ǘ���G���5dZ���=���?�#�MR�b�K@�*(N<�i�b��TmN�VK7,UߙK��ڤ��a�0r���|���5�<td۸�c���GU��5��������\\��Xi?��`
~��D��
xj@8�:+�ű>�W�v�>!�k��3�{Nz�i��͋�xV� �I^��P:�]C����@�*n�.���e[s]��#�7"�UK�9Q�͝c䂱��5잎h�|���:;���kT29D"�A���~�q t���$+ځBY��z҃'� �j���S��
�	 �1��BN���e=h0�!j�����TY[~���w+(�	��M9�P�|�1I�C�@x�3S��nv!���N�Q��~���W��E���P,F�`��wA�Tމ�0�+"t`��q]�DSî	X�M	�5�8�r�)&�})Ԅ9h�l�N���)*�p�Td�����`O���mdR� �M�c�NX�Rq.���[D\R�Ip�!;W�먜�(~;쎍�Y7���;��W-8� ��59�6����H@�	���W�`�Խ�S��Mk�6yo�'�^�:�����:˜ ��\Y���|��be�M����KT�^A�eB�!�DW��K�����e�ҀX�a\\y����N������|��낝f�Q�ۂ�!����Q�Ǭ��v�����]�E�cD��r����C)�����N/�`Sf�H���6��1*Y��유ǭ@����M�V%��{1�[�LF��k���ǖ?M/�ލ�E�ܸ�ߠ2�G�x��
GO޳޻v��0�Ѹ.z�@�/��q�1�
Y|F{TL�L9k@���n�j���ɐ��l�A-� �c| 3������`/U��N��1��p�)�|��i����!h���|�{�jcl�f���~�a
�F���%�]��-[8Ε�tn�ؿ���=#�Ю�	���k�?S9�����B"��� %�����QHC�|r�����sC������g��{��"��w���r�S�Q��6��9v���9��V���m�7Zt�̋�Zpr�^pN�:]�b�+Q���Hsd���P��-���/�R)�d"ʈj��UY�uq*�4G��'c]3z�J8�D�>����<��s���jX?����a�Oks�U��Ϭ�2��E����m�1�f���4�<��\:\�|\�K
F�!�����t<�N�K�L��-.��1�L��;�0lUF}r�c'����%C%�?���6O�;��0���{~�ڥ
^�ز`�;�����²6��17}�Ų�ײ7S�r��I��:��o	;v��2O,�"lO��8�*o	�LB�+c �du���r����M��nL���}�]J�t�.�
T[��D��[���2���Ժ)ٓ�\�/X��ǻ��+!1�Dl�/&b��s��7�=#���`߹Կ�9���ް�Z��,Y���D|��.�7��=�� �:a78ɪxW 2(�2�a}�甅a4���C�%�`��������e��c��$�C��2+!�ܑ��2(Ʒ�C��O�d���7И��Ca;0]��o��׸l�O(�O���g,���L-��%�vš�o;��woa��]�k�a�!�����M�{����-������Y�xK
��HM ��E���qD2:ؗpR�
/���_�p�`���J�P�.鳢�#"9 ��7Q_T�Ew��q� N
�Kt ���b�4�0R��ͤ�����į�
��qc�g��ɂg3?�����?�̛��t.�?��3㫝�3F@�]x"�t�Ć�d-��/�<���
��ש�+�<� �:���q�3�����D?��=K��4D�	��+{���ԗX���"Q(�/�=-�d@<�g������7��� �1m��8@��Tv�f-�t������[dm=�-��#��Į��ফ|��#�O�כ���+OM��w/�(�:$�1]�3�q� b=�Q�����
wCس����g�W^U��MK����J�4����2�v��6�8���qd�_�9,E��������I�	j�"gE�HA��A*��OQ��J�����*�(�w�;��%��Q9݂��[���1
��@
�8�,=�$(v����~�@Va�eS=E�o\c��ء��J����S�	H)K����>d� l�><���5��Ig_o�wR�	���� 1m!̭�$!�"�IS�����N��2��4��;��������P"������i�����|����c]�g��曺��p5��Gm�C����
��R��b7�l�e 5V�xLl��oc�sG7����כj�|F���WQ����1e�@~��4 ��S��Ak����Bb��}�@�z�7������d�N?��v���*_V�J��ژ���dk~��/6�e�s�}VdK ���C�p��Tg���9ė�́��;}E�daُ������b"�R�� ����S��`x��+��7;C��o�y���qSr�M�uƜE���4k]��5���f���?�gnG�\�B���f�Z��Ì��wFґ���T�Fק���I�$����r{<�d�g� ۢ��{���/ �����g?�碁�� r���+�	��A_��2�?8mY���UM��%�|���!�S� �c�������*`�f	��B8��P�_Ќ�R��	�~/��8������+���C��"\�����z�/�r�c�A��B���x���쀪�� ��m�yŦ��F�@x抒����x�J��Ȁ�Q*B'i�g����|�
T3TQ ɓ M�b2WEy�0˗�?����8�t5�F��[
��K��1H1'-u��	�}���hƛ[g�Uq/�y֑S�&��w�B9R��ҟ�,��`��Z�d�d�/�Ik�L-�'��-�mk���'jDl�?Yr�>^&N;�́��=���I�y�}0�ϒ��Zw��Q�N::����� Rkz4�k�eޘػ�f�5��EX#:z	�E���d�`����G�� lDc18�b�f���`�2�ѭ2���y��.�MNg����Yص���ˆ����\'z�qq���eh�m��w-�"��^v���_2]�������ͥN �(���bʋ�c��K����S��יу��j�����\��zd����>R���D��;N��	]�S��T��%��Ї��%
��r�����m�7V��G�GE��|
t4�ߒ՘��ap�Iy�d,ɦ�(Ih���S����E�D�7[l~� ���^����K������5[y��>́ �E�=���R��,�H�+k, 4��А���+�� �Q��u�o�^(��qn���wNF7��Sg�Y�Ok*�k仿�X�+(o��Y9��`��<~p?�Y�6���7�]��;�BA�1i�~�����1���U/q��K"LC(כF5�7&�7c6� h�.Ĕ��T�<�ۦ����������PP4�&Ȳ�����L8�#����B�༏�'է�A:H���]	�*�%��6*���t�������+J>~�}2X�ݨ�=-�T�Na�0�9x��� x� ����	�#���PaqM��Ͽ�6b�~r{.��'w�%�D��儧�Ɖ�� �S�\�l4��f}����k>�ǟ�W�������
��K��6�|���"z���"`}r�O��2&*D�b[ȈɑV�/�t���x`�r�� ��ը���St.ir�Ng�.��"?Uuz�R���!��H-�Ɔ8\��I�?�!�gYM<��6�vc�a`��������Jp��ܛ��4��a�!MT%�p�r@E~�|��h��s"�����<X��hz��u�R
qI�����D/��O7�zJI��g�9��;����i����R[�%ݲz�}�i�F�j5�.��n������pVYGavX_�����a�-Ȫ�yےsH���R���Y�=W!{�R���2��V�ʂ����?��ɶ!�T�|�v���Q�2��8�G~`�N�������c`τo �Y���D�찂��#�t��u�c�B��>$���5��pw�i.A8��B�{��3�����9�l�����{�N�l�xK�w�a(C�T��%���x�	��퉙S���-�}�^!��^���T�����?���0�di�P0ER�pE8�\����,���н�⵪�@[�>�m|�pէ=S��0cV�ڢ�?�B�t�i���GU�f�!�G���˭	^��������f����ϰխw���ӥU`r�0��3�5��a�vp<.V���R�CS���`�!��BOKճx�g���7�hh�i^y�.v�".<X�<�ui
v]��Ň�_3{� .�/s��"������0,��r����m?��D�t��&�H� 1q���7�BI�z�pѡb\6L�-=����ڣ�����я�0?.�
T�H��[�S��8�"L�
1W)�ta89�6ct�4�I����JN\+����]��±��CHN�CTy!v���1�a�O�mN,�tV�2@��t�C��s�pc{8�]:����Z���z5�S�?E��Q�GK�0Zd=�7{ycǇt�~;�y�c�����p�x�d��`��V�N=T�ED�2�|2�Q�� �ԳbD�O$Zͻ١>���S~|�Lu���^]K��0�@��[��-�?��=�\��p�:�l�.�=������t N�����4�ǹz���}����������j�NL51�4��>�3s��9�YW�s�89p?-�y�T��Xv���L ��"�%H��#?(R�*~��7!��-@���A�8�n��]��M�+�:4����c��NxH,�}ra1��i�n�gP��{3�,����BV�+��5��e������$f�9�pk!%������_�W�fA�^d%RbG��Ĕ�:4DVPfW�ٜv2BԘ�X|�G��ַıM�i�U�������g(�'/��X^�qc�"��Rc�FvǕ����(�h�RXU�kÀ� ����Ѝ&N*?�&X�Xe�R����7zH?p��3OR��·�%n� _k��
G��1���2 ��9�Ш�'gԹī�^�Y4_�L����2
�ISD� V��O��X��[�wfkJA��t}=�����ea*
�2��g�d��h��x�O��!f����Xh�����1��pD��$d����̒���\A���SE�D�d��%iо �qPk&F'�ym�	"��i����},�Bd�Ҿ�қq}��P�3�櫻��'c~���kl\���^��\�H����cE�kY����U�����{d��
d��(��md!^db����UQ�zx���{/g$�����9�������`��,۹*UrCA.�׋aP�����
�"��yǙ���� A��쿩vۮ��w��$�uχH���k^P����5&,7 ���#pv�f��|��	��g�a��>���OHv�+L��]�����뒂�8���G;5��h�5l����Y� j( q�k ;0���Im�,�o���h���˦�yk��\���{�ǍO	�a8/38bnl�~��S��I���$=�~�_2(�Eb|B�yr?��l̉d�x�`�BB�y N��*��j�>�����ms��!��Cy�����p\�8R�#E�7�n�_5Ú��)����O�?;�o���T�52�j�ƅ��o�F ��"]��D���f��QX�.�F��R��������J	�:V�ř5PC+H�`ڴ�4	��O&ٌ�O�k3�0�}���%�d$���_�B��� ��m�-%�{u�=��7;8E�_�?����}�
��)/��,*�,�����VW`�Π�n�,���iw��Ǵ�����aޡ�2�Z�	�����u��]Z�@k0�'l�ҬCe�~��S���*�L�C��]� Z���r�����q��;�a.�#��~4�j�R��֎u�&�[�cls�d�2��%Ci����V:��Kf����e�T���QAƳʌ�a��29PM���B�-
��V�I��zy���T�f��?i���Nʘҁ�N!*BO�m�د��ƫ�s�I��?������;���*&�$�d���i-�4#����P��0MM��� 5 /���[ͮ8��*�2��@����*�~���
�A3�@$��k&����˄��s�C�ػ�7����Q�VN@ݶs�����&"��"3d�!j���K/g\h�����G��s����A[ ����9g�wyE����04�}���m����!QS"k���i�^/ū���y�i/6���w�MB����� Y�'uDst#N�\N����-�^/��ޙ�͛�{A�5F�K霌b��:u&�bդF��QY��W�9���b�`�[�6��4��G���sg�Z�����q��E�h�<���6��%���0��[�:�ʝ�����O���7�V)c�@z �^Mt���}�?�j�j-����5��~%���DGj/��b΀E��W�*MMtS�HvgGx�˂�������T�:���V}�φ�V�GR�nK�SJ��@�Ԥj����v�Ulm+B;[�?�3Ia�8/]��M��	�k���\�W{��4xc�"�������oz9���[<�-*�1��O��ŘoWu�5)0� x�O�����%OX_Ё^ga�*t�tj���6�Ӧh0C�D��L��W��æ�T%�X%��%�պڎt<����֥�A����Ma����\��x��i��N~��h󾢬���o��G:8ã�}�ߋ�Z�wu����$��@�8:��,�]pԷ=H����3Ѹ�`~�$^������Kt���U/��������X\|L�w�/"Q���-E^�BS ���z}	��
N.�0'ЊJWXsZ��2
�Ƹ��3���~��T^YQ�W���>{a�i�����o݇ݪ 0G�>b���HO�&!~I�Q��HJ�ISK���)���W�r����&�$� 2Q�*k�0�Bs�'�I�h�Q�hl�뗻=�q�?a��
��@}��.Z>��!�5+>��Z/�J�5$�5:vWH�C���()܍��#����ux��N@��g)�}���� ar�yP� ���F�W���^~��b�+.�z��c�����wk�Z��Zh<c5��q4��ʕ��bۋ9��eµ@дS9�'���(�wo8T�Z��p�&�ç���Y�ޑG�3�/�V��� s���3�Uߴ�a�S����iד��6��o|�0���lT�?�-��W���ա��-�=qh������]�k�錳�Έ>���"��fs�F�d �n�r.�*����YD.�9�
�J�&�Xt�Gʒ�!cE�iPT�$1A�����5m�*y;�N�Ekd]O��`��"e�,��Yr*�\'>�/|el/�1{��GK��w�;�KUh�@��jv6_�9����W�V}MM�D���I?�WhT/M�]|��UE�\�4\Ȩ7ֺ$lM��:\��Q�j�K*P���NE��4zH�+�X;}�R�(��f$��;�@�	l���n��z̝�G���H�sʈz@��*����"`���5r�#G&�\�
�	?Ŗɓ7q��n"�g_��62��EW7����'�&	���"���)�J��T2�Hs���LTR�j�A��M�N�G
Q>�������"K]�M�����P)`�T����_�[��M�J�M�'�ݺA�II�Go:���w*W��߆��>|�!�r�4�%i��Dq����D��/�Y�q� �rLd�:QZ�����氥k��4H�A�A_I�VK��*]/��zI�h�H�m(�gk�)�>��Ɨ0����P�n��W����-�N�_[P}Ժu��5�0I)_��(��6J����H�
(�aAnB�md�������HdwC���{�۠�w��F;��Z�}6��7>!=���=f���mF�7��D����p9����c��y ���������W�Ӌ�)҂�y���,r�l�T���n����;���]� �.`�e�".}��d��B�7�!��_�

K�(Kp-gI��5N��<��J{bG(��s�v�,E��������M�D�ӏ,�Pg̀�jkq�z9��+oQ%0`ыvT���1�؇��T퍩����G%�?sKU�εI; ��QDC��H�Z�V���.���*�
[*J������1P���m��7�NDa�D%$�.\+���F�qt��;���]�g��#]�[y A_~�8k�GR���
QB�c��Y��a���ȏ3�%잁7�ͨX�O�p��<q�{�7�ݲ!�!��1];�tj�"�Gx]���# ��t��qz�xg�d��7~��%
@��t�r@��l�'���saqR���:�Nh�O�n����ўIUW������k�֚w�'ެJ9�W�jУW��4���5�
�.�I���Zx���g��I��U����:=y�C�w�˲U��fv=V���S�WZ�a��Q�B��a���L� f���[�/L��܅g�qz���~0r�:��b_�V@�v�	ЧgUng�q��r*:��v�0\�8SR��{����|$2��W�OD�GSI��x�|�'�%Ԝ���aW�J��r���&������~����90���r)z��1��H䬢�p�M׻h*<��Z�!��i�wޤ�Z�p�����V�[�Q�HU$����"�N�Ǡq�����̍���M{׳�J��OnY���c�*�mr�h��!ݤv��̙��5#*_�h<O�l%� 4�$QAE��Nץ�je�ovoX�^�����͵�/Aνn���]s��bR�
<�|�,�EaW'0�P��!��}���M^#״ �20`�m�L!:ߙڈ�b���[�o�K̵2Wl��}����Vټ���uK��L`�]��~�"	�IK.b��jE{Go׋MJ��^����L�;(9�C%~k��Xи����72�ң(��tI�p�-�sv�Ƣ�A������/�"�/���0���ݩ55K��I���m��!gf@��+T�8A��>.^�U������xA:�`"�ݙS�;4!�xQ��[ 9���7��g�����r�Ml�ҁ�+HC����jH�X�?�u�.�К	�<�5�����l�1�.��<���+r%]ݱ�����l7�W���|�����z;����@����nؼUeH�@����H\���NTZ_1�pԪ��`�|`D�5(O���/gl�Ab!�e�*��z ����leDLE7x0(ݛ��EH��3O�y��g�&t����ۧ�Sw�BR��\��dM�x�{�0D��ݹ)���[C�ɘ̵�q	�U�Z�,�~-����D�E���ʹ�E~ɶv���F��%����Kǧ�{�̜���I����8�!��Yo�~Iߕ]%��\ks�'&@t8�Hi���X���\w�����ͽ�Oû~,s�f�F�gTNO�F�D �"��Ϋx��{�;\e��ֶ��e��gI@��7+u�V7�=�5�S皪��Q����T�C+�*�j`�+�����F����Qd�3���I�yص ��߹��'u|e���%&5}/��O'�b e�kY�]�J��w�����ȣ�S��/��طo���&g�H9��Dۀe��U?��]�s/�/�l���6�����qǟ6eȽ���",Hub|b�����3c1�nV����L+�\�~�#ΩB�߿	��A@��x>i�����9�Rĉ��h��G����](u��G�x뇶�کd���1F>���;�1)@��a�?��*AS�v2�[f N�X`�(Gv�V��6�>�<�yK���%�-��Z���_ֶ�2��`���^��D�oҖ�˖I���&���<2:%�,�L�ڔ\i�a���KO
�x��i=�;��n��<�c8ih�No�^D�I'��0�t�+g��i~
�ȼ�����.�/�[4�J�a�	^�?�r� 3^G��Z0nA]?|/�{����r^6g+{V�i^I*��X���}FG\�Ci�#i�6�|U���!�P\�w�r����"�y��38�m`ߎ�oe.����:��U�"�˧A�b�X:.����@�W|�� w�\G��Z�/���7E�S��#BSa\U��	T��j�cj�#�W^9,m���[�q�_@��i!��h�\����s���gkpJ���Ǔ����{R�D���Q>Yp-�+B�#k�)>��6>�����o�[)�A��P�J}�v�Ca�ͬ�0Њ��(s����q�ɳ\����t�kV���x�Y۠�_?V��AU��n�\ÖA�uStBm�B9��)�G齩���%.��n5+��Z��Pd[x���Z�ru�0{읲=|�Јw>9!Zzn��T��w�\f�[#�c����/ִ%RT�ت��(S-�ϕ���VK�L,ʳ M]P��~��]�˥��A��Ǝe��6c)�`>� yXM��@?9U24�����"�
˦��P%��~NT��vF/M{u�T�O>��1̌�p:�Z%�`9oe��SUNd�+�%/����j���ApٺS� �L~I�LQB�{
mzo�x����b��W;)�I�C��h��+�ŸP�k"��5����>�@s�r�¡�u�(�]��XK:�0(Y��y+����� 2[��=*�?Vj!��tD8/�KQ��P�H�	������s޹��y�!Ok�`e[��&"����80"ЬϦI��%�}E����vk���x�(�TM"T`�6�l$4�1NDK��@h�c[?Zw>n'7�1���Ǟri��y�d��	>��jq!&lX����~`��~��(��M��LR�c�£%{P�\�o7��B�˗���,ǥqU4�Z/�YI�eG[l��<0�¶5�m��Ekh��D�u�iY+O)G���>��:JB��nF��7��o��PTs|�X����&+�6��<��ߊ����6ߑ«���׆�9������/�p0/��n�����D	n�Y1�|㥵=�Bm����q��1?^�E�1�M5�t3���o|,1����Q�O �@�VQ�㋟U��H��vײ�
�9q�����W����N�ն���yp��k�L�W-�IR{^�Mڅ;!���Xd�}��,ح��r�� }�\��-տ��o�9����"�4ܼ�_^KRj0�%n��
+��×�m�>7�O��l�d�c���$"�x�I���iif���z!v��fM \\wS����s�7%vر�������I���LG�A�ʃ�L��J�`9��ي
C X��v�9�o?L���6>g�Re����x\�l���b�c����
o��
��S��\�sY��@K�D�2�dZ�����ׅG/���ҞX�9��NtP¤��}T�E�i��mq���Sxۨ�l�H;�_����������B+�����"[Ij�H�Lba�ײ�[�	oa<e|:w��LF��,w����*��k��ܴa�/V����k�6uVB��2}]^�Y�q���:��ߖ��(aFLr;����h��|Y�ҍ�W����R���o.,?/=���@6�?����c��*�c�(6�Ѕ�%^ �`��֜V�Sfڸ OCN����+�o��/�=m�h���*L�B����zDp�)��EC^sK����;t�B���Rj̙��;�Y�a\k��c rȅ_�b�$L\-� (%J�yI%��'d�6�!X�wJ;��kxbH��c�Tjp�e �ԩ�pp.���7q�C� ��ߊ"&z2��S�f\�[��&`m��}���T=�9|;��'��7�8X�|���VJ�ZCzxLR����¡N�ڌ5q���	����Bq�aqip^�vC�qn�Rտ@%I�t"в:@^�����&.ik|p�B>�k%F�j���0�;���i���?��n��	0-}do�}3���xflI����7`"�;��k���V��H���"|����D�k��@�j� �]i����0�&�z�TRVF{�������u+��;Gu?�\��n�A*�w��s[-�v� J>y E�zT���3����&�MW��mH�`ׯ?܃��5Z���eP��g�:��6-rW��ܳ�T�����6mAJ���S�D��K&h��w羂�����h��� �*�׮�d���b|pc}!��E�CR��C���������ťX� sV��-��gܝAs�"M����ZC@ߥ��!��C�amJ�{� �Q"�m�#��t@��V�D���Ҿc��"2�m<�)���lT�{�)���<U�.�S�L�x������!�%��AV[ٹ�r���G0A��j���)M<=���$�
�j���~u��6=J���LJ6��$�$E�K�m� �ܲ^�g�� �7ΰ}D�x�6{y�������8%a�_�~Nf�LS�%�ӬW�c�v���e#ۡ�;$)�	��9ey����`Ah��Ƀ�u�+�NHH��P��d���jυ��3����	Nڮ��FY_���
ѵ!�q���,�hTs����Qx�@��`G�t=�ZseϾ~m��pu��w&B��'�@`�-pRA>Ę=s��ǉȂ����*#ꦙ�>v����퍣6��7D���Έ����ϭ����nңc�5�gM���<���V�8�)s��Gݗ������G���u|Cwf��N��4%�QEJ�4��v�:��+��8��t��a���q��E���q�K+�z˶�m���%�f�**ߺ��T��F�i�й��Ѩ���c��[��Լ��_���4�#=��o�£��S��ד�5*�-���Ӗa�!3��.��h��T�X�&U����@���{��O�zc�}*~�`��ħ ��c��ʒ'���S�	X>\�Gٵ���z����
�*"):_i�1��E���	�UB��'E��}���-5����~Ԍ�B���y�v�7=7�Nn��k��VV:����#�L���k�Q3��?���z.�w78�xY��R$�3���*��^ص��k�d�	{& ��C�~��\6Ig'J��g �mK�-��[޸'���|����"�)�����@~1��a�*Goz$e�J�2$�� �ӭSOL�d��!=4B��SQ����� �<� �L��m;|��%��Ȋ V��d�;X��;��^T�f�%�g�UX���G�:b[�VQ��%Kx�o1c����Ɇ�����E���.�����:d�|zG�Mg���n���Y�S��y=_��f^Y=�h���@M]N���� ��'ƅ��^�Le�W�,FCM���3"��
�Ԑ&4��j�DuDi��L��9H���X�6)�=c���x*A��S���%@�=��H\]ox��Q1AR���(̦^Ɵ:�awv`�V����Q�`�5��y�A����aPg���և�"]1PNW���
�7���ɇ*`�7Ɣv�O����dQ��Bg7h��,�����GC-<-u��?wa�#oQM�����X5i>d'9^>���_ԇ�X��!J
�K�n[�6��.�kO��!Nُ��,�l��[�Jx�J^¸@���'�}5�"�&.K�.��/���%p��,��xR����XQ!��9�w(��C�&^p��������p�I^��em����<�]#U�������m�#|>7ߗ�ϯգ���쏾���s,f?WQ�+��9}�N"%��3Z��Z�Z�e�(�{��>�%�+Q���fCS���L(J�5p�;�8Z���C?0��ZJ޽�<y�9�Oq]��MK8����U�4ء]b���������4��7����W�R�g�M����0�MB�Tf���z��V�!�%Mp�Q�2�Ն%��
�AܒSNq��<x47�y}9�Wy$aXP#�ދ�"u��G7�O~�)t�t���b���'�?�Y�nF�8t�R∗��g��{�����B���;ݴɯGD-���(��)��Ŵ��6��5��h�'8d���jx���Tۼ�]��\������MHoo�&��G�y�W�}z*l�כ�(h�<[��
���j
j$�n��$'����1�_&2n<]��R�"�������v~F37#��Cj���>Fr� ��a�9���Ӵ����^ݬ`�X�aD�t�~���t��.b�RC���Qo���/�~݋W��;- ������4K��H��{�ZW!AA�3��_�7u��|������o�g.E��b�����DF�7]&�S�傿x�E���p+ �-��w��{���Ev�hJ��I	�tNky�� �ԯ���hc+.����رD�5�>�>�<���"�u���p��C{ ��T��UKw���Ɩ��b�#}8������.w $lcލk����[&�-���Jp/��7�9�bC�-x�]U{K�*E�xƨ�p����Fs�ݨ�.B�8��hld��Hٸ��y�_��?�XQ�]�	�%j&�h��)B{�Hn/��#!c�=��H8�i�_~��G�W�SFG�����F��YS$�c�5�I�v�5���y�V��	Kf��&��SfI-pe��X��i�T�)�r�t�nj,�\��+iJS�vR���x|�'S��Fd��������l?���G�ē<��G����V����'̾���w2�x$�:H��ŭ/��ܺk�9 (�z���S��1�Q�U�N����g[C�d��ƁV���R3���lU&�A�84\C7��ڷ�'4}
�g�l*jO���>���Z�w���|hQ�Y���`��(���ݭ#�� k�B^{A�W{�-����83���E;l���^���bUEi�G<��t%�Y�
��@�0�J>Ox��F���V8M����_c��M�m��=1q��!�a;�G���P�T��zwrU��JD(�^�I���V���]{��9�ޒO�y�k��y|&�3��e<�|��!����.cPM����$�UE�]W�^]2g��F����㡽z��7b_=�� e���L%8��'rTS4M|�8��$Μ����"i�h��-��G�ϒ#w��'ీ��l������BeVi˃VE"�^�)�J�i��ʩ����I�:L���?PCL�k�S���`lȿS��9�C�a�a�������/KF�(�:R�#�P�S�?B�k9/,L��V�(O�E�I��7��?��u��0y����V��zz�� o�$�aκdiA{$;�I���m.�)Le��_�W�t^G*;[[Ӈ�\8�w{M��#N��}�[%��m+�׽`̻��xXGSH"�A���>�;�9�����\�?��ӧ�l��_�ȔA���.8�ቔ�y*�ʘE��i�;������v;)���!q�4=�9�Ȃ��{��̩:�*�>�
�ص�D� OW���R׿��a��JM�L	A"/d�h�*��8d�2G�0a³�� ,Jvy�N�:w^���dð��lR��
e���i������*fH�A5H ��EZ2� Ц��>����T�tf�6��S�Šw]���L	����휻���Y2�f+X�8���Y�^��ԕ�\^ݚ�i���k���&��Ҧ���� 	� ��?&�F:���Ey��V���<�ֵx q�p��t�>�|y��ia&zF�W��Q��������ii`�#�ܦ���9l}��V���!h���dc�BuA�Ê:e��������O�l�s��?|�bF'� �Y�Gl?�Q_�e �/Y�2�gX�Q�t�T�ÚNZ������`�/��
����b0󧓧I�2T�ZF� �W������Ա.�ʾˑ?��+�%;��
Z�������K���X�|��CYJ�#�F�@Lצ�d��Yo7��By,dKp�����$p���D�^m �I5V�	|w���^����/�J@�]v����X�f-�Mc{�6P�6���N�̰��Y�7�|��/�?�C1��*�=K�ц~M����&�J�sK"U���)����c��J���+�^���/�N�ô&���]&���*W �t�0J�.|�5�V�xk�%%z�l�\�[��+�m��W��J�����8Z����+�P���-/�t##�*���-�8�OZ��MN�{7 ����y+R��O*ji@,daѧc�+y��:��׭��@�!L#\ϓ0B/n�eh֠)�� �+�BԶ�*�Dn�>Ze��#���Bݧ�ǜ0!-�����|�r�uS��7�z��<����e����;u�m�!2,%A�[m�#Dj�l����@V�p9���FXh����5�/B��#f�R"�����s(���ij��38l��FG9����(�p����Z�ӿ�U�>D� ��j��~��h})ˁ�]خỉ����&En<	��	��-��5�}s���{T��y�r�u/�ge �9��l���$�R�RÛN�؄p��O��%�1G=��ε�	�CY�Cݚ��N���.�K�reA���q���`�uģ���
(Q��|W
��[��y�v��"�����hJˎeì,��e�m����QqH_ ��&���7r���}�6�R�ՔD�Tj'})0�-�&�lW��a�h��K\R��G�'c� �~{xŘ[WZ�C�Hڀ�
^L��^��R� 7�3����7^��ȡ��V�`��ϙ�^��+��}<����?���7$��X�!����m��1���V��j1�U����������Oo��+�u�0fr2���@��c�d0sI�����!ǖ-���?J�ԷEK�V�اǏ�\�0�n�y��"�W8[�6y�(���	Z�t%x����pBS�n�[���+P*C	,n!Sn��F���$��jFWe���x�����sȮSA,�{��C4���7d14�p�&����j�a0��	T���#�dHXd�L�����jz�:,���߿����RNJlP�c?�$6�La}B$أ8�)�7�����Z&�GT�|I�/��:X?�P
ҟ�#|�C��=k�	࡙���y�=O�J�2�UfC{�$e�*=����.V)�R�n��[~�C^�fPе	n }�r#�
����G�>{w3�/4���^K
�n,�mmˢ=}O4w��� �� "1-7�[EF�A���V�۽��_{Jz���2��U�dಊ�s�V���16��3/�oݤ%���Bc�Wb�N� �nsl?�H��R/�6�ygjvϗ�U����K'+�;a�Ћ�azd?��m�5_'��,��2��Y�P�������Y۔S�_'�E�$��"�B�.��&��7�S�"��y�RdvW�]�ַ��*�8�/�8��I1�{�o�4{����W-}��o����I�Z�/1���GC@닎"A�"�A����@��[\�����U	F�[Q�/����\��#�m��RI��M2�/V�Z��m@��h� quY���ew3�o/]�!H[��X�!�2��Thk�]��+d7BH$?�H�Ѧ�XA��.2��>��J@#���є�jܥN�ϫ�:~o�X���i���f��m�>Vxx�`����J b���m�:��D)Y�/��ffK�㍆Vx��~����b��}���)K��o߈�v�|�=�J��`h7�##y��������f��Y6���6�HF"C�����T������E�����S�E��]n��Z��UF�y@'�����X{A}:ŗx6�{�����@t�=8�䋰��K�}���'�u�z�酲SGVѧ2j�>`LyBNV}�(����|[Q�_�����RXh���)9��%��5 �/�e������ a497[���T9�gA��duO��)��蕝ft�&W��w����pϻ$sY�	E&7�����P�9p��{]�kݷ�Ȭd`�k�� �<Ƨ��5�P&:"�$� �����̛�0= ���<� ��8�^D�d�F!�̲��r��uR����P j�F!�%�yYk���+���L�C�D#M7k8R�W��&S�$,�1Km䒚1�b��>Ϭ\<B�L<�	OՂ�ÿ_)o,QbFs�����������ϫ%�EƋi�'Ed��C��ɇT3����f����˻_��l�ѕ�2ѯ�ֻ� <��$m�E�|��8�Ι�%�m��=�9����/�(~K������+.����1yX:�Pڎ;�@�Aw��I�����:�)ro!��+}�����,���L���V�/�v\G�ӭט��I.��>�q�W���u�4@K��㔣 Wv��XfBj?�%�#X6�{���n#��"ٹ�|	�5(!��iu�EP���E*aN[����]>����Ԇ�����j��kj5� q���M���GTڥ´v���1�E.���\��ҙ����kR�{�OQ���}�p�����C�T��9d���
iſ�C������, �Rj���M�z	�@������`�.s�Q>̀�!1�x���&�_7��Y� t/������תym&�W>�&�6�օU�)�� EAL���^9i��\�J������X�[W�m2'³$��������������@��������a�}L����#p��jj.Z�>�[m��fV�/��'�H�H��Q���4_�VG�"J�s�7̝��Z�X���3f�T�C�y���o�Q�2����z���K+��+�)����\n,p9��
<��}B�����"F2'G#K`�e����l���^�m��3p������_�eu��y��<G_�J�{3�w)8�_3<�9���/t$e�XU/�(�������*������e=*N�ػ�}�(B��ʀ���z����Z#Kl��^�J����8�s xw2L�������`]3���5O������"�#_����yuw�_%'JjxѰ�F�YI`�GPO!�>�+ݣ[���_	Z��s���7�p�j�
�+i!�� �J��$p�O,���Ѭ\3�c�`�Mrr�=oKp�̎�����B�鑭+��
ё�����K�x�;���'�!f�����/v�|-Z H��vN�<�N.˛�!S	���"c��C�9�G��P��(�N-�u
b���86�w�B�Q�Qx���nQ}�&�s��ֱ{��Ѻ�^i�W����d�F�vF�S�U����?>I$��d��n$q9�o$�nߠ2O_S�yh�⹙ �WL��m�ڞ�{����*g¤b)uȋ׭��!�|�k������6�fj��2no*�^��q�:��ͼߘ���	m��s�R�rӞ�7j;��-�/���y�o_�>��o�*4��Kլ���ǵ�S_s¯G�d�����$l"S��7)�ͪ}]�3/k��r�����r%�;�lz�vB��`��#�5�Ʃ�b6���6�:�B���m�&1�Z�e-'K/��щHo�o��F���Y��6�][����μA���2h�_I<Ɇ��Q�����x�nQ2�e��V�6L~#O7xw��,A��`g���hye^}=���gT��D\{f�Sm��?�ٵ���P�Vթ"��'��[INh�AE�VN�s�<�j�����d��&z���	� N��?�Y��絁fR�Q���v�E����gr�Xlއ�F��|�E	j;i���w5�ZO+i��uo;,��!��O�uL�����e2�`��-z���XǹBq@$%'3�����Ho/?L<�4n� 7-���X#�6�$��H�+�f�;¡�4��q�)�q|5M�O,���'o�)��������A����K��؄1����==���/�o*�v�w�[���L	�F��P$D��#2����rSx�۔x�C�׺&�#���V�@�bY�mG��Q���xV�, F�dzj�%Y�g���W�H�̬۟�J�D�����f%�.o
6r�9l�-����j;i��2���������.�xA�U� N�) IF~C���YE�aŔJ��Ӌ�PB�lvԜ(���~,��؋�1?o.�������'�Gr��ZjT"���H_cN�P&d�ra�GtћK_S�'&� -)Q)o	�ʩ;��� M���m5�:�Mᔳ�s���O�4�A��!��e� TCVͳTc�|�|��w%���ɕ��o.li�q��Q���0|Y�4I��}��v�C���`s�ː�h�囂�e�,�6���<�W^�Q���S$Ȼ[9h�@��:�1��$�ě����P�D��
-��m	lfgJ��0dN�2�;L�\2P@PIɡ�oԉ���)BW�)TD4|Īl'��e
z�u#��+X�U�^�9]<!W~'Lt_���0۶�[X{2��0g6:L�']��6e7uk/ٔ�<Se��I����IW��e��J�È%u�_�P�2ՠ��Ɋ���*Ck��Yj�������n}&`1��6(�2WN,�;H	�]�����#�d���nME���Э�|J��T����8��u���昭���������!m�n䱎�W�;���cެ񎨥��tE��Ë<Ԋa��W��m�����ڽWG��_?�ib'ª7���v���ܶ�������t���T�-RE�z�ٴOm����B�F�*�A���.�� ����t�SŪ�p��Z$_$7y�{�<:fY��I�Muîd�����.2�N��~�����e�,�J%f,3u��~gs	"F�١�v-�ܔ�o`e���RU���Kq
�1��R�h��u���N�G�R�"O�(�>����u޿�,.0]�p\�gx��Y�zC۽��qp�I�U��47?3�x�_F0(��Z�����n:?�+�i��8ԙV� ^>�\�,$�L}�u(K��ba~vC�%قm�p�����N��';���Fk����+_H�\�;@�`����j�)���H�vb�|���\�V߾�ܜ���g움�pr�LU
(B��/C"�%.4��qY�=εqM��l��0t���X#&�tZlá����ND]�s]��!@ ���بA ��ܞQ�a���\�J�F]R/:�����T<����g��"�i�)S���'r
f��ؙ{*�Ns9Û���$��Lː���ꠐ�a�T���pJ�p��r�zȆ���3ټ��{�6�8�c��`,��A;�N����@8FEN�n���:�P�e8�45�Å}I�'�2xWIo�QȽ`�y�=I�NV?C7/Y��/A�q'l��!"`9"I/<�D�i@r�d�Y%��������?~�@aO%�[gb�w�)xH�^��
W�.	f����.�B��y�et�������q�zW"K�G,�%G��M�)I���,v,˥�UkO�pfiƿk(��aDg�t�Z?x�7N�Zb�-��
-��.��D�n��w,~!�=���Y��3p0�d�����̦��C����r����T=����u-8�Lb�,F�{E���1]��F�<����|���0�.�)���[@�ӿ��㰽�����sHԇәx[�+K�[��W`�6��ݣI�����8���]��P9;R�,�1��O���M;� ���6.q��+#Q� ө����U9N�xʆJ��i.�[����/+��-��y�������x�A4��$~���7w�>bh��m�G��7�m�uR���0�C���q��뎃���A�B��T7��ӵ��aТ&�#w'g�$������&F$�	?�q�a@o��@U�;kb�����L����oZB���m��V\$YEb���kl��3�w�`3�9IL�|�%�8��X�F�v�VC�-Z�/�e�#����ktw<���{�p{_��fMۗ/�)9�l�d��ĐǑ���x���H6Y�t�:�$�Ō��92I������z@�`�?)�O��s�1�cy+[�����FV��L|���A�܎�KG��rGV�̽�7�8oc.�>>�X=/�;R"�j®\��+&i����Gq�4����W���)?(���-�I_EM`,E&���#�)��$9I4�Ҥ+�&��rz�����������e{ub/~���:��?��ZT�V��,��7$Чш�6�"�ɛ�%�JỘ�5Q ��#�P|�c�6F��*Ϭ�G �&`8vZ��mS��ʊ+�d�W_�0hG"���w�(�>�,o	��,&�U��Ds\L�\b�}�βEG;R�+Sp�ܟS��� 4v�zV	Y��{ ��D�"1R|_H�;�0j �x�Us���,��oW��~.��-@�5��TϽS��/�MYf亙���yI�OWMIB�Ų.�3���-��\���qJ��x;O<���=l�ֱ]Y1N�e҆�$[�H.�ׄx��D_���*)��)GZ�`��ߊ��c$�fya׸��3ҁ�eX[��I��X!���,�Q�=�B:T�r��2��(��`�2������kqPFE�Sn�rK���WS2u?p��tA���F0�����%����>]�[�i��MYR�ۚ�}PCF`��\o��MΖ��	^C��*KS&13Jvq����u�"���4��:mM	�d!'�fRC�h&�Oq�L����ūR��\�?��?�[s�������4�"_4T�!<JI�,���5��Ӭ.cJ'�rq�	�w�����(o?�?��Q��Wɤ��J!Ў�F�r��db���A)��t�+?�=6���X�]Vɰd������-1a�K$a̓D��Vٯ>H��-,L�.����7܇��LSWU��"y\���W~P�j?�u~�2ݘ���m
?��~��fZ\� o�~�N�}��o|%7�U��(���5<q�������~}bu�#Yi�v��*Pޟ*o��/��o>G	���l�BR�#f*�c Inײ�b���?_+�Pj�B:)`�K
.�㡯��8��e�Ȋ)�
*|iطL��H�oIZ9�6�1��J�����F�dg�5�]�~#�4���8�5��׬u�m�0�ı��%�L��W
�,A7�I�#7��fR���Q�)�4f��!o@�m����aV�2�N�/�0.���� @�qƸ�S�����̭�c����|��۴���Pf�ĐB�b�j� �@�d-M���jV+\�2\%��e�A����s{	CB<Y� �Z��'(;����@�%}A�[{������<�4Jf�@w�u؁�y���9�c�jS G��HTu驠�H�cM6/��6w�4F��G�ȍmIZ��c;��w�pg���*OR��m���G��QI):�J�� ���-H��걃�-k�{B�͏Oۭ�M��!��}t@��U�����q7�)F���Y�wuC��:#�J�Q
�]�� Nr�Q	Z��қ��
�t�\;S�ި)�ˉP�?qϭz�U��;�s������'T0�D|+