��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�=L��4�S���J�7�h��J�3�_�������p�t_3�ѹY��S�!����_-)�_�3s&�����T���X��)���� ɋ�-D��VJ634�x	�-c�&�Q������.������n�wz�b�Ǖ�㮡Ҵ�s#�D�P��&�tU�h���H� ~�V��h�K5F�av�N>#G�qm�HߟG�!Қ��(ȗR03'a��w6EQ�p�a��f&*��F�=��sS�*-1̩��٦�ƹ3և{b� ������D�LL�003�Z.�yj!rV�=���)Wz����U5ၳ'e,)"2����ѡ� ~F�L�I�W*u�B��c����:'�G��8|T������&��m��twπRl�<�5Y�/��B�6������Xن�W���Ys��l��k��~���S4���;�� 񰼪1c[�r^N�-��2���(O�.v�c�T��"��#+>�4��uQ
9�ٿ�{��$(�Y"�ƈH�tG8ua���Ņo�h�Ijd��u��Hrw�7VA�ZDi|���`��#Eibn.���ӫLM���"��>�测��zK. �ޤJ���}�,�$���\R�ÿ��s�3�>kڎL�PX������Dں$  ������;Fr��>�L�T�	��42Y6t�lZ����zu@n$��R���5�<_	P��+Z	r�}�Q��B#�ף����b*@ᐏ��^���3'��W	F{����=��p�X�\6Y!\i����=X��qy��U�|�Q��`)���V�!"ާ�U����@���Daş2C$��j.��_3�w��������to�*<�ΖD�Y���Ӻ��A�`3&�0i��̋����`r�h�:f��Ԑ�([�%sVi�p��@�~�[4�?z��0]4[h��6�ʵ�TN�������z�:�G��w�ps���n\�Q��5]�rg
[?Q���&���ZcE
�����P{�h3xX��{q�.��� ��\��ZՆ��&��w� E��n��ė���^�;�=�J�
پ�b��y��ۺ42��o��+����������J[(������bZ�K�:�S���s����жe���7�s�r�� '<C@ĺ&�^�,��g̔�������xo+)I��j&mڙ�'Q2����ā�v�.��sL�^�Ś��9�:�؃H�S��eWe��h��?o���m��Ց��w����d���h@aꄟ�K1zY:���b��m����'�s ��5݋�J��Z���쑞��i��4������l�ַ�e�Ɂ:����P-�j-#�����DX�b��cq&cC���qƂ'�:��VC�jV�]Bå����Iz`E ��۲o�Ef4=C��t���ܑq�|�<Cw0�%��G=˴�'�2>.㍾��ila��*��	j�������*�
N�������Z΁$��o�����.w�ZF5���m|��7�צ��t�P��Θ'k�"��'����`a$���R����~���I��?i��<
)Ϟ�x��1�<����N�ƺ�.V�|_�
0-�T�ўIݒ���z-�9�)�N�s���X���[v��
6~R�p�q��e�@��Y4��7���\I�����*��P�B�L��M��g�B!٥�b�I\�����z@n��Z�_�;�^����9�1l�3!���n�������m<U��yĸc8��LX]aɹ�x�Z��Ѓ�MsQ$ U�GI��}Y"�?n�j���g���4�˵����*����^���^Y��I�}�Rk�s�����A��x��%f/�m�M���^QQ�3����v��Xַ'P�������y�$�M�[���^�y����Wi@_H���r�-��>�埵�����}~�=�4B�|����/��.�s����^��otL�W��N{WC^c �:�Q�J�
�?f�	rt*,����=���&�~�΀���^&��^CP��6��#���Ci}	����V��� ������u��L�H�nK�=_�J��hZ�5�"�_fP��S�ˮK�/��ܫ�˿���z�=�A��QR�+-��G)���П��&�� 3�u	����u��]�����ͱ�Z����;��(�=ɢ�{���k�A[�/,{�:�)�kd�eʫ�Z�]f��U�h�R���� ��_���#Yz�G^����:�8'��IH��+���[��}|��JN8G\,����6�P!U}d�htcpW��� O�<��g�,�v�ƇGOj��.��>����]��Jg#*�|X��qIiw�F��}Il�z|Kz�:81�T���kl��S��h{����M	b���;6���-B�`2���	5�혆*��@��[�X����x����l��9��ĐN�'�%z�q�w��|t�\=2����Q�+r��F��n�� zK�Kߺ<��̯���A+3;ё�E�0А�b�ή\����Z���Ǟ�%D!����z1X%��j�ӅPl��p�>H��ý7�2������l�e�*�a���>��]`	�07Y����'I�&N|���_Z$ ��t/G%$��  ���#GHT��6z�΀�ĳ�@?C�	b��%�̬v8 ���hj)�g�wY)t�}�p�썥�]�H&�����Jt�� ��Pb=#O�r<%0+�6�!7��W%$S��Lj;1����/m��˻�53H���_��Qv8����˖�U҈�c� ���4N�k�x�'���|���\��'�\bjqo��Z�51�OL[�Om7/y��PÉ�9N���d��,�l�2�9�Z3�t	������z�|!_+]�N�ݍ����Cq��F{��:��x���Ys`���YW� bͳC�\M�.��)X����s��c&��'��1��U��D�*@��M��S�n�H��(�b5J:�(X5"+l���D©j{�~��/���c~3U����xE��m�����9�H�{M���;�\���n~1Q\��i�ͅ�̟��nmM�>��9+)�ְ+)�+��a�8����%�������a��yo�}���6A�I�p�����U��ɥ���V\�m6ЍiqHF+�p�J�>v�D({�q�֦3-��J��j��(,C4Ȗ��%x[���j�ŐCcDW^ō�t{���V����lJ[Gi�	8Y_o{�N�C!ՠ/��۸�(�}��Cqb�_�F.M�9�$"<�.W&'��!�V6�'~��A��Rn���@g�/�7�Toy���=ʊ�FIA�NN3Y'r��>��N�������p��wx��?���%�U��4��3��A�FG��þ6�}ZV�z�J�Mٴkpss���[{)G�G+�Rv��D�-���a"H�n5��,s��V���If�΂TY6�����2�D��M�>op'%Y�!@|�,�����ߝ�p�!���:h����u��e�~����2Jl�{����wp��qo�a�����&���Ǉ�p�ם���u	�}߫CG-@��-{���=	d�X�t����^v������{
|(�qd�{��Ll�I�p�eUQ@ \9?۠�"����縲.��ɥb��}V���'E�V�9� 3 ��Щ�M�)��呋#x	W��M���ўe���a'ʓ�U�}�*�gz:��v��Y؅���?kt����z� v0���e��I��H?esVF�kA���sLr�����g����o�P6�L��l
JZq�K:8��Fm̀yi����c}�`u�P1�:m�[V�e��dt�(K��߅���~������G.V��'�οeN��sܭ$;
u�;�}m�̘3����c�L<�0^)���Lh���|�5V(b��>���O��ͻ ���NU�Z{�hT��M)r�9fA=��zr�eА\JT0L�^����8����p8PX����6X�0� ��o���R6ه鿀?Z�-5�\ ���cY�S��U�5����L�29 �C�W��2*�:��?aj�hX+��@(a]!h×���Ǝ*ѹ�Jz#�)B�C܎�~���A��r�JXu�P�Er�s
�N/��"���k�����Q���w�|Ll��^��
��GN��� ���i< �jXPԌ|��kM��i	�m���0/�J��oqk�����;8�fF�'$�Q��r��)�슃�fm��Dw�x�S�7Z��-\��٠��|��h4_?����dH�����i�H�L��׸j�)Q����C����~��.u�V�~_ҋ{�(�e|3/w���ݹ��ʩ��2�7���gi��P�S_3�n�#�6/���Q��lpK���gD��)��Ç%��2�_¿��f��T�l�8��1t��_5�/_:�˴�^]j!K���#�s��ϔ�� 	��m#1�PӃ�<j�2��?dc8iK}�2{��f���
6P0:�^ʦ4$ʎ�+�Y�s��(�!샘mx�#�ȕX���-:]�e켥��V5��E�<u9kv�!���c��T"�Bѣ����]�wŝ��)�lU ���wQ�;�	�m����ʦ`������<�~��7�;��ޭyiq�s�T��-?�7��)���~z�G�'?���]G��f�fg�����4