��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���ڿ���͛�BEx��3e��g/�s�M��\�<I>��@ꔧ�@R_>��M�9�Y:&��P���#�#O�yM����A%�Q>E�SH?�YWh�&��˹�2���b�ab�
�V�@8�{���P<� =GBU�u�ι
��x����pF������=@�@�v����o��2���띸m�d߱^��zK�Q���B*Ӯ�`21+�FR�N���Y|
��t�1^��0fQef"���)�:��(�@���6�^��^8�JJ+FV�ղ'���η�S�j���G-�j	��P�)������G�D�(댷x(����}o���רE�6U'uٝ��ێ�}����me�{�A�TĄܴR��"�[F��v,���=����K��'�I!>+!_a�Em�?�kF��I�(4�S�Ѡ�A�������,�,h�N���q�
���4ԖuL���v�+���D���؅�YD2f�p��1��X-���s��������"J��ߞ�.ܷ�'!O�[L5�(��<���`XkDڷd�^/ |o�e��`�'���:�|�FW�^|36b�J�~���B�@o�u�vE�s~�_Mkc[�j$BƉ�F_ے�#D$Wc�Q�%�$�ʰ��T�:��a[\��kŻ�Zf�ƢJ}��,��������fm4R�.�@����I�ݥB ظ����?�NWA4@{�b����mQT�9t;�I�.���p�,m=��H���s�NK=s�?Vv��Mjw"��%p;m����1IG��'�D� �X;���ä�.ݼMGX��h�گ�?N��";���Y4�#��Wi�pJW/W�H�Ί��LlP�&�3�d�	Q� ��}+��D2uN �Q]������fHɶy�/E�]r��?�)yj���Gλ�C������t��Q��O3p5�����2lv��x��&�C����F9�iw>7���Be0���H&�J�:�2L�����ՔL'��Ϡ��8�C����z����!��ω�� ���n���%���F��a���0?,$&�<v�\O�"va����5@�t���ʑ~7��i���E� >քb:o5�Ń:��A��4x���M�g4-Ʉ|��5��B��!�e0\��O�H�}��0��{v�Ded+ ���B,���I���,�I���;=nG
�0(0��R�tJ�iL���P�������b�x�A�?*ȕ��G҈�\���e��a4�.�Zf�K�`y�0�+�v����L�@����<c}�Sh�&D�q/8�mV}D$��`�Adp��~�N;`d���(M;��o>>���,M0�(hx�Q(�x�(�0˻�ł�������I��U>$�5Nd�(��+�7�-N@X1�(�:�+��I]F���x����[���;5×��c���j�� t������BR��9�oB������������Cs�F��4;��Q�{��Ο�8�Ò��T����2��T�� ��P�9����v���Y[U���,���kI /w�D�c��y�Q����#�<��f�i���b�6�d����i���6�ϟh�A-'OJ�@�-	E?��DKE�)���S�9cɅoh��N(X��="}g�(���1���{PȊTA�
?�c���M}�S���-ۢ�\�������&چ�H���,����UX�_�_^0�3?�~(O�IuԊ9�$�r��* "�8�Ϛ�x_g���!���%+�M3�����tb[c�$�~���@dY�8�j������-KZf���]��}_�1�����7���c��؉��F��k%��l���d�ݛ�(������{�ne�7�� ���9�f�-�t��p�|
!�[q�3�
Gw4�τwr�x���L#�Z�^lPf�74z����6��X��q����(�ۇ�U�>�1XX�Ø%������H�Z�z�cwBy����#7j��ꋽF7����rl��S:���C�42�����a8�Y�ۛ%K~�v�eX$x�����&�ƚZ��i��R�sM��֪�U�;�קChc�y����Ô<�b�F�+(x,�IX�f���9���D�7��㝨I�����?_�<����AG<P[�}��|�&��֌&@ dQ�+����t�n��/��G��T��z��mZ� ���������/|������g%��}��V3h�?�@�C�Ի�郖IƮ���ۇ�Q���;�
��[�BS�4t9.1��u�\�S۬�&fu9�hPL][�"�B�hA��DȤޜQP�q��.odz7����F�	��Y�I='{��QɎu[�e��ʧ�0���l����h��X�/�k۟S�)�s���-�'�٦o[*O�8�uƁ�;�v�x��+'����Y�����k���a��QUBRQ�M8%���9�1�Oe[�_�<��� �h��1ZL;��P����,�!�����^�P_��R���`t$ߑ�Kh#�D�@�Ś�]��e�t!�;g�4�8��暑�v�֠]eQ
׬#�t�'� 9�K��������'>�X�e�
L��,�)q���\�o��MN_L7�#��/�Ƀ�.���O5��������8	�I��;"{9fj����g��*}	���co�_���rpP��D����G��h�Χ4y]��<�hV�+�}���#f�&[�8� �I@ቔ��B���F#bnk�稲�2+�kޚoG43�l5X�~��G-8Uf��D
aAO��P�6��x��O;ٷ��"4߲L�9�ڛ'����?O,���&qel��h�J�������Q�SŹ Tp�����@�3�:7��}���A\�F�����T�t�C����as�q���Q�z
�vV3�rGT|���')c6~��3�Q|����LN�h��|AY/m���Ѫ���ƙW�:�����K�ib���\��<�n�I����/��^T8�_gW	����5�	7R�.@H�	�s��q*�<��8Kffϟ��
��\��^�U�Ljm���k>�4��,P�r�%biߔ(\"tFx� K�D1{�n�A �r��̂c���>��1)ɲ���H,t��H1�+R���x,�׉2-z�6m�?	 |�S�U�zKH�&�|B�)��հ����̲¶o��ݚɤV��ȭ���B7�h����=��y��!�X�r���g�2�,y�u2���S���A�1j�6���L��6,fr��_-����"MI����O����ſ��=�N� �yj�̶h��2��~�Q����G#Me�V��%s� �}Z�X҅L}}�]=�ӠA�������#��0o��K���z�=�Պ��@=+�W�󨕩)�6�7H�;~�R�UD��}E2����~�����/�_�	<{��z���;�^��!rOx��0�u;q��9v\h���/��[�/3��E0�q�82�|$���e�`Sj:a]�s�0��S��]	D0I ��ћ�e�㛞m �F��l"(�5jf]L%\�ɩH�ܡ�p�����\C��h���m����)�尿��p;���ۖ�j�׍&�Fz�{Rt�����V��q����]���0+�53'�eΊ��[�4�S(m�V���AH���G�o�\$@s� �p���KM<������z�m,y�3k�1)�k)�l���A�*W�H�2s*�ÀΫT�t�V��9���R��0?7*�N4����	��{�,'Y<��U�v�#FLrX���g���b{'Յ�W�Bc�Qa����Q�A}��-�6}=N1�ӭ2��ϻ�����֧M�+��B}�n�����(�����`�=�í�೓���8[A��$��}��:P��J�0����t]oؠ��Yб:	�L��rS�H��@O"�~
jT6t���IZ��zbI�Ĭ}������l�t�vJ�G�t�/��X��Kn�pG,S��Vù�H*�_�F�؃��[�Bɘ�@���=������[|*�Y����1S ~�a�Hqɪ����u^bPY���1���$�R��V�T("I���zr28��v�5���g%��S�g��L�����C��ǟ��_ɶ�"�ĝ�m`�_X���7���.(Â���dL�u2\ ����~#�ʔ��mQ�N�s&t�ݾk��]U���KQG���d���j����ڏ�\��L��xG�3��S�N�"�0F�,?=��:h:����\}J__q't��{!%�D�3'�f�vG�X3��	��m:#�Y���&��d�넵�
84��A��h~��,���ey+;�`�����s{]#�Y�
N���Vk-Kن�N��v�,XpI10\�lݚ���LM�N�9���ͻ�l�ݬ����M��S�(m|ȃ��K�)pk�-jZ�@	�����C K-fн�}�"T�AH�U����y.��E�x&�f�i_��-px�uP(͕�&{*:��-fSn5�DUb��:�\��j�o���ߘR�".����v|	I I[{)_�=ƃ�A��ɯ>�g`3���p��m���JF����VX�/$�㵽��f�w��2	�t�^@x_�%H�8�6���fa&"8�k�gx������[�b]/G�~�#�G!�t��d�`�zv僀������1�k����Pt���a��O~ʊE׋�Ku$���wQܑ���|ZZ�^I���fχ�;�:�9Vv/w���ʨKr��)���&�M`i����������.�B�_��X�K�YRv�va�F��`	��"+�D��y<}���Q^��0�n< j������i�A��FgG�i���V�:p��	
����w[|�Pۺ -u�5�ڛcw�}�x�{۞R�;a�S}�'�.�>�������j=�q�*.䩗�\��u	��կ�X���]���@�����~�[@�b.B2�!T@��+��O/�q�{�ű��{��(�ǬE�:�.�<�f��1�y��e�ҙ%y�s!)����P������/��U]��[!YT������P�{�1���i��T�H..���
x6^}�&��ǘ��Z	���$�~#C�ƕv%k��|-y{x�̭5�5Ⴉ�cl-��J�	ц2[�O������	��
�ۼXXR�l3	VT���Xl�Vo��]M�u������vT2��#}H	�N�$��/^D�I������I�a6��9�Wt@G-�u�Ũ�&���
*7`���,�[?��2ˌ1��Z����1�R��H�ij����u����� s6��H(��`��k�E�;/�����v�Y�5��w�	�[����J��MF�>��Z���6"�C��Bō�o�F��i2�F��e�#|c=�Z��������(�O�^��*㣟���Pb��U��*K�E;��?�^%M�?\�U�h�B��W�i���7^�6��.2���wp�Ph=G��B����"n.����̱頭�Q��1$S�M�S,�f`�i�LT�o+�?hg<4���Z���D+����Zj{�A�y�fp�NK�Z��l��(�U��S��2���{�Fm�a!�x�<��|�Y�?nt�{{>�ŝ�O*�Yt�:�����˃�0;/�����i}p+�7c��B/ZwG��`����8	�딫rP<������3C=�'ʸ!V?�x՞(�Gڅ��ˋؔL�F*���Ztt$N����5�i�(�#�#%�fN?B"��T$��2�rT@t�[]�%�;�]k�
 `�T�	��1�C��y$fC���_�V({ޏWͥ:� }��;�bB�ݗ�i�/�"y����w���ӊ?�-Q��;ޮ|Z��ǳ��_=ĸc�"��_9��
ZW��*L4-v�|,�;N�	��"� 3XL�Ȍ�I���)��.�S����(;�l����&��M�H��F�wuʩ�^��+>K�(�\b=�h/�� �`I�5X+{a�<��u���I��3Ʀ�ѻQ�
�g�j����].���pI��W]=��X<�8>�ѳ(H*A`���kX�����G�k�F�����Nv;�k�.�6BP�:(Պ���}X��[��%B�J^P����!�/�6�.�k��GtX����#V�:�+"ͯ��M��w�=�A���]��6rl���Q�[m���(���qz!�����W'Ў�Ǝ���� U�&QF��.��C� ^y郌Q�i��<���S�6�I�xt0����#I](I�rq�ݬ=�g��u�7��ntL�8���
�ѮŎ A5�*���/E ?�zL%�W4�u$z>�=��x�d����"���T���e���1�A�f��4�$��� <*=�7;�ק�R��CY�l~rvʲ������z{��]�L��8ΏH�[Ys��4o�.+��$�����Zs�e,����3���$;���4N��$E�\OO%lm����wݘ�嬬�,�ς�BwG��Gn��ʌ_�LK����Vm�⅃���qW�7�������{�Er����!O?7�Q�=�o6k憳�o���C
k9�M�m�^�_F0���X��B<*$��0��W!��O���j��|�}�Iyr������f��TА��W%�1Y�*��i���������jÄƱ�5F,ļ^6A��Rr�LUZ�2a������JA���E�d��A���J�$�ݫHY�{Wf�X*JP���{&�57�
V�f���Ю�խ���C �^2� N�7�7��ۊ�d�2Հx�=��.��B����R�R?wI ["8ڮ�8��b�ꛔó��'�z^v�'$����۲:���u��V�R�Md�ͷW'
�1�cE����:gz:I��ϧ'��>xct,�+��4":��6��)��7�M���w}D҃>���TJ#�	������?���j�2�h�{nfj�Pl؁޿�� Qͯ]�c������"�c-$W���E�gV=�Nze�SWBx�n�=�֑:Fm����uksV��_���@�7���dm#����*�hdO�:����X9
�-)f�W��:���$�)F����<�M�M�0������JS�W>�������E��0z��Y�Aa ���
�C�>ߢ�N�e��&�D���m�%&j���vXv����d)u��o�t����� ���L@<�	�6��_�)�1� ;,!,i�2յz<o�����G2H�A	�͔���p}�E{ 1��=�}�x�DQbB�%S��5��J���]W�W�EPY�֖߬�p�|f[���{i�=.����-%�nY����{�0P��1��#3/�ٻ������<*�<�
/��Ǌ�X��o4�GT�jK �9�L�a�9&w�o���>'�֐$	�.�ǝ7y�zcb��X�dEC۶�H��C_�$���6q߀�~���ɝS�[`>�ZR��q0?��U^x�D7���V�[ՙe��}R9�����5�9QsN�G����O`"��@���(�`��t���/7cY��5s�t��Ix=�!�9���+<�-j�	��H̷�jF�ܷ�1�Hk&u1�V��y7:<4�S��� ���#+�,�;fJ}�¶֬Њ!u��߰vl��:�H��p��;�Y'mx�6���|_��l>����Q�,����ы�SY�����o� g�cP�OǊ��u�j��V���tG{���&��,��Io���X���x���W��hj�������楹���RW@`pٟعȡ����d"�(� �����t�$v��F3^DtX���P�T���B� ��*�
��(���� 6Z��9�r�Xܕ(<��@��䦓�J�yR��Ø�+�|#�n�$!D���#�=Mc����a��o�ty�TFܰ���)8�k���7�H�-�!�C�a����?l�M�'M�f�쑒�YLR�C:e���	[�?\�Z���ݩ0����V�MW��Fx�0�F��ջ.lפY�t�Eˢ�yL��{�*�节Ή�l��O� ����~���Z�uȮ�r�(?�6R?�9Ê� ֋�i�Њ+��zR�t� V��n�.dO8}H
�J$�v��,���ą�*ee*K��զyu9
���C9�z��5�"�}������{�N�h�-�?t����Q虜���ϰ��Ǟ�~���=��y,���?����I��=.�|�kY�u�@z���ⳗ��R2/��-��׿nBirv�.����RozQy�to�aeu�-3�Ӧ��,qw�#^���wU)������:@�EC�Y%n����f�g	m���Y�q����� ��2`��K�.A�A�b8�&3�y�����O]bL���!�3ȑ�B�
�b�xb5@=�'L���A.0�M�������me{��A�8�^�6�&[��s	u:պ�++f6Z�z�9�RY�	�c�0'-_��S���Ҧ0�6�C �&)��;{���q?�o�eն���C�C�B7+����ti�c�-�.J��ܺ����'�3��'�&T��o�q
riM,�T��Y���5/ޚ�K-g����]�h���iց�.��q�=�#��s&L�C��VjgO]4�W��4n�C�vT�&�r� +���P��MT���bv� ������"z���x�;� �jRe�v��-ҍ�4:D�[��;���r'��_��ǷrN�w]tj�J/��}W>�k������c��k�F"&��E��(�����}�+��$J���&��
u��JF��,$�e�ڢG��1I.%>|t���ч ��!�+�D|0�K�Nʩ+��W�	ċ�6@-W_L���(�^�>ߎu��,0��C�2/ɓ �l����V���c�(zRl�4�`��:���5���2+��-F�2�"O���*�oi�G�~�e�L����)�g���}T��W�󯀲T��2S�Uv��&�<�%���Mv�Q���P��:�)�(ã6�B��Fp�b0�Ws[56R�@^?�Q{�%aIG�?�WL���sC����C�L�Us������A��tn<B� |o0m5Л�
l�(T��䝡mM�T�O��7�G,ZvE
�"��6ac�z̓��w�b�d'��3�OM���Ψ�Y����T+
YӸ���Л4U�����f4j�9;��v�2�-��S�e�� $	Z���������;BŴ� 0(�/S�&	�K��xU��w�w7�5nWs���z�\��gȏ>��pf��E� &ڈv���s���Y�0߮�X��/�\�)hZ�0>�dDx�X�;@����8R�퐻͏.�C��_G�@����F��u�y��i�2_�/v�S���;L`QVEWiYYpK�<{c��F�� � G���n�� �
[B.� 1\�+���L�_0GZ�^�c���6�O�(�hMv*��-��R��.�ؾ�����]�0]�/�3�ȣ;��'\ѻ��`ɏt �3
�,���MJ�H7M}��G�*Sײ"�M-�����b�3�3�׮۲����3�Ԝ ��yhJT�+ș�ñ�=.��5>�Ee%
�N�= ^�_@��rct%F����:��q�I�ʀnM��7�`;�S@��ݪ!��ϑ��3�^&u����h�����V.�bB��2��ީ~�m���Y�<����Vy�_4��trU*����&���"����Zk���_ܸ5�����O/����b@T�)��p�t3��^��qWv�3B4R�|
!�;�e��'��yu�.3���cX�GݜֹnN���"�B"
�S`��tǿr6'���GФPg!�>��)۸+L>h���]�����M	���뙶����a�jŠ���a�E6!�e�k ��� �O�G��Vp�=�Y��Z+(bX���֏,�Op%?YM�v�V�8ք���^�n�z�<c6�Px��磠Z�zS��ௌ�.����њ�7m�/H�U]����'/3;��93��8ЇV 9��Y�Dxn�RVD` V����ޚ;��m����3�R�&)�A�z=�y�O���(��M�[XqU3ju.y��~ǯ͂PE>��|��[]��S��k���6�xsG5l5H�Ԫ��47w��:�\.ª&��d����d�-��J�	J�pA�g��f\��Ճ�`A��Mo��_���LŶ�����G�� �Mގbقv@Ĥ�@h�
�6��q8��`7��s#KK��a���A��;0E@%h��(!�]�䑺Y-�;R[��=7O7�t�^��j}r"H=5"k�c�$m�lr|i�G�����"#6*"�}�I%w�+2V..�bOaJ淹>"�\|�z��P�@����;�6FTaF��yJ`��|��cJ�ر�{�AҮ���d�_��3~�����s�}ydB�̵�^��M������/���L�,��ݍ5K��ŰG�x��XE�c�`�)���YLۏ��VxM��p�C�Z���Ua��d��̓CB����":��fDH
�@I�{s<�e�L)o��(���i\R+4���L`��(�F���2#�/��(��;b�� 8��:y8fA��3e�d;��Z�,��
C6/���\��M�^�8S��'w߶�٠h����컵)�-#��/Y�"c���V���r�%"/��q/��r�a�I�ȜBXٺWg�b� #V�`V���[�Em. ��q-BdEC�5��b?���΍��qM�I'��oח�z"�wO����8M���He{�|��5��+L��j��t��9p��uh��`ٟ�_��K��e�� �.�~�G#	(�R�W*
����)4 ��Ԧ�c�a�3x�7}�]<D��-ݨXO��a�%��C3Nf�(yD
��J������G:H�4Ek�?2�k�M�o��Q�Љyb-uV6����t���*�tѕu���$��g�0�vguj���s 4��<lA�p��!jL5���o$a���?I�{|���A
l=� *7Yٸ����*���u��}}�v�� ��N|E~mVJk-�$Z{��v8tϻ#�䮗W$��R~u�2�.�HτTb�픜��{vC�Du��=Z��2sS�wm��D�h`V�՞�ZPN���Y�d��x��ܲ�h�z��{ǲ�0N�j��T��w_*�͹� {r��RO�C��:��7�4����K�蹢�$7@�����g_���ˠ��*K		|���{eE�0��l^�����#ApVً�1��y����A���K�' ޏh�E&����o��T?Լ;SD�!`�dd�&��9���nb�]����[��=���ǆB��v�S������������GQ�׿Cd��~�����|+k�v�A+2'<7nY?B��[� |����Q�u�;mNX�.=Sq�Z�M���dۋ�o�#U�hɉ� ���3�2v2�2��oV/�!�B��h��PP[���M���Y��a�����ԣ��(������V�'6?��T�7gR'A��*��b�o��ց�d>���V|�}Y����(���=�ZgG�\$�~
Og�|mT|�R��<)� �}1�^eu���ȧ����1tak\�71��p�i����E*:�ȩv�\�@�7��|c����R�/�_i���˟[���y9�9f7��n��[�?���T�+m����ct�=7�"�͠")��6ԉ���Y���+����'�-������{�Q�K}��#�v~��uӆ^�c*cjB�L�^,=)6N����HrW� L�Z��ņ�A��*��ӝaޓuz��5K��<�9#��M��H�Rn�A����-���KK��a��Š�3���CS�8Q��$��U�.W���k� �#�Jq`�ռ!��2������sg!,��}ݟ�� ��vZ9��4p�}KV��a�G`��B[h�����[?�z+4������9w$4-�J�XN�go��al�ɉc?�^��n*��%��0�_��'�9i�P�Ɠ鞵bͥ��2�Yew}�@j5���5h�����7�.Z�`���>��
�#3���a��4�/������@��C���?�f���@	F��Y�!l���/�š��J��/�%��#�R��m�W�o%��LӋ���N��
����7Ϗ>��"��4X���ƙE �I�[�l\7���2-~���
��ѬSY���#2���=1�	t�wD/z];�R�f׸D�sũ�fH� !�#�˂�͇�!�������������`������[���~��z�ʋМ#:��z?8;����	�,�����+�Q����-VJ�+��1GhL����<��\�ȈI�:mu�]��Fi��ib�Zʺ��N�+riO�U�5r�yNw���w��	)�| rKH�z� C^���e嗮&޻d�=];@#Kbz6[�}+g�IZH�zaFJd�����P`F玡`�K��ѝ������kZZ�5�E��Kq+�ie�VQl�nl\�Tq�~?�3�ed	*t�뼻!�.�ݓCr��Hޤ[bs�)�o$�4?��D���)��p�B=C,v�hET��L��u�}1��VԴ޺8r��_�i�re|��B��C=+]��R���j�@��s�+��iXT'�4�v��T0�Dg�JM?Rk�1��)�gtզg�Cƈ��0����`_�E//��Xry�m֒�5˟�@�6�,e�.��I�\�fb:�g��<b��.��t5:��
l���d�Cs�,y�*��2��[
�)V�BV0w��-�@�;�J���G*���Sl�s?�<���iNUh~˗�N4a�h+��AM�UU�Ķi_՛��*цh~~ŭ�	����GJ�g<e�Û�L9�w�s�Up�M���P�|_"^��h.R��q�e��o�@���=U�k4[�řѮ�]R��]}Yԃ�c$k滱�1"��z?	�����P�%�h�hͼB7f�h�p58<k��2�k71�w�)�o��������nk�lbB#c�{�vo��?Nݔ�e��=�����^Lgs"qbW00^�������6�A�,nNh]C�"�Hh���>����L��;�a�5d|�'�Au."FZu����V�^�cm霯h���Og����n9<O��������x��8%^|�O~k"PSP�]ϠXF��˷��S��SH�W ��$0���s����	��\G����S/M��3iC⌨������9�6�o�Ay��R�X4��mU^����h���Afl �u��,�P���%꾼�E�:+rA2��"ƫ�,�b��+����e�k&e r#��N����z��RL����-�|�fZhm��C8|1]ၩ�F�ԾS7a#S�]������_��N~�`?�	n�"�K̯s�Sٔ�6Cf���1O�����f�]r�רG��x����'��3���J8��X;�<��3���`�V��l5��d����`��u,�/N*�|���J�,�C�[��0�\!E���TO<YW�뻿4�~mi�eP��Q�F�\���ח����;�����=j]���\u�$]��Hi�6���ٜ��\푻o*_߁�d��Y��v�'#m�Dl��d�Җ $�����AW���^��FM��E�`�����X����u�g��*��Z����.�_9�B�B�P�ڠ1��8-���
��phR�lZ�t��<��� 9MЀ��4I��b�T�k�.����`q�_�T7S���N�VX�A������N{Ϝw4B0Vd�rfm�HYN�H=��d{�7	�!b�QG%G-�p���r,4H��s���K�$��g��Q��H�ݔ�`�J�aIne�PN��������oޞ�!��ݐ�=�ODh���@.��7u+>��_�!6����T7 l۬�wp����l��I��F������~���G���UiT�#�i���v֑��#Z�A?�h�l�m��t`��-�;�^X�(����{��?�uߩ�䋴D�i�x��ȘG�Mlj_ɛ�,[s�X�L	��D�s&�������S�<	�ON8t�"8fQ��pf1��� �CJ�7�ì��Z.'��,��#�P�ڭ&"��)9�0���pv�jD��e9�-�|4�&,��\��Ez��C:�*b�V�j��5?��ki3���i(�%X��rz��,u��xT%K��~�2���:�A�ɀʕ�T� �����T�AT	ɝ��1Ut[��PY,&�����N\��F]@[�E[��[�G������=�G��l�3QӗQ{���@R�vs���q�;`��;�x�*�Ц�76�OJ
=f�k����ځ7�U���6�T�.HGh;��Ѫ�� ���E �H)���WY{��X�&|>^�Q7�+!]R�TJ�?I�/F��|��B���#�Ԉ�FX����-�k�[麟zh�����ɍ�o��A�#��2b��]��{�-9rNTM��d�x���mHBPA5M����$\����#�i�u�ͷ51���êK�dP���I�7��V��ׄ2*�5��o3�uu7�o�
��p����di�;c���<��L1���l����J�ýUX���~9�_3��#�Ti.I�=7 �hKE"�굢e�8�#�k�_y���^9ԭ���
wiw��In�%2�>�D�)69k��h�qѐ-��_�{���Ve8U�����c���Ni��E�y#��+��q��оܮm�ʧ���	����gv�"n��&1�-Hk��?m�N�5�.�8b�#jPph������By$s~���}�.�ә�xƧ�BԤ��O��`I�N����uKh_�
��ivA���"�8���Š�_ɲ5��W�"�*B.Sr�4�O��0Sύx�i����?B�^�=�.�^]'p�r���M�m���O�s;�`�w#�1L)��M@3�w�l<;�^���q��L6���"ܓ�+.b�^GP;�z) ������#;:����pU�!O�ԉo����ayTL���m�G�2 �}�m��l�H��˻a�7�_5F�P'�<-�e��'���%�>[��(2ɷ�S]1��KIr��KSQ�&,�C,�?\��y��\=�w��:�7�D�z6'�-MWy��R��p���xq��
)n9���o���P)�S��l�e�_�]�g���9x��J�g��`�S��-�vj��\����~֠�)�v���@^�1������<�*���`����l��D���SŹ���B��r��oQ)\�_��HL�YT����t@��v*��Z�`[��M��d��^�{��#�Ơ�R7��̙i�M�d�?����~���u���܏����F���d�\ړ,/�K�k����S2�/��+;G���p��YR>xC|�~���zx,����槟?��,�%��~D�q��)oj96�(�F��N�,p��ڑq�n���>��/*��D�{j^��-imq�N�5�P8�
��/��)MNoǞ�ߎX7�����Bfܲ��V+/SG�g(�]��Z��V��2�$b�K�r�)�6�O}o��M��`������B�j�NÊ"��H����m+B������[��N�'��f%϶ݛ._�D��B�`���xn4cyz�.�d��-|enr~*$y2�7�������}��z�����o�=hZs�C�+RT�����W[1�-���&�_݉*�f�L�`�"ES�+�����b��L���r�7t�uY�@=L>�0�P��6�$i���.c��5O|������?����a���La�5�	�a�|�m��߇R�!���[��\��*S50!�M?Ai���:=}%kQ ��![g��,��g�q���D1N}��#�aD�GeA+��������w(X�]x%Mݧ���uk���������÷[9�P�2���o�5]�I+�{���b�o&E�P����B��G�(W�1�7�-���T�
�+��Z�9Y$��:c�$����?&[�qߍ�X{���tCV�X��Z�v�x�0%�L��s$pI�:��:�}����G�f<�1�
("���5�|Z*�kP�&���NP|p�<��h!�G{hq�x�rʪ�[���h �8�E�zfr�W�I���R1O���	�,�$��5���^��/E�}���\���:��(I��E^53��r��$r����f����ᜟ�ʀ����C1�@�!� wO�Tj��}u�9�}�1W�G�㸝8����Q���7&{D�5����H.��٠����K���$�漒N%f]�� W���?%m g�ĐF�ŝ\�>��.ٛ�jL��;��\�l92j�u�w����eh�!}�`����X#�K:2��i���!���ψw+aH *���cLPa��[�D��(k :�A�~&�����?C�¬�äK
�j�j���1��0ݘ��.H�%��s�vƍN���/sf��J]���Q�w�=�\�2b�EF ��Ws��ڪ�\���9��>x�c�b�3��}Ps�v�K3H�R%%󆰯]yj��R}�\��`z� ",Xv4�$�w�e�} <}1ZܤD��������Ir��xR>b�Ow
8�~� ��k��*5��;��l�vMT�D��TD�Du�,U#09y�3kLl�g��s��2����$.�&B{�Ǐ%,��f	��mI;�W�3��}�gZ�c��x���,?����1��������*$t�+ċ=���݇n)���w��$N0��;�q�EP@�d��w��;ut��u���*�f�:��^�/�(�N��9�gr��ʳjFR"n�ɢm���l:%�xa�W;3e$�-��rQ��;l73�:�֮x>([Ś��;���p��g����Q��r�^��j��W�<#˰��U���UK,5W��G���Ö������+%�O/v	a����4�����yd	�3?^�܉�,�����T���a|�Ku�yÇ�QآdU�������W,N}s=�l�~�>��+$?��rp����1���6�2j��I�l�#B��F�Oz�@s�F��'"���o:��*��F.���)�>�#�%�H��e��\46Eʓ�,�n|i l\�E��� N���(Z���Mﯹ�h0�..X>�WZ�p�ɑ��t���]-��d�u�"����ųu����ߛ�?�K�>!>9܇J��[���)��Ҿ��T��`
b�£�� 0��-�{��p.����kn9�7z4`y6���~ծ��� ,a3�&S�C-�G(�-h�<T�զZڪl���A�Y�^�8,��t�)D8�ҁ���Z���e�Jo�?*���J�Ͳ�X7gwH�k��7^;t74A�E����Ķ�f�������ᢽ.N��FM{����n8��y3jtϿ�Y�,[��5�q+{^�0[� b����'J%e2�TM�]��R��n�|�hf��o��CㅸE�1�	�?�w�J+,�S�wRѨ#O������}4�0=��**���T֊��H��n,N[�^K��g�s���%ʰz�+�v� �j��O�_>rS��9E�udgh�O^�0UY*��=�����+�?e�v�Q��w�<�s"Ph*��	���BRY��hgV�Y��}`��m�6���!��}(��6��6��&��O�V���1LP!E���cX!��Gr��f�Կ"ɍyʜ���ٲ¾��ȉ!��X�9|ZI,?���]��,�b��?��q+2�Rd_7����z(>ޚ�b���ե55����9���sw�$Z_��M�*Fsp]���?N��/X��O�E�����Dlȫ��Z$2�LSu|�a�d�lK7�.��W�� |��-;D���"u����Xٚ����.O�!����6����_�l�XTQ+oFC�O�f��j�~���uS-
��R�p�0�-K���9�3G��D�+��9��?A���.sZZڶ=�-6�#Y��@��xO���uL&�`m���>V�{���%f�7�Ib!����F;��V�O����W"�U��ɦ���Ru��㿯�>��Τ�ќ�F�Q2So4��P�h�A��Gy*�u��n�y��%	#�F$!JM����|t��u)ݘ�#hq��݈S�oXmL��ٕ�$��=Y��ڠt0j.�6y�
"�q�nuf�앪q;./��#3�sB�t-��rL�V$3f��=���;w�`�+�c��:=�6�uƟa4?��:�'iH U1��9b�m7���꬙fsA{���ʌOS1�y�]O��]~��[����N�<��j^���K�q5 ����x=&i�1��Ր�u�}n�|� ��Y}/K�%������,���O�i����!�-�s6p?�%Q�=�M]�I4�[~F�nޡ�������V��Az�>q~���ǕWz� *%'-�"�c덊�l� ą_�o;�y	_�=��k��� �_N�8��J���g����wu��S��1����;}�a/��_ꑾU���Du6����ʖf"�3bD�둍�W+v���v���ﰆ$QFЖja�_~>}�B��n:��"A ��ܚ%�v�g����!�M%�z�0WrOi�:��ň|�t�38��y��K��=&r"m�x/q�-�ʑ�1�F$�'8'�'Xqs�uڛ>�U�'�%���w��%A������~ �1�+P���FH��z�j,�ل]B��ܶ����>>����ц��.aS�g�x%^�yB&�A�|i��`��Jl4�.=�m�����=o$V�K�vC�݅�v��b���"��Xf��vc�aEˆ���/"��&/u������(��4�~�
�d���o��|�NxҤR����L'����d�"�r��JD�L�8���KV�y(�P �h����.~*T,��01���O$�i��wh͝��9��s�������ٽ��C��JF`敖�A��S�J���l�T�,n1(Dv��GF����ue��X��e�,$�5t��5<�,_�8\�n�H���7m�RD���Ğ�0<E��y��m._�сr��7���0.%��%��#�T�"�Z;B�aLa���Eӎd��+|�V�v����_��v���&�U�ǩ�<-�?4aQ�,`�<Zm21�Lc�b��_���^�k���U7���O�>vi�Ș��[�c/���9ڡ�� !������d��)�1fwj�[8N�Ϛ�mmi3�"P�p~�#����G/��1P6�}�:�=�ᘮ��~�t0�0�g�Ć�X������q�{7U�����#������\UQ��I�b�r���ҙR�����^�q�3��х��a����/#�nmCbV"�>Ў�_JB����k���:� {�{�^eb�3���`,��/�����,�-P�nST�S#��7F��_���fJ��ä��@�rz�\�?���顨�ZE�!��v�uc���I�����n�^`��'��u�D��~����Qu�</-|�`_���3hP[��Ώ��P�iɄ+���V3GŃK�ę���&!h+���S�j���C���K����D�8X�OG2��%z`���p�:��.�S�Z�
tHT�4��Ǘ�������lԈY*��?�k%p
�҅�fO��}/<q��q�U︅x��K��ph}�*q�k��"�N��<�.�;6��/���Ъ���˥�����=��*��foX�c�{Yh�M�8n<�|xC�-Dԍ�Z���H���|9��E��M��Q���'�n�-�0�5���+�ھoD�.\�n7��8L�����[�� �2eTWA�[�#Sꈳ�����a��;4�R�na�ɽ��Ve��$.�85��A$'�	����Z���	l���H	3�ߜ$���{%���M���>��rAWt��J��`�$�#H��!V��n�xR(�hG$�IqՍ���H�ݍ���$6X{X����Li�L,��!dXֈ4//��o�D�M����Vh�=b��{�0}����h	;��Ӫ^&kP.��0n�)k�=O�d�e������3�Q-���D�ĳ־.6ECr�1��{13
4Շ;(�?��,���2�<5�jɘ4�v
�}!��#M��2�p�"�Q\�/��8�~d�[Es9|�'����ݶ����_�d�C���|�U^�x��̆Ә�7��?�[���F���X`���c�<u܃���� z�9?,Q��pL79a
P�|���g�����ER ٖp1�iiॠ8fBc�}�~H7�D�/#��;�Z��(աCm�S�&��*-�抟�7�y����ז�r�J�,R���X���u��l�t�a���)s$���F��=u��O��d���<f"�h����̨՚���7��j<�
�T�h�8��9�Q�:�|#h�}��/b+;I�.~]T���d��fF̿��G�(��
�j��)�@;�ҷ~�K�_oZ�N*�����|�s�S��k���0ls�%���Y`��_���t��W�"��9^��R�
r�	� �{�o�r\3 ���s]��ҧ�D<�A�oi&q�42e�\1���JV#+Yx���(����?6w�,&�hxyR�Q�Ԡ
pʌ+p�T����[wQ=��P�h��M5%:BB?��ڡK{P4]�
����ql5Q_5ǩBPp�O�d�L.IqZ��� �U��o|��|ƭR���*��t�/plUĄ}��A�&��!�Ncк��OZ�)�z��qg8;N�mX޻�+2����Q�t���i��>��?�'.,4Ӫ�!z�x�)@�#q��r�p֧f��_�����A�)�/�����Z�[����a�A,�HM)�D���ތ�1Ks!��4�j��<w��kO��@����Y�ȳ��=r#��a� �G��W@��%�X��R��snڦ�7�+sj�q����1�W��8�ڌ'�<��j�I��mai҅��ae���e�p1��)xY���}jѵ�B4j�o #4�K��6�6�B��ՠP����@x�jD�X��Z�k�Xk5Y�W���΋�Z�*���5XU%���J�(��UIҺ����69�@��1�����m0ZV�h+��&��zGA��,OԷvK̤:v��������jfg�_�4�w�Ƈ�R ����7�6�7} R��$1�ڒ+�-�Ҁ���m�S��������O������$E���&(~�'Vf���	)3��e8��
�C�d"
Mfi��Nx���U\ˌ��.P����r@U�/��	��`�L\��M���]�$q�楚�MI�q]Q+�[8�}ҩF�*Qh{�U�F3CPߒ �MQ��}��Dz�6R?�:��K�.L&
�<�.���w�Z$9�o�ȁ%E#8�����#Z�U6�CԊ���v�L���J��j&]M@��@U�� D�Lߦ�$��;�h(x��ε��?:�{C�=a����	����L5Nt�B2�m���@Dy�����b�M}�uρsa�]������B[��v��Z����e��J��ұ�2���e�Fx(��X�P"G�����3�t�3��4�1E�hߺ� �����:l`T]lH����H���:�i�ԧw�&Ȱ�`
��(��K�d3�;����Eh�}~���S�\|��4,�!��DU�	��y�|��E��.l�q}�6{mM�"����?) ��'���V�6�o�(�Pݶ��x0�ۘ73�� +n��D��tZ��4���隟���?��M9�u^́����_��
|_1/��*k�,���NB������$nE�a�)BMæ{
��$W'�u�n&9�mE�)͛ �Ȥ�6l)?�^�u���;e���e,,]�/=|Y�q-]S[YR�����k�gh�y�� ?��U�!ҭl���#w�I;���I@y}��9u3���h���"R3y3c?��8�&}T3ulDXz����[��c"DR����@_�i-����XP�F,�8x�?UCb�q+�ZJp{���H�7�n`Q�M��ge^V�LG��x�!{󪜣.����I%�A��9�f��ֿͳyAh��%x�*0���ƌ���	e��L��ww�P�%X��܄���Nя�%T�s�t��e���b.�\�ܖ. �O8B�ǁ���6�W��A���@�P�A�7�E��i=�ri����v/���郲��p�z��&(Yڣ]�mZ��"&���Ր`�q��~�@�/���[�3�����Td��x	-B#��&p�
��Zԃ��͢�c�����GM��4g�=4س����H�7(k�/�[�i�� C�n��R���0@�P]���-�����P��*@H�
妑�i��$0�V��KcO�N�:�	�s���G���$��78q�B�r��Yq`�&�3o�5>@�},1ޕ��3`����Z�;���/�*.kaƜ.�)?���aƖGH��r���,(���Z�m�����0�HT��-ۑ1|W�BHe���l�����;5b!􁈽h������:.Du���?�/[���i^������K͵r����wEZ/A���(C��2�ղtS�NCO�%xزbb�uT�NAO�o��U�ϥ�-�	�^Y�:t/l����s�'1��UL����7�y����+����K2ؾb$+v�K9�[��ݳ�w����V�xlx$�V������'�A�v�'D ���0t �}A��oF�m}�YH������NA���AMK�<r��r�>ܽ4`�U �J�L�@��fb:/"�[l�&�/W.Tˬ�t�lC�~��فf���l?z�a�P%ym�u��O�!���bSt �R�RئS,��xV|�o�*t�>�JK�2����C�%��6���y nI'�Qf�݈��z�6s?�cy�������2kR�0U�	n�Esu|B�����r�ܳ��4w�I)�7�ԭ`49�b�,C��.6W����6�f���}Rn�,� ��>m$�K����(
S���ޝ�(("Ѵ���r���@���{L���a�$~���7�q�93)���W]��Z.�1_�"r�Jow�܊�b0�<�ǅ�bw�Jr�(q�1Q��P��(���fb�R��-��2�͈Y�r_n���zmzE�2��B�h�ʅ��+�&f<W
,�F*��T���l8����b�c����-9M�|lR����Z������5,ّp�#�+yR�b��e�A�����މ��0����2Z��ef<�<��<�/+~{n�s�G��s�g���8'yg��,�5	R#���ntc�D8�����&�:0cϐ�ߟ�/������Y'f��W5�5�,�x/9u��u���ￎ�G z%,A]K��U�K3�QW$��U �wM�&3�.��모�/Kd�[���ɴ�@D��wtiEq�l�|�A�������Y<�O�*��B:a��<|J�^���Me�5��UH��q�"V9��<s~/�^�������GT����㍴Am_$�6���3ofu�:�o�Z��9�Q_ �K�^<�2nï�EtnIL�6�j7���xz�Z�e׸��=�J�z��#F�� ���;��&k��}�!�I�jD&�29z�^?����5���:w��ɝS��Y*�<�	>��m�&���P��$�L���}�[%~r��C�r�)�̐{{_�X� Z$1��4:<?�Nht�@A���]E�,wm��\E�����τ�Ԫ+��O��X��?����dD`gɞe)��h]0j�}�Sa��ĸ_�d��NK";�=L�]O!-Z����xr����jx]x����X�[��uF�4����D0�T�j]�'ޱ�L�R̅2 �T��1YK�H�����~�h˴�w>a<q����洫-��r�-�q���Pca�(TȓL���#)NګLbǭ`�8��vh�]JYê���tXPG<�w;|�-�u�	?���0[����i�r�j��X��[��&{"�yg@�,%_�pH��̬M z�7�2��/�1+�
�e�}�TK������ �%s�Ȝ�v���� �5#��AOn\�j��o>�1���
<
��1�1�l@�#$+�^�5��R3(�m����>�o���ۮE׉L�mo�����ǹ\�f
�.!ݣ�@Oz9� ���8�<cy���v��z�o�^d]rC��Ј���Dq�U��gX�Uv3;���8��ƺmjf��1��^>��A'݅5X���&��8���4�uD���ͼD�}s�s
�8���5_�����@��}�	��^n�n�6��n�4�*�Jh#�RʜbA��^2��
���E�r0�)6R�d �l���WQ]S�阎��px�Utx�gN�G��W�y�����0��&�_��B:�^6���z%����w��鍒�?^4+��0$��SҺ�����Q�������'Èʳ!�Ql��A#��*A����O���|��Ss��VB�� Tvu���y��/�V�S3�էAy{� �W�)����l�9C�'���[�Dhu�Y�S�K%E��|!� j;l$n2"%Ӡ[&6�_�:y��QI��ʏK}3��s�n��$|���[��j�H!�F��|����3#m:�n��;{A��QW�+�?(��uH��Sp��V��>g��p��s	�ڑ{�T�7�u��@���%/�/�Ed�����SY:�����֚�,D�2c�U)������`�(Z���� �fƫM�v� n��,^��o�,˅�YjzMPt0w�'��ȍ[�c��(��
��7T\��̑�i�X)�3ɡ{,5_|q��Q���?�&����>�,J�CSWU����������x5*F�ur��7Q�N��7q�L���S%BM��g������V9�Z1`�"7e�ɼ�bj�5('vl�n�\�U�R8�L�v:m��四�g����������^�h�j{���QQ�%J�ݺ��hu������FY�U�uW�Z1
�����͚*?���2ٌ5L^@��~��Hy@Hǖ�BWkT@�v�/2W\�}�_@�������ߜ
0����d�Hɔ�w�A�G�h�`�g�z�G���C������#mɹ�>�n��TH4�I����Y�ED=��kjd(�7S[��:_4k%�N�sQ�Q�Ԋ�;s�{p0��Xn����Wj*����<{'4�{3=��x��Y�X��Ǩc]�/��
uS�#I3����~R���۩Y��:�Wk�=~�y4T~�JՓ���x�15	�{|V�5�^�H� ��r�j�e�1݁�#fe�؇C�m$�_���1F�����A���p|F��O��PF�z���Ux�߅�?��	P�	���2/������TM0��ƽ ���; =x:�쳆خM^���\�Z~|�oj�0FfNc�KK�7�V�ߠ�C���ȇ����#�i�l�$�$�}��ՙj�X?헲üc ��lA�#UV�=�����g����,E��<��/c���sOg�8۞���w�$a���9I}��Q����xu`"����k1���(=�H�����N�E�� +s��*��%����iUm ���fA]�����ȶ�ԶUMG+!w�d��$e��YUt���2�u��M���*$���ӣ��/��g��<6
�h���2,���#�*!aH��(��C�����>{�̔r(��2m!�m�t��a�g���lI�"$��[�E{*�?���链G��-�<	�)w���I��/+'��R�+���������w����š�<Ru(S����Ue�:�A�?�z����^�ab8�d>+f�.Hķ���'舶�I8�Z�bb3"S���z��W�R<7I��A,��hD�wZ��Ւ%B��v�s����w%���삅U�>�N>�@�b�#���Q�V���?ӻ�_���ir���i�����`o#|:q@�`�ן�4q��Ő/�������b�{��MÖ�� prJ�q��Z�������&�'���\4�X��y��t��r��D{Uī1w�G���S��v�8�8ӢE�XW�dx|6� ���}�>)`�	���40<H���9��qX�A���}�2��?�(��#�����|���Q��9�4"m%Y�^�oDl�����b]m�J����h����u���(�qV��֡5!T��P��S���_Oh��DTq��������\��M쫧�։��w������?��ky)�;n�:G��8�`��4�?xTѣBM͢��U��z������!w���K�@�V<`����3��~Ub�o�VL3-Un�1�]�LF��Yn���x��?`���~��
\1��!A�UB�ڑ��X#�p����j�O�,���'�&x�9\dB��Tj���\�_J7��Eߎi�4Z�Jt�F^2Kn>�6�Ya�no=�]�D��Tw���2�8�Ә�Ч�jj�J@�C#z)X���9ro��˒Ϥ�����UZ���v�F�3r��j>�RŐ���m��`�Z|��yȉ��pq��Zٿ����m7S���l�|\�����T�>X�w���.1����W�V�`����LPYn�� w���2*�#���H���f�� ����-�m�½�52��ӭ&�g�\8|�9���`p��[��5G�Zv�����&��cE�����RA�x	f?#�;��j�lC_E���k.1��ؑ�5k��+�����D4R'H0^�ԁ�L:2\=7}��-*YBw�^2\�w�=��@5ͰI�L��WM��Úu*��Ԭ�nR�n-L!�&�uD�Y&(�����R����y.����(L����?@���1L�\�]�����?�^�}<�R��� �ً�����m�Pz�il^�A��.��:UXS=C��Z� �M����(o��mſ�K�f��I��b2TFm����:�m�񯖱��t���W��;j����1���%�X�)
����<����`	��[]�3���@f��rL,o%��R:O�MБ�����E��.�.M��%��G��s�N�`L�����!�F�p15] �)�j�IT0��j*]W���������H6\o��`ܸ��a�-� Ur`�@��F�
��̒z7k�qp�u�0���r�t�%�����y{9�bE��	퓈TH`�����.��ed�e*]��}����Y�m�$�h#i��MS��M��!��q��:�p��i��8@���Ϸ��^�W{)OGf���Z �%��*o��g��˰��9�}��FS���~'�a� R�ni��E7���t�p�X�L�����4o��؝��J�d�ԡ*|����٪f�ϻ���|Iӱ{���Gz =�g=�]�	�Z�e���H�Z���Kmq�E�(W�@�E��OG��EA�Q��Y!�:u���4\����P��ca	m��{��g_�i����f���0�C;K�{�
{��܃�Y�fUu�r�:�/�,��F{]+\���^��	n��N�������k�)���l���0��z�F���²�� 
�w�Z���J6`�&��u܊����-�LA������xn}I�N�<1���i,�Z;����g������8I��'k�׿z[��E�}C�Ԇ>��Y�G ��9&�I�t
�=e$/^o�y�.��4r�G�/��%4m�`��4Q��t��������s#�(�`�
f�7�x�c��:�,�K��6��j@���N�����Ag���}�M=�E��u����A��p��ٖ�@�v#�:mS�*������j�j����N\��j�AܖO���ChLd��}��]Q}ȒH�a�~i$t��_��4�F��t�����#"�+<WC�D��C�$�	'�0T��t��yzEoڵY�qb­��¡��	k�ϳ�y't[�\��8���dl�9fF��s펐֣W�p����4U)ByZݺ��X�� Ay!�lm�Z� ;��v�����k_�H-Y�)��װF��a��!�z/4	|��z �ѡ�`����Ҙ��������r�\R뒮��s%֒��t�%�v�ngd�@X�ٍx�L�6���0�N��w��1�k)�Q03��RU}��N�� ��H����7�:�`LB�n����b���۞5,�-�s0�\k���	�}���/0Ц��=��RRPL�ro�<Y,;s��!���A:��ԤL4��c��w�	�O�'�|�����3C̱���S��3��}W�2�ݵჭ�Ң �U�LU����if�_Zh_c�Nw�������OJ��s6<����;���,��x�1��/4�������U�E�:/�����!�)���&����<b�	w ��#	h��H{�r=𜑜�捄����=��@����uÖ�&)]T3�d�}��FH]|X� ��B�]�V�|�y~�e����o^�K�!כkA�,oT+VG]ȃ!����n_h��n�!_"�AN�kQհy�q8�>���ǔ"4&�V7Pn�kEm��Iƴ�Xrq��Ϝ����������`=l����*�|����"f	�~qi~L =����k�Q� _�ji�R������OZ^2�L���D��{��4�F�Fe�'r[�~�����@1;���"�?X$Q�|�����2�
�Qzǝ�&9��-M M:�*�üո2��H�Z�]\�p5;�k
��c?� ���M����8�bgI�� �sh����a��X^ �	)��6	�2�2|�oFƬ��'Qb���y�\H_-����|ϵo��ؙMTk܇�ו� �TFO64ۄhր��dj��X��z�5����l�wB�@���<����� p��fPT�]c\շ�OA���{d{�_�ro6؁�벝c����j� �/㳂B��;�wq�dC���֚����裸�䁊Tzs�;<�hAPk����3@�0|p_EU�B�h<��Ń�/�����S�"!`�� ���G�p���eBg��3�]������S)�:�%�*�{x�6-��m^�(���0}c+�468Q�V�^o-�f���'��%�e9��1!�n��V0%�{̬ڍ��-0R�"�s�x:��E#�.;e��`�D>�!���`�;5�K!�[���W��ߐ���g���):�â�o�D�.'@??�����+WHB��?�7�,��sݣ QZ�H�t7,�b?7}�����;Y����ڍ�5�>%~]�b8霶D�p� ��Z0��ElK� W�����$��L���>+3/o(Ĺ\���~f��Z��~QV�*#|�ٰ�eS�\;B��ǉh�mW�.�00m&��?/@ RF���_y�I�[��YokW,�p�*̩�&���z9-P|<�8�j��[���g��@��_���F8�Srvd8۲X�2��6�T�?Jxړ��i��4�c�t���ξMFu�z ~h�N
��&u?J�%h݆d�I��,W6�w&��C�(�k�Ϯ�"n�����-����6��o�Ç�o���E��f�=�@�̄B�xv�N
�l�	̰�~�I����)-f��77�b�`�g��q��.�"��Y��EJ�D����
���4�o`^e5�F��w;�mqLW+���&��jVu�����Y�Au�����A�(8�+��ҭ�DzG[J��C��B����jp�L�A*��E�� �׃�Ǔk���Z&���
cL�oߦy�ūe��0x9�gOsӏ�0��H1,�["#�0Q�Ŋ�D�(;�s���+q����s��t���y~'���&t �Fĥ&����_�H񲵳���D����^�G󯷗��_*؊B��N-��k�چJ?�&k��	���5��UN�����r'!�"�1��pc�5��ԛ3�G2x_F�kx���䲓�����΄�Q��n:��ƄJ5fa�l��Mg��2����B��\We�]Aa�
��n��˚v7�s��{�NϸO?��lBD���um�U��Go����B�]75Ԝq�?�^w��"�ۧ��9&��+�^�7�!y�%;��j����'p��	�U�>QP#J;��o�y3x��B�ߚ���b��t����=���W"�Z��F���%%A���%-]�X!/�r��O,�,���a��hM���;�Ҟ5ct�MT�ٷ��2�pc���n���Āa����T�����{��M�+�0���4o�0�&��Tw����p8@�sj�~ ��wP�[��[�8����v�F,�RA��i
��������5����\���r/%��%K�$�ln��NK�C��SE�Z�f�M�.��"�*�2ln�11�8&�H�e�1��R�6t�Y�-Z9���Gg�{
r��w6ٹ��=3��,�H8�%���<t�86)��&���%:�SE��� -"dڮ\���@�'K�QZl�pa�E����P��XR��'\�q�s�}���rK�Ep� �A���0�l�X��F�����!���VΚ�~[ful��P�*�8������'HgBJ��4�Qis���:j�:K{�x(8t�{����x:�eO���r����9�8��I`"?��^�������d?;�/��<֣�@'h\C�>�2��'b�ʔ��R���:2D���c�mQ`/@�&=�j�����t������FJ�ZQT��5D�|+&�nz��gX�	2O�[�3Q��j�h���'l�4oH-�e��I�q�h���{��!g��~�&�/_���n��׹;�Z�Kٰ:������'��ue!���7^�k‟�y�ᚄNIN��w���tF�ep$��V��*�U�CbG��T#��� �&���AY�,��&Ԭ�Q7Տ�a���e����k�TѦG5A���5�N\b J�aTQ@aF/#]��������V����'%ǳ���A��4�
M&�c@�lQA���<� m��]�{ǧEߧ[�4x�_�F��w]	,I
Y��}N�w��5��@<���[1Fy���t��~!�u�h-|=|�2�^��Iu�Q�Z�zaH�F �ĥeF��;L���]B�Z��gs�d�x;� Q�@�C�X�k��l�G�uc�K��<e5�G�́��li���.T��G������L��q컣��j�;��F�X���*4�PE+ڌw�yH} Ŗ5�6l\,�M*p�F�-���/�
������z��"8Hz���x��W���Мh`���+�@%��r���)_J#��r,�$W���ߔ�����Jd�Ҽ�c��Q:$^>zihHM�Lz���y�sE�[el��>��]�f&��dpd�M�>-�"wdl0����n�ɬݓ^����Z!x�YT��gX�^�����N��T�m!>=(�q���%�G�D���or���f�G"��à�`H�������:+`��78k�[h�^�MC>S������I��������\U C�T�"�##a�D����>�Ϧ7���51&��pB�	��U#)6���"�oΤ��TC�2��"��WR��!(��!�تAm�}�m�C���AT?N�,yo\��Y�&R���霒G�JqZ7���ǳvD���B�ԍ'@ޗA��s�v��Yw�}�z�Ա��ʱ7f��T�u��!V�Y0��4+���
uWCN�c]�O�Ъİ�+C�@Һ(�D4/���;��9�Zt>K�g��c������H�ƾ�a�Ws���2��=���\%j�6 p�[MeR��q��	���^p�,�ƣp��+J���P�&�mW�$�g�r'��Gv�m]A#*��zA;�vs<�dP@+,��>.�(�t�X����]u�+(�B=pr!+�/f�]�<zֳ�k� ��J��,U���L����q�w��j�J�x�R,*��xr���=p�Pf84MR��`��HZ�¶0�&�y'p_HG��A�����+Z0�-fs��,�ן�+�=�⻪���Mgcxru]͋� +m-�)�M�������MʀԖצI��kZ&l�O9��`�P��N��	�	�)�љ$�F��5JՂ2�tU�.�A��W��U��i����憓����!�5�)7u�`��p[�E��9+�3x�D`�������B}g�c3Y���.vX\p��Bw�X��-k���=�J�>��^��1*�ܭ���D�%&o�,�M�l+�UɌ�q��,  vJ\��;� �SΩ�M�G�]^���>y��N������-�)���Ta�Q������+=�{2�Lչ���V�G��j3ݟ�)�b��g,�6#^X��?@ "��3�*��VV��u���S(�U�����Gԑ|� 6����d����C��iϞ��[��{>q��ica��O�<��%��� ����#���wڞA����K�k�������=!��A�Of%�u/�_;�m�������/xD	}�@B�'R?AV~�P6�Ke����^nR��Mo ���6�;ı�te�iwT)���k� ���e;���\*,_ޓKo �$��-~'��e�iĪұ�wYw��9�~I���?"�� �E�S�?���̈�e͔ sd2Pv��a)٧pV��+�4ݚ�+��~�駂�hc� �8��E0��E֩�� d�i�����8�w���4�߭{�V��`�v!�W��7�
��p=��1f��.�
 �.��{  _�`��	�Em�V�lK^�f̃�����3���zL,�[�;��gg�뱝����9��:<zP�����gN�JHy��G�:�}񄍝^�RpzhOT�d�v�bu���dJ.�q;{�Я�TI�]����L�\%3��K���Ϻ7؄=���b	D=�{��ch�m���6�4���K9}_'��V�'	�4c�h%��|L*����n��$�Y3�g���H�q�dĆ8X��YQah�ޝY��ӝ_QM0�e,-����QiPY���Θ��Ie���h+�,/*��r�Z+�`�߰�kΞF5D�����7�A�����5��ŋb?7�3�^���`eGO.Q�8 wu���q�iz˂bř�pt�p���R��˿��k42k����+�a��ċ�h���NY拁7���Uj�q�[��`qm��C��)��ŵoL����8�w�z.���t�D~̦`J�O��ĹN�G������G�Ȅ̐DRf	M�>T���5-�c!:|P'ɵ_����Ԛ���5�6I�u�MR� ��^k���H��S|:��N�	֍�2�3�c�G_�D�|�[A!����������X�yI�n�/���ڢj�R4��`+��.&#'غ%�S�C��b��k�8F��r	�U�I�w��Q�=�%�
5�Τ�t�����S"�bmq�W#ٜ�b���M
���%�6]hZJm�6�������s	a`C �����}�����sI%c��"�wB�L�o�T�!P�9ͱL`��v��IW�����<���/�Z����),���qFwn�71C}͌7��}�#ىn��Y�E�O�\���k�B��G���V����S�zF�6ae��q�����'��IN0�ns���D|4z��j���S`�󞼯��>�eW?��5'���(�ϣ�Y�b��'�sR���kK݆h�������O�U�2��rS�c�v���u�*��3��S�W�w��ۺ��
�0�,�N�ПH�O���������vI0�!#�b@��x���|�;mN����^�~���?��`�TG�	�o�Q��?�r0٧Lz�D(�0��ؠ�ׂ؎�)�/�_c��Z�pd���܋@��:<�@�?1��#
t��a8�V���D��\��&��Va�p�ꑑ�K�[[�ϠRa���J78]4tu��+����'7D7��7����V����J��*sKi�y�郆Ja1MT�������6������+����h���q�i��i'��Ty��Lݳ�m�3�rW���(��4�F3_�Ö@������	��x�Ӧv��0��,�a��ݡ���~��a� ��E將�@�2Fds
���r�j|"r2�İ�~r� R���&.mx�/8�@Ql��y���H=���s�hdw�B6㡓p+�Y��1�+��I}jY�7�U���@�̍�&�Z1wP:��~)}0M<8��0vw���j�#�cx���g�>�[9�UߔmK�=H�U?8�a��t�t���|�0
��Z~y���;
�+�r�o��Tp1UH�^[_���2���z%�	�L������w]7�<��-��n5A�Rm�
ɟ'�6�>J+���e����9E��Oy�X��1(\���`8	<�z���gP%p�&��,����0RZ0�.Iڊ:vx��j�(Y�Dп�asFf�&�*�r�<���
7Ͱȕ������XEQE��,֘0�Y��aV�,�<Pd����O �a�x���+�c���i�c�A.\�O�hghє��^-3�h�m�����yG����K���Q��;���	�f7�$�W�H鬙d_�ExV���O�O�Y�����V�5��8��I(��d�߹����t����(�#d"4<��|�Z4�GW�'1�E+�e�av�/�T!��h
���BsS��̌4�
�B�S ��k�Ik�3��4�P�L�ȊтS_%���3�>�i_]Z���j�X1b���A�oN������.��%(`Fx\@�W���N:ι��e��~�� :&��2��0������L�����Ѝ�;�%f>F@�ùE���[�Y�,�&���=�q� l���L�{����L�q��Ʃ�	װ@��,>Ϫ��Ƭ{e~�A���M����<0��X[�AD^N��A���iDB/3��&�%�GPO_�ly�%::�*+g	V��Ԟ�ͥ��$̅8��4���Tz������؛�f�������Rz1�G,���c�g����4zc�Ʀ@ ��{���"��M U�mH�� �N�w��#�͝��8<>t�K2�i�Q�6�EQ���K�{<z|�k�Ҳv�e'���$��,Wŗ���r��Z�7�{��C�-�Uj��;4ě��e��K��8�=$��G<J�6;̢w�}�7R;Tt_����N�Ǔ���݈Z5SO�Oe�m��ƒ�;��aD��� �����Kq�-n�ϣk�K�~��D���b����
�
�ɼU�J
nh�Y�՘�@�.Wp��W}�]��v�c.M{����bA��/m�+���m��,9�з=Wu�0'�<����X%�@�T�%���&m��tڠ���۟P��b=���V�2���X2_c;���!��P.[�-sNI�š`�9���ੜ�J�j�#i���1d'���s����'��I'���JMݺiU��,��������bZRK
�r�r��ztM�]3�654�_|6�\�@N΅��O�J��9�zUQ���YU�B˿�yGE/����>`�xKdR��`P����x�<��I�K��6H@@��ǁ �,C�{�!��R��.�đ7Q9��0��k���սTZt���Nх��)�&Kv���*������9,�[2��캼��W�;őxe�'��4k�E���QM�,���G���Ṑo��G�{�?�`7��$�oz\ǣ�!k�)�@e(�(b�Ӣ(.��D�П���E!����E��~?���^<�Z=Xɉ�ˉv.S#Cqc��-c�1a�����5�x�.��́�a�t/ɂE������������c?���^�4����C�c������D.�2��l�z� ҝ����A��LQ�@H�|�!���qc7[�)�B*_��?z��{Nϥ3�L�̝.��=��J��bK���kI�#L���2k��L �����&L����� �9�;���Q"�g�7��4I�
#D�DI�*��Y�j�\�q����������� ���h+�B�̭�Vh�~�.�P�I}�ý�Q����罈e _Zg�[1jw_�I �&��##�O����H=*�ҷ��X �����e�?>u��uՋ���0��L	^8���H]�P��t��bҟ�ov��_�O욦a��@�D�����(I�n\^]3�屰L[�48�s��t���������I�}t��������\/S~���"-t?�����߱5�/�LI�%:� �F��#����9�!���5����D���?:;�6s�Ah�pC
�|ɘk�uI�L˱�J2k#jKo���� Ђ�fz�����'��g�a�Tuł;����a��z��2=q��_m�a���iN�f�pn�E&�B���+r�d�pO����t-/�3�>���!2v����xW�Gܘ�/2�+-��S�<�/��cM�y��O�*���]����v��MЁ*)�[�r����*g�0���K�M�#�l>�dvQ������H� <\A�c� ��p�c?T����Y� �=�\Ȕ#�1��F$L{������1h�*��_5i/�В�8��g@Lb���EEY,�ӝ��<B���P�?�(��ڹ2����U�����R�1 �����,��7�I{��E�� ��.�O�bL��ے)D[��L�p��~�៻9���u���7PvXݱ�]�l���7y�&���E�b�
�)Dy:L�o�|I�D�:5InD����6�G> 8���ߋ�>�u�&0�]��ȚAP����s3h*NE�.*�OS]��`��9�Ex� {?Yb�Fq���qN�D+Eh3.c��TN�w�0���e��>�X?�؀����4�'` ����aQЁ:E�&݀�k�a�1#����?AB��h�té��P�7\Fv��:j;��s��6 <
�����C�ZA3��b�SE�ɞ8S�ߩ�[�V�����U��U�:�H�\fuQųݙ�E<�]��<���v���&*�#&�1���"D�|�
d�7\�~sHm��o��7L�1Is!�PW^��������٠6�|WA �bR��t|>[%�N�c�Nҳ���)�g����Q*��k2d���5v��?(����Ɍa�G�o�h�D��ޒ.˸m�G"�@�j��y�;ѿ����Y4�����n��y�M�)��-vݘ#����a�+����KF��4��3t|=
�͕!��`��p�h}��m���j��̄@�gˑ�n���^�qv�e��*g�M�K�!3��?A6�(�)&�X�T�tG[��KB�({j�@5���8a֙��"��	�^7=����-=����0�=�g����R ָC�>����M����3�r���96�8����t�+D��^��@��80p��SQ��DĲ���?���%p�+��uU~l�k��G�2��x��Ӫ��i��;�`��o�&d�I�H )����i�,�aP�9���6�B�ek*d��w(s�/r�wrTBǔ/�MC�ɡ'G��������~�^$��j��j�б%`=3H:x��5�6)�-�m�~�c.ŵ�jF��Y�:7��ܻ@�KđT�l ��+��"'{>�7㳑7͟�'��J]��'ʼr����YA~"xM��k�M_��y>�|�(������4���>wS9X��k��Ҁ�*��X�5�xA�� ]sGq9(�Nq�e�UlB��z��l&X��q�y���u�DQs<�ב�5�[�9��f�H�򰧛����Es��G�!J����>��^ �M,v�B5�4����7�%ސ�@�r�;�u 'i�S��>�����r4y�j� ���o��.��n��޴���<��cE��]�����%�桩�F&ri����t%�K:���8�� 3��E�fR���Q�;=9��z<s�l��p@x��� >����¬AN�J.�l��7B�6�R�K�8K
f,-�h)9K�=�Q�6��*1cV��if�@}�+5�;��H�/P�r1��av1�E��#C��z� XgT���.�Ǔ���.o4����I���bU~�7�n{�U�Z��Z��&v��ϱ�I�g�N��"b��nT��l�¢	������l�Ob�G��T��>\>T{�+�"t(�������W�k�Yo2�[u�.�o�����7!O��A�����l� #"Q���ٻD��#����M������8��X��R�u�����*��Fpҫt|�h��4�~��Ӗ�'�� _r�Lu�r�'R��I>c�ݏ�a�pK׹�1�͕S���/~#��	gy��d�5h�1U�ੴ
�77D��P�7���އ��u0�! �{#˹H#�e�����8��
`�Y0�7GC�4����y�6��}-���`=��/��5TB	�_�YVy�Uü�]%�y�{��k�9�����e�e�Qb�"_���m��9��W��
�Ί���@o� ��`�Z3���	�0���S�~��UpW7��wO��&{���Fp\�h%�׫���&��JE�a�ω�q}�VCY�)�FQ��,�&3%�-�
��[���{4	k"�E���b�*�^�DhXv,|�����h���
�Z �OA+v�6��EhO>�p��c���2�M�<2)T��B��bC�'�U2�f��IY_�1?�'^&W����;�+g�'n�ӏU�;s&;L~�������3����'�hdj���P�����������Z�w�Sժ�{�f���+���җ���b��2�a��J�"�Ud�&�G*�y�C-�aÚ��~G��!�0�dG��Mu/Ċ��A�L�&I��P��Rp����!�Uʚ�d]G��jM�6�J��/��L����.��!���/�iA1P\�h�P|���2��DG���U���e<��%͂�f���o��(�J���풚����+o�� ��i:ZU�I��|���_<��b�S�s:H�Z?% /�L�@uS�@r99�W� ����ytݻ�quT1�J�ɼ�2a+'u8b\�b	$h��d ��ߨ���L��Bw@����;�H�-�����O~L��-�5�U!Is)�a�i��~���47DK�}`�����rt�a�0�s����$L�G9����8�^���,9�[��ze� ���oH{Tg/}˯A��TE��Cr����=Di���+]���ǩ�+����6ׯ!�7]�Q'���� ������n~K�"��(c)��'�����l(-_yΠD��ɺ�>��x��k�Sx�[�����,B,����Q�Q�J-��.�{�繲!�"��cg�v{��D�D��NU�ڻ�w
�ײz(����!��D/#�.���/;�A֟/	$��t�kw�܁���JD��R/6%-V�;��-ci6�("����G��S�quJ >�x�{a]�*��Ը��la��Pf���oB���>�[Z\��c*��9�(h|a)�v\�?�k|̌�9Un%������c�U�mQ�EUf����fm�P���:������7�9p�z94:|��E ������$���������})T�N���/@����d��IX���9p��E��VH����r_"�0�M�~���c8�����S"�:� G���7?u,�Pz�ixr�l�8W������V����UɄ�m�k*Ґ�j0�|nɔ\���_�ZPf0L����L��.!�l$8I�A�����p*z-�hI�Mv�����B>�3�g���2�ų�����q��1�a��C�g��b���,L��WT\xBp��X\+��ɼW�f���r��bO��/������a�C�D�i��a�B����z�,�g	r�?�.��"!�I
S�V4,��-���bN�_��>G�p���z�r�fq����)^,U��_�4f���z�˛��&4<�.Z�"�-A^����m��ڷ�␘��}�p�v�f�Y0sҥ�jr-b]�F��u�3u�5�c����q�?M��Ul͂����x�E�Z���1�q�mADTD�,D����k��G4��}��J}3����!�^T�#rud~c
�&[qؒA�(ү���(�k� �~�24(�{~O;(j���I��K�K�$nC�%X;��[_���7cA�=]�s�x��E�s[����n�����#��ކ�� ��Y�j�	��db��:YH᧵��!9�z�m��[�Ŭ�%0�����g�7!�e^Ɠ�UA�*��V�/���M�����@�ax{��W��D�.��@[����)��'��R/�v�:T�<���.�'�T���S�������:'Q��/�Ch8�P�ǯO�<�`�|����u�q��z]�!�1�l��F774���Qb) ܛ�����=#���f��j!��mٓ�YjLj������[��{��qGQ��*�s��<�!~:i_v�I;S�����M�7-�T���j��Hľ\F��,�C$�I
���N$F(W�r�[�ږ�O��`�R�L.2LɄ	V�J�q�;��HJ�MU�%�o�Ba7s��iLms�^C�I���dO�h�2��=��}p���㓙J�F�h���K�,z�m�lÚ�+s!N�P�k�D���儵�N��
���L��l���Q-��N������	�W .�)��U]'p�K�R{Un���s4�/�V����[�-%� d|�� �x	O��PiFߣ�ds����(��J!��'и܇�h��>��Bk3�/�j����GI��QKD�[����o�C�E#���w�X�B!�� Џ��'F�O�a��,��,.y�(���M��c,���uT>Y��'#5Hq~��x$ҟf�Bz������dN S�`������ӀdAcTx���6��۪Ith츳d�r����W�U�fD��v�F0p2�?��(AO���R�Q�R B[kS2�Q�&�j&��P~�㥿��w�6�`�"�o�	=�w(�E�t�D�#�T�� ּ�%@����TH���bk��߈�P�3d_�㔅:A{�|sa4a�I.r�)�)��"�pJg�_:�� o�f���{����#�t��Ѳ��FJO]NڊHz���Zh7-F�-��?.)����Ԁ��&�C&s.�^���5CU�S(�L�J����ǉm�Ls�$�����z�/H�Z�?x��<\�Z�OZ�Z��~)x1f� �sl���̎<�i0��F�������߅{�C]��z~`<�s:�	�JO�e8��:^�B���&��,ՄZ3�������h�{f��K�1��x�����1��	ō� r�'S<��V�k�iN����8/8���X��� ȅo= =�JT��เ\����'B���$n;qh$���2kV:e�~2�q��>iQ&�W�m#�js��0��B�m�.�F�Rha�"w�g,�=�_6[�ʗ���ya�	_�������5םԔr�}�MAAg��O�߈��y���T�y���%���m!��>�c�r�_�\
���(^0��JlY�7��P}��?�	x�;�l�C����91!�?��C���:CK�L{���T�$�TX9J;�l��K�9�
��x�Z�+ӄڑ9�鐪�����]��`���tH ]Z)�:U�.a;�Z���8S��e�����/qv��kP��?ZGä達���/�����a_��x�N���8��,���$�S���-�x�d����J0�ĦMD���خqm;���-/>	2ݗC�3q�)��(96�˹��2#9��:7��R�Ç�#����Z9�x ૊����x�i��v]~����~{�v�<d͉r�}����Ǖ�tcl����H
j�V3�V�y_�TN-��_��m�a��"���+����-��k	�W(�B l&n�w��^��r
+�H��g��o����^"��&�e�8�U�t)��/���������$a� ���<̗��Qcp�E��;ɀ4JS�]+s�8+]��#���?TU��7�I���?���+K�gBǉ)7�÷���#*>�h��2�uK��wZ)�ճ�~���ջ\��ۜ.�l��$vk��J3�r��Mkb#�}x�*�H$[��ş��A%�����gc���g��/�1<��[Fv�,�y(��ˇ�F�T�̻u�IA�iH��e�ZӉt�t��iF���V�������}>�d����uY+���؄����2�.3rL��� 
'�Re���Ϝ$��U7��]���m��in
���ٶ��?ت�A��
����6�c�}D��m�%�pOf�ЅU�A��B������-��K�nv$/��.l�ce7��0�5�BI��r9�(Y��/lM�EfP[��������٘Y�,�o�܏��Qf,��p��B��l@��f 8�C�������U-��|����y��k{\�y2��3h��P���(��$����A�ŭ4���&����^`"YC$m,�$B�V@��}-�ο��ܕ~����6��!y� <1�k�W�̰���FQ*'��ʷu1�uAM_��� T4g���֧=�Eӟ�{��Nᣮiw8��Q=q��S�%o�>^��UH�W%*��^�d.�2�Q��v���]��D'O���,�v�iP� >U������V��@��`��%�e��2��;)	�;�=���G�E#N ��o+'���� j��Z��|y��|���:C�R��&)���i�: P"�+�n3�r�p�:q�+���Hu�x�f} e�Z��2=�f��^B�P�{{͘A=�"��mW����+��{Ūd�%��qҋgȅ�$â��Z�V��_��d�]���P��˔	�Tى���ON�B��f��a.�\�0��!y��~^q8f�Q��k�����A�b���4� ��Euij��z�k��нm�C�'��Ef_�]\�9o��V�y��� �d�oO����q�������p
"�r�7X����wګ��؋���E��jwP+<�Ĭ��xr�N���\d"��q�q��&�Y�z��q��'b!O\9Wk*�fm��t��->$]j�ʻj<дz�N��ӱ$3nw�fZR�s�4X���"A�����U�8�g%'W��z4��4y�Q�|����կ���X�V�HK�,��R4Bm{�+ٷ�tR0{���'��q�~�������5������p�'K0����U]0��w����ꏰy���1�c�a>!�wϤ`��i|�n�4��C��P�4��|�^	u�Y��h'O\`��[�Q���N��3t�����R1Z�w���]D�h]���'�,r���r_j���S7�gW�L��)�w0�_'P�L��`�&��c?��=�`�ڭ+��|fj<%0�~4�������������^�#�y��!�R��a��N��]�.�M��g��͗v$�v3�k=J�*�^p�>r`��ꉶ����7��\�l,��}�d'�#{�Þ������sm�1�7SJ�ǚE���W��f1b-�6h���`\�8+���31�\Qb�"�1��m���( ��S�/?��$�����Zb��3�y<�h}5�Y���x�$
�ecK�	����Ep�:�8��јVQ�_�|��T�Z��d�Io����03��4@Kl;��L�N��㧻W�3j?)��T���n#Z�YEm�Ŏ5&�#Z҃28<���*b�Mbz9Ϙ��:����B�˶����B�Ӆ�C�L�6�5��%�n���T46s#�xB���d�s�Cд��[`F���.b����R�[��w����8��9����k�H?�qd�_��L�/Xk.}R��
8�LC5j%�l�%���	�V�*�~�6� ���4��+䝖$�o�S�0��� �����x�����R(W1��Ch0?�-}:�C�E�z�#N���^�2+���_��d�cC���\��$�գ���Ë�Qoڒ7�%=z< ��^؈�;n��u��+U=­�1%��{�[QN}��g|�x�kq�P��K�b����k�|�����/d���x��q���کkPxA-�b����=��
[��7��k�9	��+q�a�ϠZ��8��ϰ�T��|�.}�'�}ib�b��&�>m��8혝��3*�%ypkgM2��ݠ��1y�p�֝���j�yS�,�������T���vk�?Ėc_�!�)#��j6���}K�y7	#�;Gq&�B3����F��Tl2�αj�W���&CQ	�"�a�H쨄i+7Z��/u5�/-�l��F�F����o�b΋E�
v�.��y6���Y*2�� <f4��R1 �[�=!�&ќF�%���n?	�ǵ��'��K킄�J#Nb��j��f�t=��G9J�[��%�}ﴥf���"R�m��ᬭ�c�ڨ6q���@�����h-ߛ��'����3�o�?šjE�vt%\|<Mxk�� �ۤ��� %���T
����0�wK �B �2Wo�k2��/�� NaԽ��+�g�V���ը�Io�%(^��S�W�l�w2!/~҄ĵ6Xs��!y�R���@	�T���#z���H{o-�Z�d���p�r�%��y�A u���x,����ؗ!6< �K��{���x�d�@���9���/^q�;�X�,���H� �ȳ7�C��L��LBF�@_C)'#=�#��Sv]J=�)�E���Rh�a��6h
����p]�Aʆ`���M��}Ͳܿ�jMRp�h{sk��̵���ꔄ|�C�$�2��{Bwv?����V��a1laoH���l���vw��h����5Z�:c�b�v����\65�Q������j�!G������Rn4����!���ㅨw���-�I;�G�>�~�� 1'Ġ���L�ʭ h����#[ ة����ȱ�^H�3]��nYH�B�}�L��1~�6~K�m�W���l���t�t�!���j]n��1t>*��CcnD��5L�/��j�,W�|�K>�C���#�g�4^�b�g��%?���ӱ�����֤t=u��H,��?C#s�����]4�_¡F�<R�L��)��`��&�����"�-!h��3`��_��y��ad�'���꠶�c�W����	ޝ�]-�'�loˢx�S�����$���`��G�.�Ӫ��1(��u� ���"�Tg�*��X�p��:�骦stA��nq!�z��M(�r��d��@�B\e���Ţ�{�3B���0�[�;Kp�HX��T���.
�/���'r�r]`Z�P�$2�T��������1��6�'�>B&��o[��ծ՘%
rd�O��wÐO!�q
*�B�?�+��q�GM�e��2ą�_��T�	� �w}���S��\F�}/b��$=����, �Ï{��C-ݴ"�E��~ޱ~d�֩6�-��V�>P^ff�����DS!Uke� �R�#CF1t����Z������6��L�� �������y'���]&�3*�k_����~�^Eo�����;��ǮE�i)��u�7�P8*UR�4��Ht�Az��*2��~m]���Tӄŵ��y����E�2�����h���R���VE.>ڔ�$�Ce��Keȅ %��֑�AV#���j�Hh���ި0݄S)�8�Oݝ;Zݞ[�� �FV��4�k!� c��1$,�F�c�$�/(v���D��*~:{����q'}-��MCuav�4���']6��jB>���=�>���|���*�(�5A*aK]�	.�[�E�=�d��-��OR��K���3[���""j0���f�@}�e_��17G��>�}\�3y���>�+~�Y&���q<�E�h�y���@��#�>u�2��~I��&������Cq�N=��RH��|����G�2��	��2m7�}9���S���6�)��3���)�Ƕuݘ^)u�SĢ?���)R��x�.o��8�`���>a��B���O��r��UU� H�@�ڲ}�pE	��h�1:R�����-������a?l������MI���X�#U
���n�t�y.�mS���Ab�ʝŔt�ȃ�?`=Lo���'�o�hڱ����[��N����s6��c
������R��	A�Ғ���X{���"��!���)���	>1X3�uU[����y۾�Oa���8G�$�:�|}��2'9:���-�3�X/��e�=�HfƯ�8�T�_�
q���`�ɪ�l�*���A8�au^d�A۽������=-�I��NT�y|��7�צ Z��l��6�꧟���1v��D��v!:����O7ŌS���s9{�	�%n܎��ԉgbV�x�9	��g�	I/�XC4�O�)�j�p��Hq^��e��]��x�/h�.cA��hp+�~�H���I<µuɆB{/�J3'yR��/y�yV��H���-���l���(?tg%�����Y�^�,�aj�f$�1�h���ϊ
�R��;��s�x[��D�HE)uU��X ���˰J�UEuK�>d�K��9)��?�jO�r��A�c��G���jX�����؈����n������I�+�U6���������o���;5�A�b�a����W����`�b��]�� ��P8���wLN��e6?	迼�`Nƪ�Z0;�\���A�S1 |P�Ǣnɛ��i�Ro�'�� l�]r���5�*h���"f�bG}��F	6{a���0��,r"��
�Jyp�8�#�P�n).�ݙ��I*M�҃.��yS�������'�dź!�B[[\��.<�7�ب2,#��*?�j4n��*���O�O����{]I�fQ��r�ѧ�i��qkb������`�^�תފ'�)��چǗ1z(��5�p�:���ic��=2,kBZ��LKGWeL��Ԛ���[BJA0*ԇ�Wp@j�̩�T�B]0�:|9Z�cR��Y�X4���Yr'9�	;�a�y��B.��l�5��mr5z/��������uC���Y�a����6�pQ��S�wEpj�SS��!j�Q�"�b�?��.``�v,��cn6W3 	=#�v�P�ό]�[��馔�N� 2�J�3a�ZB�|��+O�-�A�}���ݕ&$�{e˞i�F��~�U�>$̅�ϫ�}��Ep�����6u�{���cb�F�#��`��Ĭ�N �_^����"2�_}rA؊�F��	h�Ŝ��`&�NOr�>0[�*���㚊�� � <�D��{��z�O�У
�y�,��󿉇��^�7% D'TN����?EcR��y��3���N�y���n��pF��Sʭe�ä�R'�ޡ��x�W�	��b	ql[S�S���w�C��㞢�{��� �<F��N�x�5��qr�%���ez��'���_w.j�_]��DB�#�^0}+V�#�HZi��_0u��`��~_��tػr)��6k�]�o�踕�4e����7�Z�Q���SӺ�ur*�)GP����/�Mܓt���o^��p}���vyh�0�-+����!=��C�R�-�S�Q4���������Lc<޵������h��C��\k�z:D���7���C�$t�c�By�k�k�~k�JG��T�7�W�kث�J7�У~�{��V�m��	8XP�?W~�7�~�)Ξ�B���^0\ѭ��F� �o��x�pY�m�9�`������$G:`
(l�2M����%u%](�.���t�8~��3��/��^�W�̘O	>��R9 q\���W���*����U���6�_��Dj �C����m"�!�=�;��AѠ ����W �T��r0S����6q�Z�8��~c��kB��+���:�RŶ�6#
Al���7b�qE8l�]�t���q�A���8H#�㬑/�7������2,�� �Ô�*4ޢ��4͈X$B1ܛ���XGj�K��aW*��C��[Ho�\K*>�����֤�>��,.������H�%s!�+Ma��PG�d��^.n?��'���Ο�4g7�q[w�!����`h��ߍ�-3'�ie�J+V�%#7�s}w���SlƮ��@3�x������h�e͕�s�y���d��c^ɋ�����1粨
��y��(�s���ݚ�7.�%4�Y�vf`r�O����i?ӷ4q�#��	�Π|4�Ҫ�K�OFQ�_0G�!�Sl5�v<��)��`��`g�&�e�B&�A���r�>sL����a� �X���>t��.�����3�Z�!�#<%\��[k�O7�Ī7�ʺ8~_K&T�)�J; ���f���ϘN�O�OCࠢ��x}s�b!����Y3��A6G�E�U�O9�T��
<!g����"~2�d0�z���Q9�̡n`��Ҽa�$cgI
"��}m-x/���(@��Z����o�q�z�Z�ţ5kA��/@�s���n6����������w+G��Hb�}�YÄ��d�����&�mw��Ѩ�D�����0f�/mb�����ꤟV��-����-٣M�@N,���J��{Ǎ0�E��A6�>[=��b�rq�6Lu�w����@9F	7��`Mo��|/W���'��:�:A�j<J7;�8Q&�x�R>��^Ò փ rL�ś}::2���F�q�\�Y$St���@h���w,�N����l��y���1K�E�	u��#!��  �1�q�S���D��t���#�^��׷��>g^���4�!�t� �^b~��T�9��1�.g�\�0ʡX���8N���T�b��x^/�Ղ|�]�A��ǞDh�/�pK�����zWG�X��ۨ��)Q(]!$���'��W��ץ�t��k��KEO�(`><��>U_��Ux��t�Ů0�s�rL3n�g�J&����-�����G�݇���|�Y6:�bz �(ٹ>z$���b���x7S�� �^edTr����n��c��!��-HK�㟉�<�Yus~3�:��YSoѤ�~iyF�[j��]�CN�ZZ���y�wiH_�5��W���G���4����m�5���4,V�H��\Vs��������=Mn�f\_��F�(�C٣�LɨT�`�� M�xh�{s2�)w����m�Ӏ�K���7����r�vr��t^6��#p��V�զ�R���o�����Y1�����м�Lp��=�a��i-�/�����ie�N�PW���V�z���s��Ν�X��?����)�Rm�Z��ѥ].�6�GM�v�X�$��◉�B0+<�k�6�u�1/] u����l<���Zo�=���l���M.���3��|a}M �s����1ľ")��L��7d+�e1s��}ΰ�oױ�ʼ�����ݼ��
����u�-f�������\��{�����7J5���I�Fn�\����1��H���Z��T��
`�u��GZn4�*���t��L�
�����BL�x�$�͡G�M��;A�K�8�S��WzA<�
݋V`�-��ѡ�0����W�63�'��B���K��|T�� ���C�-�"��Z������"�;"��*b��1�;�!��r�>��[�w>zpl�V ! ���k��u�x���Cx�z^vqG
����t��UG��ږ�:j�Z1������_P��XB��]Ζ��k`5�7q���Y^8soI�- �ը���q�Ƿ��9$��\dk��k�[�-#���Р���ԭNJናP����S�f�I7�h��E鱎���,�N�{3;�[걤l����m8�vQ��n�Z��T�������S��9.<w��T�!�	�/bX0TPX�����ۙ������?�GpF����
cV�zp| �e*S�:��1R_X��2g�5}1.�S�c�80���];�������@��n=��.4��O��X�*A��4)��M�H�������c��/E�%E-��Y��2��Ӡ�� K!�µ�k�+�b�e�9,��R׷�����e<� 	KeT�2��n�c�Bpg�1e�EY�WF�>i�os[8�u��	���yc�M��{�<I"�O���L�A��di�=�B�4�r���R���I��Z�"�a����H�5Z)z�U��A}Sx�찟�����R��W�|a�|{�"5q|D(� �W˱��?]�&���zD��<|��1�	�:��3u���y6qmC�r�����ڈYz}�wk���H�%N�e.�@�
{�1~蹿<���F�&?���ȑPI�q�$��c/���V2�l��h��ĕ/��VöG�.�avp�
91"����$R��������x5�F���`�<K�Ϥ����3���D�}f��A�)^�a�ޡ�b'U��=�WE��+G@��T��Y��$��4ޕ1�iJ�Zޘ���*@�����RZIp���"c�5+]3�w���h5Г��Mf�1~���V[cU��w�;�DE�2*�}F��@oo���&���SM�xb��EN�`GO� Z��)���n��.n�,���ܴ��F+Bii	^�<n�Y���.�=,K�n�zg�������`�
@k�)kp%On�D�<l.���M�$H�8_�`m븪6��{Ξ��-�#�I������p�gMRR6<�W���U��t�!�j³�=�?��`�q�,���
Z��v#�Ʊz@Ě2OfDά��mޚ�ݔ�*�"����|oS3!;���?�i̥�n��9����2�1�LI�f�M'f����$�����-���1�B$?Q�L�?��
	�� 
vLn��*cY�sB:����k�������HԳp%x�F��@*6 ld��V|�n���i�_z�[翊��TT��(aj�%^����0�o�FMx"r<�L�Pj#	r����J�!�<�_U�m#'Z�~JЂ����;�2#�72N�p]�ސ�����u%��L ������tjܴX��MG-@+Ö�=.�G�<�1��׊���q���i��<f0T@p)���2��Y��`�&4;�P� "�f�w����cX��ą����g�
Ef*0����}�T9PMx�CA��h����$ Z��S0���K���Mõ��H�0�S�z�!	��J����Q\��7�h �r�hM��G�����G�T&	�ӈ�[a����a��I�����hTٕ�J�W��6;������m�ՙ/"YB�/1����DㄑB����%�>k9�+������=���& .��j9Vi7Zw7��F��la���`!�>��Y�=��yG��@�[����t�VOԻ��ѐ� l�UK�^���ğ��h��v\bi �A�t���L������"($�E�B5_~��4;�̟��b��Kp��}<P��7\,F�DH�?}�������� �%���
�2.?�q*c��w��I��]����� �'r8�(�]qC�����LU¦�70�C?V�N3���A%��j9��"� 'a�:���⸲�ǔ�7�E_#�~���6�Q@`2]3�@`��;��Dh;��y��'GU�|縠g̴�h�	fĠu��J�ZxOf�軋L�e�c�JF��[�����{��xP�Tu(d�t*>����G{�7�Y���[�[��:l������)��G��$�}g�$��~�YppR� N$kF4P�|��Ea?n��?��Y!6�x+r�K�����ʭ�r~=�P0��a�z�Z@�%t�����I����m�~g�
�5td5X�g������';n��R��T����.����!ZBr2�BW]�����,���ն09Z�8�o+����c/RD<S�6b����� �*ϗK�ְ\~�e�z�◍�f��Q�Bs�U���at��Ю�N'?�
��oq`]�X�!y�x.hkjpW�C(O�+쪊uVh/��%-tJ�Xx@"O�JÇ£�;-,oJ;��$_+�CNGa�(#��"v����R�aP�dC��d�7ao���Sj-��8|���H�u���{�>+c'�ܙ��5%zc��F�3I�4* j<�yۏ������B���cv<�f((g�kc�6����`o��`���<�Q���!����'�fX�ҹ�!���֔ȞiPq �m3����ܱ�	@j�u�����-)���-P��ߚFi�9�vs(��}X��#�,�� ��mP�_5�<p��Y����u��<Ka.U���+&L�"��\"�2������=Aa᭸�7���0�˟�<a�R��.w��^�k,�@H��[�4*�l8�Ϻ�y'<=V����U�|���
9�ř�$ߟ��w�z3@���y%��}m��T_n�\�#�X6��^o78a�R�W���B��xi֘���x}��ْ�>��m�fg��m@5�g�U|�Җ���P�U0�%D��\�&�0��<����ce�W��P���a*|�v�}��(L�<�L@bQ��
�w3� z�<�]���~�.����^�mx���P���0n�'<����Y��Q�G�7�����1�n�¾�n*6�
��S_��j���њ��[�G:g:��c�vG��e�?�,C��{�}l�j��u$�����Y���b���#�h�jZ@tiT��!mUt�M����	���I8?�b&���މ�|y`�_���?7s������� Q�?J��ܣ�~a������E��$�ˆn})}A�=��6��'G���ꢚ()���_ڵ���S0�n6��,[��@ߟ-�k�����A���_	�a�ggŜ�y�W�.MPJ�ob��*,���1�kohe|~594��#7AT��b�����H�6Eg��6+o�Ƕ��d��<?�}y&$�qЅ@�N[ *D��C/ZF��\x�[�2�Vj�o� ����b m��i%�_��cis��d���n~aAk8����s�r�s{�=V!�-�����a&W�Vk(#��b�������8���Z#촣b$*"P���7Z{�o���`�+x:m�"��RÒN�>u�i�0�j5m�*@�K 3���t������~���QeC����/�)x4�������e}!�7~@,���7��"�5�:�b�)v��c���{;��]4���y㪰�b����S��<PB��0�A���2��&�h2�kE������n����"Tù2���נ!������Na ����C�khTn1����@���Ǚhi��a�GHd���I�8Io=%`���RVK�2��N1R]��8��Y2��Ma�N�/�;�r�iث��q�*Pl>�ݑO�hKٌqt:��K�r19x}���'e���1�(��3HP_�D�g�%�XvA�����h�<��1�Ξ6��5٨��[�>�]�0o��㨄}<]����[V�k����[��a�Cu>�@s	����iH#����������:W�(p w�I&w[Iq�|�P6���Iݶ���h�z��Eߠ��O���+�Zx�^�*���2��c�ʴ���$�q��Kc���&�o0�u���;�2�Y>1��%�L'�^��QWeYx�s��e��d=��x��$�do�[M؇�,����Z;sOX�ٌ�Σ��;��� 
h��MCa_��3b�a2���`Cd�QI�����I�l~O骛�m�����ڇ�W�S�oyU��KB�94���nG�?X헇��<��e�fGQ��٢Z���Fc2h������Ƈ�s�H�������[,z;]��q���f� ؁DA$_J8��nnZzZ��Ɲ��!.  ��åA�B��D�F[I�ܡ2�Mu�������� �`R��?���F��w��%���j&��B�����+Ya5�ڮ��I���2��L���+q	��i�U?�c�I���������'�9����"O���}ʔ�(����zF��G��]��;k���je�'�g���G��[Y��wӰJsX�B?T1N����� >K���{�wB�w��[c�De�l�p���̦*�\�o���bK��|���!�S�B��~qf�g������l⚿⸹P��@ɜ��	����gQ  ۧ
E��q���I-�:���mS��/M�ؽm�x�KI���P�y�����%�H݂OK�B�U�G���j/o���������
�|P|<��h ���`2�K��Iw�*��|\0G�#r�o���_���[%��x�!z؄,<��u�����P)6W��^�']������ gj��s�Yq>Q���4�J�g���$��z��6�{k��� Ԟ���^���S��ц,a�Z�?�q�V5
�u��� �ReS��Z!(o����vb0�®
r�Ab{�0a�g"�5R�63��{�%	��=�z�6�3�lC=*v^�U�d�x͛�9�`�,���oF���Oh�>�A3���C��B�Dw��ˍ�蕑��}���k�h#����-��;�)_)��	~�YM�����@�\ø���7}��e�p�i�D��.r��b�z/%f�.�ɀ"�6���k�l�eW��=�7�^X��|�']�\y��ɋ��m�i� �$7w�ipb�Mj��ٷf�5X(_�.�,�{���9�z�c�UU)�Wm\V�"ݡv�B:�S
����TC�!�c�=H����s�3��� V�<i�8����J �H5$�4E~;6T8~���K$�}n(�`e��x`	�5�˟��&,gî�"$�)�ǋo����Y# ��Z��9�~{nvi�_؜y���mf	~��i/�� Ww���M�E�����ms�N��f
��~9����+E-}Ծe
s��g=Od��FQ:�c1ܫ���2[�+�Uژ͵md9���[G�Q�ڤ����J�y�#V<����[�����C�<��������࿵uL�8��:U%*����($�r��wy�RM�W��ܛ�Q�Ǎen���5bK�e��T�xy�!�X{�޳��,�?�J	�>pb��[�mP���(ƉE<d%l[��Uks���
���Vܐ�"�
�_�.����ٸrD�6nw�׷�Am�D�X�%i=0�$�]���E<��M?l��"x�5�Ǯ��?=���Z�-<v�NTgn��MR����:�Vebn�jr�0+R&�"�#����q]T�%{� xD����PM 0ڼ&����`��7��Z\{��Ay�=L���x�Bz�܍eN��W�,�p���ʚ)�m���:�
Jϔ�:�oD�o��2|����]k4�T]�Ng\���ߘ:���]|�8R�D��僪��7+���҂����Kt�+��?X6N�?��o��|��%��@�0M2�1!xd�P?Pa�&=|�_�>��9��G��D�N���0&P9��o�|����(H��R-�؝���Cbyt���+����d�����-�F����iA�f0~��5V�3���@��N�DM�̀�#�.%/����9UI���?�[��0�%ft`��ק�I�i&_�X��P&	%:��,�@"P��CהϽ���&�E��h�@d`gw�5�RŎhe���v�Cj��&&��� l�g�-���a��)��a�*����ntTӓ�afצ�U�h�O[؛�\.��d�ø�3~U�i��r�[�g[P���z	4W���s��4����"���5k+(9����q��������2���>a�K�	o��B��3pc��_�������+��_'9�$Hzv&0���f�ÿ�c�s��D�+:������ �s�I��@.@����\'0�N ��-���:+3�K���)�ɫf}?��qT���dz,D��L8�jY~�i[��xjzd�?�"��\yS-QMCc�k�A%���&}:eZWσ9 ��{�6�'�4d���(xV��E�����	�C�GrN���JP�gK���M����r}e1<�ǣucu+fK��i��B�A3���ZU�B�S}����X�Z�"��tt�(>s���fu2�>���k%�5�s�#S�Ţ�(��s��t}~�Q��7^�w��C�#g�m$K9�.�%�.�0@��,$ڟ���`cBЛ�s4&R��O�0<]V���l�/ǀ t)�5�RP��Wo���
/}��Մ��净'��`�h���r>�K>EH��:H��Q�-G=��[ �	��l2�V8���� O�Lb'q�!PC@�H�M(�����ǵ*�����6L@6q�<��>�v�GP6Q���a kˋ8��>�ެ�d���V!�B��cW%/�<C&����)����w;�,d��쌮 �8�>��LD^a�FϚ�o�a8�5�*ll+���"���������5�&��F��~�L��uQM_���#ʒn%��y��(�6
w���\��ʞ�-m M������D�wA߰+k��?o����e:ё(��9`|�p�9D==�Z�E��x�)�i}� T^�r�\��ds�N����4�e ���
���j��a�� T�9�h}WY[���XIu�X����K��?=���9�m�{�S���KLz ����W�f��S�'�|���ڡM������)���LR&��\���ҥ>���үXֻ|I�p��4�\x1���k��]b~�u�����K_����{1�O.��y%fS�<�Ϡ%=r|�g��x7V���̎�@�@6�>\U�1���b��{��l'�8<D�QC�zZ��MהDn=.����=��tP�a&MM�A�wH渆[rma*$?UpF�OJ����/ҧ�	�ׂɳ ��[���g+�'���;��[��r`�%���2~S%��sʜ@��/���O�0����
�>�ԓw�D�/\�51�wO��79YDg�-�S�E4�5�V\i����nn�cL]��s�z��RҔ���efL�$k�f2�,B��Aa@���g�7�7%CG�v{��#�n��	�e�5Vv=:yp��cd{a���yt�{�^��?$�P��������	�?���V��~B0���S�P��{�.5����8aL�s��6ϼ(�}��l�S�"���� n��ˤe7�������U�zf���Ř�O�����{h1z�-FO���i�r��.��6KB8�䑑���ց�x�N9y������$�.�j���;�j���m���������@�̂{����J8;�6ΞX�� x;�<��˴B�F������@ʻ��`6v����@�}>.��=�'ŠX����jw#(�Uѽ�|���J�U,#7���][1lIh��t+�`L�������ב�̹[\Ղku%̴v�4�ee�}���\S!c�E���TL���?^l�n|H�"���u��@\?��A��	�U�L�����7�gL�B�p���5`�L�p�����sI{Ot�_�`��o`i�Γ�M��B5Z��,f�:w����b�����n��-~*���t'���Ì3ŰD�/2��+r��]�=�<g��#	+/��t���0���2P�S ��Ib5&�t�KÍ��y(�|G*w�{Ͻz������'h �f��[�;
��	��;<<��Z6��[���N�!��[�C�T0��q��'z
m�9��E��ϩve *��Z}/0N�:�ir��;�e=�M|�S}�'�Vm�����ӎ<M��qS���yMܖt$���
}��r�_-}u�CU�a?��L���b�\.�7YC�W�j"5N���:ȝ1���>�Bl�rI6������C۬�ͫ_%��M��"�G�u�zR�1^#8��P	F�Tf�N�(�J�sb$	�����Il�8(�����Aky��Y�i���c�������n����\8�B�ٶ�a�r�7QY���o��4F�B�;�Kb���3����4ʳg�z��7$&9��Έ  E����Q�e����iw-�/��-<s&ʶ���ūp��(S�F���P6�-&�b4�-����{���(2��0�j���G�b�����C���M����^}5�o�39Ņ
���z7�2DuE1pD����'`+f�h��OfBm��`燋6�b�lǵ�9�	2���JvY��� ���+�S�� ̃�侰��}B��Q�� P̡�|x��x�a��峘Ja��O�� � jQ�g�&�3�����]3B�_<g�I��F��ph��m�hH����(AD�Cno�}��N� l�Eh=
� �*���aJs5}깏N[�3�d:�,���/�����6cZF�[w�'��M�>pKJf��8N�`/��P8�oq���:�Z�d@7�[ʁ"���m]~���oo��:I�^n���Z!�LB�٩l�j�%1X}�7��T+��Ӏ�#���Ƞw�:yW'[��무�:�Il���a�q�
���]L�>}�&��D�U����	��}�������փh@��V�`�����Ywg�0z�LZ�m�5<SQ����Щȴ�[�pp�i�V������ �x�ݒ�<+�Bҥ�_o#�
���%����2��e����5�;��� ����S�Nda��22ţ�]u2�δc&0�����'l��Z(~�_�> ����L̓�J�*%c;s~����tJ�඲� ��pN�+,�Ө�.Fgà���\GḪzWXƸ?R����Ŏt%�9���L�c(a����4	��5Ǳ����x?�דҼ�_�}�S�j"������RʹxT)��QBDO�a#�U��C�i�D����цN�6�����	�[b�1�N8��5�������E 8,�� ZP)����U�b_c.PD��$N������9�����@o�a*�����P�f���B��ֈ�c��',(�z:��z��u�x��a�n�i<�,avꮻ^�-ٿ���cJ���]�TW���,�ʨ����4#���!�}yݣ�	Hpq�(4x��^-x���D��?��xl�/��(��pjłpD;Q֠�\�ǌRj���toVm�����b�;I�u�u�΅�nqZ%�GXke-I�9���J
�M���	{�c<�c#������o���50�n�����
�����	iרJ$��?�ԯ�8+T'4��;���U�M2��N�pS<jgٯՍ�ɨ~��Wp�9h*�n��l�}`��������O���M�̶��L��X���[T�c�/v4���w{8������Du�l�8���a����Ns�[�7K���7ofE؊2��}��$_K31+���?a+���օ-���	��}��*�����F�c�Bq�2L�����&{&D:$�iH^��#��oqiщ\9�34�ZCH@�>�#�t�/�� ��ڤ�����P-4d�ՠ�W�}�g����P�<k���MQi�:�nׅM��n�1��=g7֖ohC/ђu��gp���zP����8O�{"ڀ��/��\�����P^�n~���3C�
�\<�{բC����Jʐ5�/��b0C6���:�F�`w�!;��5��7����^0F� ���ܧtd�h�纳�C�/J����Q@^��V�e�b���O��3���>`��4L��H�Sk�����?�Mb��j��7��	���zη&2>B��1��PR���.�Ӧi{�=�Aǖ;t(4 ����'�h, ��]��y���Ytz,����sC��RM���9�����i#7f��(��dT�Z�����t�RFY��-�I�	Z%�Ї7���H��SU���Bq�^ͯ�Y���n�F���B*Dq�^r]���	^/���<��L�cQ��!_l�so��}�>M��m���z��s"�<�k����I�޼ȡ���Y�D�eOg&3�ָb���(l~_�M���P�d���+b�)>Tz�{����ɂ��K��o,>ʨܜ/8,���M�DE�S����ݓ��mHX�l�Z��M��x�	m=�,FҤ��u��� ���Sh\� ���Tt��@]����_,3�[_���@�3�_�WNu�}��$M�c��OAG��A��N z�i���������K4�[��i3�ER���IԦ٬�CT���c�-���%��5Sݾ�6���y���0G�%R�F�E[Kx��wu���Ã�S�g��tx:�����n���2� T�թ/�� �׭�&�]Y������z����
ɨ�(ť���B�Ws�e��e\_��l~�$E^D>!��[9���^HC��N���EbO��ノ�?!t�2{�FSd	h��P�d����]�&ۓ<r����}*�=��oAY�l���5�^�O�+vQW�A[�Z��*�©���Qc>Tt�5�&�����Ui�×.���hѢ��}��\o/�1C�����$����VHNZ��Dl	�Ԁʼ�v�����;`��4�ѤNᇸ�u�Dʔ`r9��_���i�t{c-4�h�U��Z3φKz�Ɛ��9�1���&
�9���/��Z����쪎#k�v���
��1eE�}{F;T�2�w
-�8�ٙ��h� �3=���~'p_'?n"!~���ݗd������$�]���~A�VpO�	��8��eNN{Y+% ���lA�׭r�Ǥ�C��:�vHi9��&��	��$B������~
D|9Ջ��0f	��<�fB��O���D�м]�a�F�ގ����N�}��gl:uy�e?+�NFW�#F���U'������;��|�+,���VF�X4��P���aD�j��_I&~���Z�gݘIM�"{��j\S�`���u��Dp	D55�>.9<�n7Cr3�S��G��>��5���b�N�����ڋ����Z���Dg�s������v�Eê�ə��"�a�
��"�IC����*2X隅�^����5���?����A�*K���w��s�^>������ӹ�ґ��!�#����.�:�!G�<��a��<K�����$��0>�R��g!8�ǸV�����
�7�[ſo~#4���ک1� &P�|��z���{F���?l�5j8
(�� ;o�+_S	/��EqV?��x��y��YS�ܙu3I�b��>$�L{�R�Zg� � �NV%�q��=\�x@^�w�Wk���StK���X�9q��J�/�R6�<�N,�R1+l�8~�ӡ��]H�0.�>E����3s8�7`�)Fƾ��)uЫf��l]�6[,���aW��B�BxP���ϙe�K��?�E#OQ����BcBQ�_���|;�0'�}�)�����Q��Q��k�D�}�M��.��ٞ ���`WAW所���M;&%<��Δ�t.P��M�- �@̨eC�>�]�;܆��W��CE�eyZ�';�q<��=�_pz�D�T ��q��J��{1�w����}r`�q3\#D�["o%v��uG̴h�-v���]���؁T��	~��-�P��t�*ZD�nV�S�:"_�|7�1d�d<8ڤ�2J�KE�/E��0�=ǖ�gs72��C�י��	�������a�z�\�����]ä�YQ$(�ՠ�æ�9����џ"ph�"%�4��I3Oy����Q�����z��hk[`�q9���C*:�M�~4�e�	��Ǯ}s
aoИU��j1~zk���xK��5���$fX������A�!�XQ�p�A����ѥX1
��)D�Q���}�"��7	��	���m�q�8�W4��Y ���!\�z�̂�I�y����]�϶*����(��J[�����W^k%s]6�r����Dޅ�>��� *ua�.p	�L�"��UV�]�n`�i>q���6�s��%,(ӮJwb��b���
O���&v,�h� L#�U�[z����h���rA�y`'L���sz����f6�e���
�ޑt Q�*pH���V1dT�9H��%�,�r�Z�qϫ�����0F �X ���GS�+Ҁ�~'��&�~(RW�P-]#s���LƳd���mj����X6�r�a��5@B�B�;-64��v�;���|��B���(9�Lc5�gV�$�  [ f܎f��~�
h|���a�P[�7�o ����==!Bʒq#N~��� ��bO�$�������o}4�>�jx�v���� D�� F>2�w���O� �\.���E� ��}r���3��9y��~��\JJVJ,�(�c9g��q���DX�%�o��L_C�s��מ� �o�b\�����h���>�#on��h`���"�)ޏg?�aBG��_���G/!�`����0����dp�C��^qk	b��U=��\S���_λFC���z�"3�6�K>T�K�ye��+`oV�yo��za*�z���Z��'��1�r�0���]yu�Y
aO|� b$�n����K%��%��M -��A��6��`�9X=��6%X�Uk^I￱������į�QeԔ��Ҷ�u�Q��Ԡ8��I�$E�/z� ��A�{"�J�D������4��ŋG�U����h;@$��yW?o�	���U��\^�n����I�3�n���Mo!���%���2�p�͑Αc�U���V3!��`��o �T�K΄��(ȱf��H�Z�#
s���:	wG�u�$B���R3X�l�����߿h̎�]-6����`��+�(F(�3�~���o�#��r���^�g�j�$w�`��7'Hf���y� �m��Yf��^��F�߷ͼn�d����A�����/
�Т0$���p��
�z�}L�L��ssq�n� Q��-Ôv�#Τ7��1*�SW�Ġ�w@BH��鹺>+M������1��LC��06!�>��}�����y3�M��[^Щ3r�����L�� ��Jy��O�:�H@O3_. ��,�%o���3D�~��*�B����s�1�x9���͸�n�4=
�3�
n�+v�ܒ4C?7k.#VU������{�!0!G��'�LZ�Y<����㙩�_�e)�Z9����T�n�f	���P����7��C�4�e&ۚ_�ʻ�BlNAS��T��;d.���hOP�q���8#��m���E���o6V�+�vm�6� �H�{�C�̈́���i���{Zw��"��#T6w��sh
'�r}�s��S}C��;����O��B{���YJp��1��#�����F��.�D�S�����E�2Xq��!2dh���5�޶�uS������K��^ѶjR1�梂C�����槡�Ա��y��:�fhB�LgY��>qOR�E<A���B��(����j��3�(1:ф�T ����1f�O�,��"�r$���a�z;�"8쇄ؕ�ݛL~�e�`����&��c9���]j�4�k�l8�`�p��O�	���Ѷ�kj�c�2ƀDB��ζ�G�̂��`'\�k�j���眿Bl�V~��B�؃�
�(�C�}��s�@�hiad�; _&�ȟ�#�-�>��ǧ?��o-8U�}�Z�r4�k����G��F���s��ω>�k������슘�I�ur�g���\�6�i��1Z"�ޯN�s�w~Ɠ����O 8h��ux�[���wAV?T5�^zQ���u�֟��,�'+���H�2��:��A�Sb��\Б��K�V-E�1�q��S�x�{R�&��Jm�pI(!�ޔŒ9�}p�ͳ_r��,�k)�����+��iFo4����y׿}���(�*v���0�G���άK���1�:��ΔC�˰Yr)���e����-�3zT� i#Uh媭��:�����D���`H��.Fs��;�R�Q91�C~ў���,���.�Z�ښ�HihRs�z� Ԧm�'rM+��}#���~��.��6l��R��go�s�2�t��3f��h�Z�����GD�����|bn���Ⱦ6���Q��"�i\�~�K�麴x��o<��A�b�Zx3�܈�w�Y�5�,yU���H_�/�<��r^-�榰:Z~>h��P_��
ںp�R�����2%�?�d��Y	��4#F��-~��'���M�5~�2���y{����BA_�([G��G�z�+�w�����6X�A���~�j<���� R�3�V(��>��/ q��P�#�bm2ʪ$�Do��1�x��N��~to����*|��q	Hy��I��>�D�Z.��+,�U9�艞��f���Ij�OJ	;����wX5�m�.s���YRF���w�Fl1x[�)�SX�a��^�Y��(b��n���q�6��G��S�0�[�eC���=�H����JD�� ���P�fc_�X�!"�t���*_�4�'¾;��`���3X!����6�o#�~pޕ��VPK@�	W-���ϼf��Ъv� W��zd�p�� !��e��/
6}����mcB&����O�+�t����`x(b�Q4�K�,ϊ�h_�ʧ$�i�ڇn���T��I��t�*k*��>�8C��5�~Qq�E{Ƿ��t�>d�fã.��v]u$�@���M'�h�z�\;�鈐���ˎq�
� �|7�-Rũ��[N��ߟ���'�)J�2�W�5dj��0$��"B��.(!�|u�U!K� 5���1����e��`�O�M'@,����]��zZ[L��H�V�H����4x���]/��"�40��'5�:��a���Fե�����5l����`^��}tq���ѻZ�(Ϡ���r�W]��DM�	^GR�����[1�w��{�Γ{R��0ܛ��(��K�Q��b%�A��Y������P�G���/l���F���^�1<�.��>Fd�S��	 �G����;�,Ev���m��A0�N<V���3��6Y/������ �p�{Z��cp��C������^IB�	H��Kl��"���ܯ��ߕ�k=l̒�� kW��}�}t �#���Kh�=U��g���ii�s�v�T��/u��l��^�}���7�yc�S�f�((!_��;j�]���
�â+��
(��a�?�@��꥝?�K%]X��=��y��R���j;������uJ��t��0�|a��D�ۏv����%�8�"�p��ܮA�}�r���h3�o�rAi�x"Ѽ�ch��9�%B����k	�+��V�W�^�������p䮪C���@���5�i�N�erm�o�~�C�b�S�q�)�P�n�)��e.M�U
�LO���EO����|FF�H��d�X�F;^��O8��1�c\�����w|{X���H�iI'Y�}��48���������4-�y���HI>��>�$"�K���L���K�����0j�P1빧�SVs�(2��m�z�d^W5�1杹�c3�[KG.um�詛�F�i�kݬ�-��E�3�0l^��j��!� �H#�-v��^�5���<i$��v��������tJ����qep!��/���d2�3�.K������_bf����8~�q�f�Ԁ��F�ʮ��F��n[Mro+�!s�^d��Ғ鬄w��9d�"�/�3�d��B0P V��su�'d�KϹ��U�(����JDƋ�@'���p��U����y 8`xt+�)�Di*�ݡx鯋5��%
�0�M2ܘ�U�>�?����=T܂>~�].B��{��λwz�U�-��
��ջ,3���5
,�V� a�1^2��4��K*� M�"��d�U��S�f?|�di��C��Y�#��_��� d;'����B��{�E$��?%��ж冲�KU{v@�e��C �;$��-Da��}���u�\���T�>��P�+�	)�83���[�5���Mj��̶ɍ�T� ��
�_d6�I���FzJ,oe�<��T��I3���m������OM�É+�Z *P#�q!3(o�J'2���^e�r��:��:����}���^��xXE����� 	�)����Y���(��	��4ZX�I�#�Q7�����2�y"Fg�H�òA�V��KHO�ű��E��cqh�2@�}��=�#s#b]5����j�xTO��I?��-�5��L$�wGa~0��4���l6������.��np^�F��?�C<%����?W���&h=��G��ɘ\P9ᗔT�G��y��o��n��ae�O)����M�%u
����g�̐�IfdHb�,'u�w������Z��*��z���8|������+�$	���R]��E�E�2������pȱ0�:�]��B}�� &(��	��������e��=e�;�(::�!����.�ws�TV���F�p���#��j}��I�<�%T
�8"2�m�}�Nt�8S�AB,�J*�:$��W�1��g+�� c�.�y�L�Q�m'�A��� (C�|���
?	k�^]���̺�YW;�:���x;�:�:�QB#k7�B�T"tk�7Vr���ǧ�X�I%�veT}�@�aѽp�����G�o���Kg�߾k3o ��<ql�2%sKu� ����C�)>���f4
���PÁ�3����3J���/C��#h�:�t�.�8�ɒo�7���֧;魽�\����������4��q�V�����E��H d`P$�U'�9�]����[�6��s�{�S�c{�p_	I/l��D|c�,��T�]Y&ә��« ʇ'���B۸U���r��<�תH��˩��ث?��aI3`%.퀩�)���&�%�ђ�E�ҿ�Z5G$X�M9�qF�E�j�n���4"qkgG�1�׮a �ϙ�F'�#��;�7<�㮤 �bB>�4(�ˬ��3��;<ނ�S>���!o��U�1�l����~�Z�;jnjB%N��T��o��zpaw��zjL -�+T!%�΅�M`��4��S7B��A#��P��Ť�b8E��L�E��)m��	y�� ��g'n�-�S��o��.}T�θǞ�]d�r�,�K<h�
��|��ǭ6H�~֌��ךJt)��ވ��i#b�lIF-���4B��Su��]�w�ʮ����Rt���mb;����!�ru�倿���+ꚰp.�k}��@mY��m�&и��Bw��g>��s��{���=�P a6R���Y�4Z�v�^N�K@�J���������N��1Qi����C�46��*�
�a��#&�@�;����,�O����zYp=�>�.��?:8]E�͉\���x1�~hC"`�L��2�K�l\�ȡo�RLm~��)�w�m��K�a��;����)��Ȇt���ǽ��o�h�e{ŖiOLv�_A��?�қ<��[��?�A����~��8Qz�C+���
�� h}U<m���Un������Rz����~̪b���/��v���x�f�?�g�6HU���T [���7�)�/�����~'��30M�����%v �
��M=��ܮ:~���a��?M��ԙ�Y��9 �}�Jp�@y;	�G��	�*����[�4��W���fޫ����JR���^לC�ٹhJ
�j�,&��Ε��Xp������3`�R?��o�K�Α���1q���@�Mt�7�8�	K�����yY�
���"J�SM���@gR�W;"�A7�����<1l������f���Bh�ן<��`���r�/�pO�3�^�q:�cZF���p{�~�2����>��9�To�&1�&ԯ�ȿy�e��Lm'l����P:T���s�T ��6+���$uu۟
���R@�'=��|no�~w����̡�P��fP�e	izgz�T��s?����0R��)���Uw�x�O��o�����5���q|����q0�6�9=��O@g8� ���,+@��(w�'-�X�՝��dkQ�
�kc��[RC��DK�ʬř�<!\Q�B��V�D�6STny�h=���۩�e��rW�h�Y\$O�n2��p�uV1���j����_h��^��4$�h8�����Χ� �l�Dwxj��8�-2B��H��\<LO�	��	��5�^F{7ZM�����%��4߮]�X�|�ꉤZ.5�t�r^������-�	�v�A�+��!�٬|�n�����~��PA+儬h�2����.ߢ_]��w�t�tVr8\��mX��đ� ,�<�, ��\�jg��n��Dq���>���w4��;2{Y��_ߡ̫L�z�`8���;X �HWS-n����S����\
��~p����e���'��2��&������!�>rK����z�1W��7�ƘG)�^K*�D�H�nH���r���2^������?˱����O�6�
�څ�9����=�ݨ�~
WU�P�d>t٤� Ud$�l9�վHb����3����h�����fD�i�
���n_�m��<$_����&���y�1*��KU~L��ȼs��3�!�S������7�@(�ľF��{�B�G<`
o��qM�d���U\c�l�:$|Ql�<�3q -�MQ��WY�.F��� 6L=9��5�d��ˀe �1��f�s�lbd�@i���je����1�k��;���(xҙh���������`�.�m�g�عw�W4	���ˀ�Z�J�_bZ�hP�3�+��%$��ȳuU0��DoՄ�Zf��S�fǱ��2st
w���tN�;�e凡��6�arpdB?�e��!Z��1�/E딷�K�w�f8h�7�S�f,˯�^ٿ�LSX"D6�SO�̓��sM�z/��B�u�&�����`W������C��'�&�~��H�_�K���+�8%:Ĭ�����ָ�~����;G���W߀Z.��8�}�*��#|U�>C��8i��hZ�U�N
8��c�PR����ykEE?�}�;6 ��f�VW�ƺ+ôM��m�*�{���k�Ĭ�paΰ
�KsP����qJ�P3s�s�F5�B��WS'��vꭂ��Wz�h�ӌb��y��3{����v8���|�+	ǖ��@������Z�#���O�J�>U��Ά������}���,;�y�)��=�z��*�;����vvը����)8F_;������݁O�ٍ�?�Qǲ�%ߴ	�����\�sh�.0�ܦ��v�)W�\��R�t�S&2��a3N�Pb�JS�m���M�Б��4�AW���;���e2�9��ߎ^� $R(�dR#�VN2T`�>_��c�o�ϸ]xk�W='T3�֍�p[�@B�����yؾ4v��1s��Kx�Jo��:�[<d�m�O�d	�ܜ��^�"�?;�bX���m{��o&���*r�EI8�C-#�5֗�4k��z�&��^� ��H�������[͕������w�y�8`LU��cd�5bp)���ҿ;+C���_&��IH�s��'e���� ;-����' @�'<�� eT����t��/H�%�*�j@��z�t��$�U"����˻���(�����as��c,��q���N�����?����B�3
Z7O<�hfʊzդ�(�$�MC�4��n�т<BRu�dD �Lʐ�D]���GӼ�s��?1\���N��-�t��J2�=�A�*^�p��<+Vj(�F_�Ma�B[�ۢh���H��[�](JVr�!� �o��(md|�pɉ�����`h����A�t(Y��r|��j�2��$���*�f�ڷ�r��n�lf�� ���GD~/��51����)WWܘ�8���Ezd?G�U
%�F�k�\��� ]�R�t ��6Y��&���'ݟKk���v�"��B��صe�~�n��~�؟,q����o,�2ЧAkĜ��
��I,��o����§�wK��+��x��3)�;t�N�v\���xʈ�~,YZ�L1N��C${���ɭ�&x7�&ad��ϗ�^M��*�S��|��<��������㬨��ή1h���9�y<���4 {1 ���.�;��{�����ej��eQ}󾔻ʢ(5�e�MT2�̢��\(�p�s�+�aJ�B
��ۏ���v�a�At�-3%d�9������Gɯ��;=՚��5�S��J���D;gC����ܬ6-}>O�f29�#��RDX��;^agz�U�Ye^L�F��;n����v���ѻ�j�������˧�!�%*<�0�����t��.�I&��#����
Y�4�=�VP���]�����o�-| U&#�/ �E6��{3���������zܥ��Mv�(�l��[��̖֨�E:��V���HHFU��x|�����z@N�J0M��t1>�fm�9��3L�n���b���"�h��X�`QNe	q��ƥ����u�큳$��,��m��%�g>�=`ԟf�"�,)�?G8�Ɔ�g��܋�Ci����_r������_ �fp�H�YS��:��%n]z�둤�A �&�9���B�	W��t�������X��L��/Si��:�1��S�j�� �L.þ�([)���b�ڥ6v`(`��>���t�HZ:9#�E�Z���WkY[סE����쥢-53.���e3�R?���%�F���ե���<l��1_X,H$�I���R�� �#U�y�/m��EÏ5%!m�F�P{�&��m�𜿦��:�65��^r��%��b��e�ĥ���p����oz���0��`�������G��5i��Г~�Ӳ �M����S�7�z���~В@l����m���!6����`>���b���m������)d�˹X��~��s���R�Kٽ��K�=��H�18G,���y!8�:��=Y7Hi}��N�f��D&},�5�b���_"�_x@���pF�Mu5�5�����~Ghx�CC̎��ȵܾQg�xb���������ӝ&6~��!�#����x�����l��(�*U�O�oB�O�\�w@�����7o�\U��X;S��O.ZY���َ['Ȑ�q\����@	ل����_��d1A�p~&�(�����y\rb�����y+�4~�����8�/ R>��Oy��G�~�M��H�Ge$B�p9!����G!޽��b�\z��5y"0n�Ct�����V>�c>�e�ō�E�h�'޿��)O�$(�/�h���H%��g!�X#=y��i�^-E�,�����9���y��H�(�q����zro�0mqns�l����j(\�� ���I�����������?$�A&Ыu��x�U�HN:�W�� �.�Z��D2���LƓ~1���bx������̫�e�|�>�X�pp8�]���V�w���I�Q7�f� ��Ȇ��U��K�I������Ԭ-G�,�yOu��^�Jʂ>�8b�.�:���uB��]�g��9���>ܺ�ΗKQŮ]�}���B~]˼��jٶ��M8[���F�MQ)����������2���Wa����]r8�����k�r��:�j*ꫨ#��ch;���������|y���߀��	�x�K^mv��;�K1�r�;g;�H8P&%H-�g���`*�M�x��TEk�se����R��&���k�H�X��^��	��氐GP�»Q�㒽
X[4R!>�C�6�ʉ+�P��:7�ߞ~z�0�/`��;��3A��X i�=N�/#�����`ɢ�q���R.H�Ǥ���{�7Z�?i�Wܨ��j=}���>�B����h��J��ʖ��j��ć}ʥ���tѪ]@�җ����.�����袉��
�uK��}Qƞ(�w��^��Q�,z�K���������q�i�gN�uM�������+�ƩBN"�.���&��,���*��i�MQ�� ���F6�Klv-U���af�>�0a�����~o�� ���+��u���)[�рC�^�F�4؈�ha+���(�1�5�~�j�$���=�!����~�c��?ˮ%���lG��������Xiɚy�y�%W͇�"��r���(�J���< ��Q�*:#4�,itO%�4 �N#�l�"�������q�d#���Zs�Mʘ����R-{����ۄQ4��#H���XZ�'���#p}��0�h���n]�� )d��y�v��r�\@5q5E�/	�
��t彗��xc��l�J,;��}ٴ�6n����VR�z���g���`����ʶjm��RB��y����n�X�+*�.DFF�2y٨�k��Y*�5�.{���ǰ⑌�fmT{�����S��Ĕ�vzG�ˮ�t&l&-���8����dz8�t�8�R	�kb���j��t�h�M�-�����o`)"�iɟ�c��"���[3����B/�B������ڵ�Q�+$JJ�šf	+���W��7�fL��!�����_���zDW����w���3�������53Ot�SIL��?����rc�mܣ�얢aE!�l�㋞Б�f#�
7?$X�l���� ���b������<�)υn�O�$8=�6��~)7��R�d*�M���\Vؗj\�� 3f�9��Uo��=� ��˧�EQ��C�Q�̯�mi���W:��o1� �y/��dp���GB����rnT�v���k��3:��>�dQ��E�4����	���'�Ρ]T�-���gx"F�X�\qF�3�]�T+QL/����ԋ\�Sn��-i����}֨ �a�+�h����,�2o�^³�uA�ώ��h?6uڢ
��`E�F[G��ٛ^gD�T�A�F��5�	�j��^�ΰ�o�k���lN?g������E�8�-e��;�j�D룡�P�o�F��_�>^6�k�c�D���d�7���?��p}�s�g:�;�a�aWa�r��^6�W�9��|�xd_�6��"�Z��Z��(ZI�'�ގ{��������ex���PR�wP܌����i�j �E#�y ��*��O��������k�jê�u�[A�e)�>���Ĩl�		�T�k9��GiWp9�VD�G��*�����et�E,�-���V�\]�^�z��f����P�Ҹn�CsLF��Z��M��YNE-�aF��-����\�9�������K�H����Jr+�7��v����Ø	a0���1���[cڌ� ��_�'+��(c��A����n�c's}�W���B�.�v�eO��e6cI�[4X�1�]N3Y�-o /6��w�I4�=Ƒ����Ha��0À�6,�l�ܯ�5�\���Ò[�.��ѧ'��e�,<q#��u��L��@��^��nK���=ߜ���������z��M�n�:����c��h�����W��g<V����A,l��MN���'.k�5z`��t��kFG`���A<%u�s�	lQ���V����{C�!~�����9:0"-Dg�G��JJ��?���O�`��*��D|��)AQ-�Mi�}ɐH���(Q�{J.�w?��ť��*��2�8�H�%F0��0b��
IA��b�/
�;�ALʹ�R�
���)��qF�������P�v�y��e��u�M{�"u*>�T_iʹA\$q���}� ��*(,�C�'*v9M���SARN���6<�8Z�ΐ Y.RN�-���&c��l{fKQ��ܺ��tí"IՀ���j9�����(���@u3��@=6v��I�\�ך�혷~m�%ǭ�����o۾�"���=5$�c�@:C&0�q��A�²�e�;�X��z����.W����=�^��F�<.��Ed0�����_�Y�E(���%����3ت�����4WRW#�Upk{�o	��z:��k0��a	���Ϣ�KŃ��D��v=n�i�v�~ʅ�v��5 ����@1Y� 굮ps���C�}tO��y�:�v�`���vǃ���g�P��f Q�G��9���V����Û��L!���T��J��x/JUA4��l�b��'n��#��K� �:֠ESRZ���w�$%Gh&f��\�RR�b�tG����*(��$m��?:�F��������� I�Nџ8��2>!u롆��!��B`L+`�培O����!�Ԕ\�q�W��m������W�ST������-`�Gt��b"#i���G�'�i���h��3}�9��\*VK/<jW#��\����=�6$�@�u��_�'oH�hp�0-����#�N6hTlZ�Y~��	ɝ5莕�y�ҵ���%C������O� Z�-�<��0y��,<i�g�#�W��Y�ك�����/�`;��I\�x')�H�@�������X�F�Pϥ�ɫ��uw�T��&��x���YP[�Z�/��	�i�c)�[��C��R$��M�2�u�9.ܐ7�S�9��^�o���<۪UtkSi䱨�ލ0��'{W��&6������Q��A��-�@@���Ԋ�E�� $��K;hQW��7��oG C<V�);G�2�V�u�@���c�j�,͔��PJ�jk���r7�qдR͜�����MD���K��7l��@l��)D$�=�w9�=A������5�,��+4H��6�z~�69k�(�A	32��߮W�z�N�����T�B,Y����oSή�����٦�N���Z��\���8����.P5�����p:��Z�ꫳ�cyS.������� Y�;-М�v����ub.�БR~\}���qY�T8�\����9�]��#���l��Mb�ˌQ��,D?΃JQ��0EjN�eH�VT� X�����j�:$�,̻���By�[^�o�
�;�N���P��%|�43f�&L���(aʰ�p4���؝0[�:���0��g�R^����f������y��֐}�2p�'{tx^rL����G]>QM��v~o��6��wnA�a���m�
�4qMk����G5iA�E�)��\��/Y�H#0���㉱��̜�N��'n;^]	�&,�Y��^�ﱊab
C��&ш�ؑ�'���K����/�������x���(�vF��Z�i�%k������}�M�<�L�1V�Vz�A�j����v6�=��yG�ˮG�������CN2���*L��Q���[?�˧��Eg���7�6R>�6�b��ɪ���p�����s�O��GR�����(�3,�N!K�lI���O�A'������On�|��#S�䯇�K��Ao��f�����9ҷ���d��ܰе�rܸrBz�o����)@�T����a w�>'TT#u5; �<!ǈ�:!J]L��ūQ(�n�V������;{��SV��g��?MVA�sw� ܚ� �7���$6j5)�J�J���(L��z&?��m9 A���X���z]J@\�{k�Զ*�e��V�L��`�4@t��������f��-+�����	&d1 
u(���ʔ�O��2��m Sml*�Q��
�
�j=FD/�!�A]Z)��?z��u͇N�_cW����2�ѽqb�H���G�{ŕ9aԛ��cf��,T�P�0�0=��{E�Gk����5�$i���Z�宝�����S��N���T �֜� i2�d�>pǵc�@ĉX"���t��I���ؕ��h8��5�$�����/���5Jďr�@da�B���v�˓ʎ�d�Q�#� T��2D9A�����"i��ʷ���ܥ��>�q�?7����8}�$��t]��.U�]E��23�\������0�Vp�zI(誻��>vM9¨(�?�B�j��}"��V��x幨�Shn�ؾ㑱��?Ν�@Q��6E,܍��)w�B[��@vy��پO;yω�_��ux�� ��ĉ��k	֐��Du�*S!@2V'�ɮ䴥����?
=�Z �y w�²���Ss�/��`(�n����O֭�8�\µ�%qi�D@h��o�����S��A���� i�,�g�x;�ɬݗ���{k��H��(�	4��$��R�Qn�#��F�3@E|�RC�"Y�RԤ�\,"�z9!���\��d�'T��N:+; 
��s��ȕ`1��Jf�������,�n�o��%�����T�\����?�_�`HD��L�g_ޗ���9L=D��XPo�e솂�0(�������XlUJ}����ҷ.~��0���6y�e���/ �Y_�l4��ѩDq���mM���-�Gr�pa�M�^��o¸���~���m���<;0�U��%L�J�����H��f���m#~9���Mbv�c�J�P��2��+2F{��/��aS��>- ˈE�f A��2�?*��s���| c_�Tm�'k���i5`��mqf!��Q��؛�A<��"b*�4�>D@5F ����"F䚼$��gR�I����ʦ�|��?�~g�=��G���G��ʤӦ&��z�hJR�%vp�QR@���M8�H�L���ٕ�%ˍ8%��=���+�uK|�8Gz���l�+��"��`3� ?���#M���ޝj�q�	g�6��Bu��I�jY�>O�h�n?s	�2���&&����@�~�9Rd>�f)@ҝ��Y�ď�#L J�Y�D�.������z�#:mP�f'z��������^�r =�0� hU��S�9����⡝�׆�q�H��r�1%E\��aa
��P�S��2'���v�-�����Z�-�+�H����K�r0\�c�\��@ȑ�e�"�W=�?��NSk���-�=V�v�I�2�FpҜ@���k˕�F��*�R�1t���J����3�QՐM��rѾ��^4��+~�/����ruþno3�T8&5���*Z���{��|���,��K�ߟ �&�#��o��j�w�w�@�@OZ�z<�}�o�A��/>��(��z�NB�j5ז����o� !�l�����Jq���'{gp� �I�H�tc���c�9�&@�?�jF�U��-Q��v�] ��.�K��ݓX�&��ds��wu"�����kJQx��󛫠���o�K����L�hɑG�Rj�]����h
�0�x��Wڧ�����������*2��ߺAσw��ix^w�F�0U�P[�c,I��!��uG�z"��1�_;pgM a|2SZmǫ��j�͠y���!6������&�medy�W��]�ލ����?�}
��V1���g͸gK ,�4�����h4�j헜*���4W�g�v�RO4�Vt������k��2�^�Y�4�����wwp,ث�[ M`w.|�� �d��Ǧ8��M�^z��S�+ג.�u�Se4;�f:"xӕ\tB�v�4m|nbaM����$+�s��� b�@�9���]F�p��~�؞\������vv�U1��������V���
P�)KCk��b�{"�n� 7��H7B;/ ߓ���D��٦�#ļ���T\F�Mm�Vh�5!;mz�� .���9_�v�G��ƞpP�����²��G�v����!�������f�>��0��pX�5>��B;���NLv�|$!,����3h.��tR������IC�� ��VS�d�9W�$�5��z�N�%�����&r��<�����K�/�����'U[�rr���O`�l�Y�ս;��<��I!>�8�_�?�V�!����n��ZxD!T�Q���gM#Z�`c�]�;;��Y�Q��p���6�c��S=E���#?*)k�Z���Q�뉓���(���O�d=�<[�9�Ї�K�QC2��֒�O7�M�2�Uu�V@eaѱ�N#���W���R���<�U������a.\���	�R!QL%�����59oD�0���/^��x}�ų�Gwm[����qfJ���ʤ}�d�g�P��n�Ġ�̦��|����8�a/ν�T,��t'��ڢ\��
| ���/G���2`��������AB����y��n���3�,������6}��:V�%a̾q��m[q�=�_�k���sc��I�]V���`	m
_���H1�Y5�TＶ�d<��\�c��Jg1��W��g5�te��'����]lPf�w�O� ܷ�m�P�-U�Ot�{'���@�xZ��.b�~H�h��ENɇ���l�0����t���DI(S9��l�>�u�>왓%*�r|ĉ�Ew��¼!��)T��l�;EeXH�7}�Qe�:'������H%n[�z�H��o�#���*[�6�����%�Zh5o�f���� Wu8l�T~��Ĳ�s(r�����I1&q�/��
W�(ސ����2+H7 �V ������FFA�Xϟ�M��f)��U^:��f
�YIO/��� Uy�Ɍ`O#)d�(8zufP�^���N6�|F���M)Phf?�9���rx�+VF!ܴ�g����z�������<�Z�Pe*�H셐��f��R�@��� ���Lq�y5���>A}�'��(�f��4ɔ��{�z>���d$b(6��-�f���n�#��:�N�>�K|���pX��7q�1d�buR��^�K(� 9��[������/�(N��\͑�&bdElaw�5/���Ul���w��rτ��k��c~�*��'1p_��1z�٥/k& �'�s�LH��K��pN�4����T4|������"�����w�ۘ�(x=AQ� ����	<��r�J�^��J)��(�%�/���п\��ls�:u��O&v�߻�GT7��
�� 6���*"p�tT(���)�A
P'# K��@/OUK����B�DOQ��""��g󇠐!���I^��)��/�v�� f���-�^ϑ�A�Z�X}��_sB�w����H^�'(�x{�w�i�:!ic9�T��L�އ���`'%a�@����9�ޛV����L~���O�b�?["n����*$P���?�Lit_�����H��p��H7�<�%�2�nî��G;.}���u���BA�QY�lޘ���If:�9⋷�� ��}F�
�U=E�kQ~�Q���M��R�`͙e�Z|�9�&%wM⪞���d>���lA'٧�Q�D��3S¶G�^.��v�����ф��͍n�ڿ$��C��X%E�����X6�����[ϸ.A�R��������S��"�9FK���`dǠ��a��+'o��a�'�A��`�n��RF�@뚜�f�2C�E4�ﺠu4ضޫ���Vcc��+�5��M��M �sti�w�7ͯ�y� d�&��ŚX�� <��E�I��h�ƃ���B}����
�9�^/]Qm�*8l��T�ک�ϰ����:H��۶
Ha����C����1$2zdVT����'��<0;��m������oڅ'�M�1�S��w��\́}���,iGP3�4�'��X�N��/�P5p��f~y�2ogL�e,�Z`�#cg��)��g"J'�}�ߗ���iYx1������#1�[k]v,�bq|��k`K��'t�o ���z|��]�:�.����b�$*A�M��.M˴��x�[����KaܘI��ZL�D��0���������tη�˦�T��W����S��ݭ��K²�^D��Di��F����슁��c3� �2aX_oG��?���t���7Lr�/&�V�/�"å�lT��a3T�
��IO�M�����t) �E0�,���Rֶ�}��>:�\�`�y �7��8����m������Q�j84
d������{Qd���w��*�Z�1�H��Fv��a4b��b�҂0�שa�7 OQ�'�@[Ea�J�X�ˋM��R��٨�N��l��u�9z7�>���@q��O�'�E(m��;k����h�ުP�l�l �Or*���\ɮy�<j]w���B��X���?���DL��g� U
��d�\O�2�d����--��?��.��d}��u�<Z�~�#�����"d�{t�;��c��4�{ѹ^��ٴ�R�XPW	_q�&m�2`�O��d=���5m8�VqͅWW���8~�*%�h�K�v��b��Ou�hP���"��\��(���H�)3��t,EYR�*Xk�6=�P�ףN3� n�"*3z��_�!	�5�`�(��5S~t������Ѽ_g̢'���M��BJ���g���=�kC����Vj�ǽ��r��|ʰ!U�6��s���u�<��Qޜ\�K|&}�Dps�3*�n!1C�[�Xv�2=LX��*,583Nk6�E8c̵0��E�+�$��ب��dv��&��ЃQ愉2M��O��Pm˚6�GЯ�34;*Q��(�B� M�+�e-��t-�L��{���Z骀�̲O#�1����L4��҉p�D)k�-P��Â�[z�<����TϞ����b����r� b�T�_C�X�-�����ע��p���������w38`�#b�7�i�pok�|�%I>�S<]��B�o��*�uE�!A�+R�݀��|��:�Ux<�֐>|��Q�['w��	'$ɵ�_�0�0����.��1��	�	�K>��v\�k��$u�m�3��0U�	D�sR):A�9�Sm�Ӂ�7�Y(�̕>!�9']���T�;���e7�)�[).]A����pۼk�˲|���	�W,�Ǡ��"]��{�C�(	�H��^dofX��
��ӂ/`0�w�#�jcf?�&D��28E��-����0��w��Z�F������s�{}s����5�>�$K�ؙ!�j[�#�3�($N�s=f�:�>�#aO�s�3K��}]#d(�x;���A�P�)x�I{k�)�f#0�0��m6 �{�c4+z��"�(�}܀b����ck�܅�]����$�H��Όh�
�w�I146@���b�{��c�V�T��
��O)�RR�KHo��j����n|��vET�7�~K4h�3�7&��%�� ��/��
4M��s�s�#+��T5�⟘4wB==�]�c�J�d{l�z#�'X��Q��s�F�,r�Յ�/9��~�t���r>])�����ދn�<�JZ�&ݮ��x�_�|�����_F�`Yq��Qє.���o�pO_���Ly@��������=t�L!otr���ٟ5rQ��ZwN�J�/�����H�_M�YA��>��_��>4��ns~�����T�` ���ԇ@�]H��]6lHj�/�p��	d`vw���Kj�ey	����
��y*s��u�ue��_t,�Te�Ht/���9��q��Bʄ}W�Iѐ� �.a�����li�}�@���,8���snq2���b|#�|��6~�(b�u����h0�~!t�C�Q�'#�9߷��qɾEPd���a)�K8�6=Z��� ��p�ɝ��[���˭!^*{G�N�E<Z9��������*�8`�����*�b6�h����$M�;o|�DHK�TY)�Ţ3���԰:}�Y��%D�H��t�h|V��Mn� �\O�dw�PK��1�'������P(aǧ���C#�6�@S�k��y�␷�g�,�{�`/̓���[fƖ`��"
Y��o̧��~���P^�򓼵�� ��vh�i���1:��ж&	�n���m�2/d$u�?�����3�>�C�o�r��I`*�*ݶ��:��x�z1q�iǽ�4��PM�#��w��.��������QHӨ��O%���7�?w!O.�kT7�5���&oI?�n�xM(l�t�b�%(T��
��v$�R���0R}]i~���vr/�������0��SP� �O�Q�9T{�گa��t|2)��{K��'�&�;\��+���.�L6 ��e�oH�ZQ�IV{�����B=*�=��ҍ �j��\�9���7O�c^W@���ix����FL�}�����]�^����lC��� �+�&���~:���);ZxTr%H?�	~���k$�BF�;f�f���*�IT��p����䢄�	�n�(MT~><�̀du%;�&aT��QJ�s���J#j�X�.I�4��4�X@�	�oV��\��9�Q�X�{a��L|J��]f���������Ӷ��24�Ů��z�o��o����6����-���̆��Sj�1�7�2)���BޝӢ���e�f�M�����{�R�^c�ķl��2u���Ҁ	a���ě�AQto���l؜�����h���tϬ,��ZާG�H��Բ�FI���)q����)��Y+Y�v��*~����v�\|��3���&h�۸l��z�!_��N2\�ׅ�5�!���r5��i"�r]��w[>���A� z��MZ����?Ʒ�lU��<U{g�&\ȍ��Sc0�����F(
��K湞a��CAn�|�Æ4]�( ��]!��~ָ��F!� ޡ����_������0��W�7	�~�@�U�������n�肔�ZJ�f��j�y�.d��㈻ա;��`ٕ��j-��@U\��|^�em������ߎ$<��4_����MzS�w42Q0����U��ǯ��/�$ǥ%Z��7�/Ee0p;��~;Y���iUL��B�s����8�vU������q�2�4O���'�τp+���)X�TӒ WB ��8�לs��?�鴹^�4p��U�?�T�b��.Ax���|i]	'Tςu��6��O"�]M�݅���� "qՀ�ЁN �U�<���Vƞ�9�̊���fg��9U�Ԇ=1w�ݮ�Q͈�I��s����rAC���K��3��r����~�m��|�a���(.l�W���o��!������ �J���3U�h�`�.�'7�w�vm솾�
��;�Ȧ��$,��F��%��F+(��i�!��m���[B�	�3�=W��Ơ��F�/����Y,R'�h->�+0
�&
��HQf�E(�C#2��Sbo 85�?�P�9�lR*�ڨ9r^=Q�T%��:�Z+>���+S����Bn��]F�l��q�R?A��T8�1A��-d"��i�|IY��-0Q��P2��� yՈ0p��PYqQ��>�6N+tb%P�k�?������� ��d;��Np''Q�r�@�p��-�N���aKQ?_�_�NX���6�l��8_נ��& �d%����R�U���Ԍ0[�Hn0ɹGq�TO���,�:W��y��sq|ܫ{��N�=2�6����Rn�;��l|s���WOD,_WL#C��F�7����ڌ�Z����u���R� �ú�4:���c���R��&�n�� �>���NF:�<'��j������^�a�dx��z��38Z<����b0�٣�z�0'E��6���:�CH��?<S *��fT�4\֪�_����F��m�?������QREM6C�:?�=�"~�`�7;J��B#��z-jg*7�G��Q�"�ꉂ��]U�a�y���u�=W�\K��k�f�II��C��J'Cw��8��*&u��QM�g,��b�D���$���R7�E�T�)87j��cX�����:F6��|#e��7�}tq="�p��l"z$�0�F2YjW���[��D��;Ҵ/�]�3]^8ۢ�^��X4!�u�|z����b�٫���^�q6<�7�dH�&��q�t1`U�}�G� �XК�1�		T%���X�;ՇG�[�)����/�9v4,�9�/Ε���3e2"���En�mE���3l|�cX����+A�WG$�)��ڭ(u.��s��Z.���s��e�9�q�(�MMCn�.�6��֊)�A6r�q߇� �@0 �T�a�s��.EM)���WD4Yr����D��+<ϫco��k����M��'�V�ʃ���K�Հ*���������%� T��)�m'�4_�,=M�$�Lr��xU2L� �Di�#R�����ց�.\�U���R��I
���F�n;��<p����|�_�F��:��IUf,��V�h��`7�W�N�4u�,���y�и 	ѣ�^y�� ��GÇ��f�JZU3h�S��&�	����E٫��� TP:�y�[�4Q�s��]>odp�8!:H��Z���k}:)F�3�f�y�J>�(q*��kj �xj��V$����]H]��|a����>��7v�� �z_�呲��\&����3ݦÿ����LQ�l����o4n�t�ab���3��������r��(+���لC�ަO��َP��s�������yEp5��?˫w���Pq���?��(��1�Ǘ��Evr����(��n���v�q��Fk�
K�0���>%�y(�˄:�yYi�7Fy���8N'֍� WI��V!��u���mxp����������Zn��=LB�m�җ��O��w��o��$v�Z��7u�e�b��c�j�#-�a琨�����r�.�cr��U��_�j� ���� �$�l�q����������$���xö$��s+e*p%*�|�N�&�V�m���)+=L�ݜ
�Lf4#�� �6~���$y��m��a����bX��C�b�bF>h�hs�^UQH�T"A�1��m��p�������|�c�tn)(�	�L����W)��n�Dt�������U���x~c����"������N6�����U��K��8S�� �-ʲ�;<�m���ڃ������o�/Neߒ�U鈑�d�
t㩅�t�#{#C�mC�V�� 8K�����]GiN����ﯜ�^����cX��>�/a�*{��𵀄$�֦�X���}���r%�<����*4X{%��$�]�DS��O`D�ׄ~rk�|GY{�\^V�G2�[����,�I(��$ޢqIވ���Zƃ/R�/=�|r�m/���+��|[4Hp��C���c����"��2m��K�[_m�ޠ��m���J�K ]�x�蓰�DyC����e4C��8��2#+	(g���N@�)�I�,�l���l�DKb�p�O��%�mO
3��>��^a[��DٱU��8�� �h�-e�5��T��/5i���F��R��7��G!�N�(��'5�!N�"y5iP	:B+���Z]zV��_����4�O��p����
�t��-����LR���mnqe�\�֎0g��F�v/��傎s2�����߫�(G��N��y�ЦPyh	�抝����(����3}�#X\��-!/�^8W��?����A���ܿL��/�ڵ5�e�p�6����\�We�#�<y�U�����J���yFR9H���w� �0�.���w@gg���BiZ�:4�
R@����	����*#�Lsф���|v!��h�êӛQ�6Ag�`�G��/�H��m��I��״_J4���Ќ�02W�Y�/�va���"~|O��a�[�cQ��BI�U��0AELı�rgZ��p��t}��).�C��e�&5u�yD���l�*�Z\�U���&G��^Z���� �;�{�2>I�-�Z�<�*2P�-�}�>OH�a�>��~�� �L����#�&9�|�Z]�� ��e�)��3(6�JJ��&���t�!�}�ϩ�d�u��6�xiX3��9�<Z�2�0���k��z^��� ͓R��I4k�z�}�+}�'�4����#� !��,,hο�����9�-5>��Rio�����7Bu1��R��
h��|L�u�͘�*������ӷȄD�^���t��ڈ�/!��1��LO#)тб�j�e�O�V��� ���R�w�TN�_���)�Z�)����kο�j�]bZ�zR�9A_�B�Rڤ�����l�����N �9�M�iz{1�5u�.�z�v�V�0�Ȧ�_4�K�&Ԉ�g�H�*��*�N5�_j�{[�nE��� nA#$��X�����)��d��G��܃ހo�
/0���s���6�g�:�JSB�q�#{Ac�=�V����d��񷡲�;��5��+�]M��eզ�h�P����C�hc�.�1μ�����2r���}(N�.A�����eF_p� ��~z)�CǄڡ��o���ၺ��3~XE��
1]��_2}X�	�z�G����P��p�2"0�'�F���/�8�(�N8�銢��U-6ض3�9.
�l��a{�K�Ռ�����]��
���.)ޝ�6��D�4��2�&���&�}��P������(ϟӌ��* |��݄H��M�9��淯�A����(P���X�5mʹ-Vf3$̅"[]ےRwR�`h���e��~ת���������L�i4��'BoK�yn��hd<�v:�ޣD����T"q`�wj�}��`�����r�"Yb��E�&]�{��\�����2�s��P���I���Y�m�1��]�Z"�b�h*Q'q6�ab����2�d���'D�ɂt�~�_ry�
�9��:�"��#8ՋpJ2|gJv��,<��Ē/�}�����X:�6��Q�eS��86ӜF��Mj�P��e j�ցX}ng{�7l^#�x��r��"�jЉmB/���A\|�n�����*NHL�v,��
�X�v�/�E��\�X-�{W)�zFo��4�q1;K��B9�FB�fm`ֹ{�
�a���'�я#Y顔�>��e� �D��%'�^e\?�����cd6�"f��<����\����>�����i2�Ż�l�ɝ���*�o���>O�8��F�_7����܅ym��(!h6��4.zP(+Hc���S�is"��&�1�ŭ@K>��e�
���Q�=��eU��tяq�`diS���|\fͯ����aC#+}������[���w�_��Q�a؍�+za��NYG��/κS�����G�FDB'�dh4�7�Q10������ �c%E]�#��OB>祉���;����F81
�"wi�Ï�h�e?9�t����X+������˩��l&������§����n^�u^��O��ǻ��;��mβEԶ�VP��#˹*-�uC$?@p�t~$��� �G`!�':݀{�Rc�i�Y)]3�w�2�#d�n� e��Ʒ 8@�@q�?��x��ȡL��·�[���ʟ|��|쭠ݲ�hb�*v%�[Bɷ���F[�p�(B�葙d�qۣ��'�e]����m��&r�������hG�iN����}NE ��t�Ň�uo?�}D�\V)B���������P17���Hx<�@"/4V��AS����l��8Pک�Z"�r(�_�آ��j�Vy��)Jeo�pYH4ֆ4�~2���(B���xR��� ���y�$���������/Ε䋦�F�]\���C)$Kuw���EZ_��Vr�Z�\�AM��#b.C&EU�v�d1�y7E~/-w������q��70Ė�0<���;[��s�
�6�L�AAvov���/-	��c��ٕ+�
!��F�� �Ӻ��3���v�iPI�;�J�����:��ћ��t|��m����3�+�Llnc�:ދ�"��R��"�A����O�ؕ��������Ab�B4i�*3/��ࡓ0��Ɇ��R0KX�eSW%�!�ou��̼ȅ(+��7�-�TLEo�"]��s��]��2fMv�Ζ�w_���/�&��K��g�0�����)zy'�..h��ŭ�G%�v����HeI���F�M�o���v'M�Մ%�Kҕ�wd�r�P��p����H��9XSy��01D*�;�"Bv�9������x=0�a���A~N�ԛ۫�ÊM��<�o;�����i}��<�%��Nt&��_�j�y�Xlִ�,pE;y�����q�ʀ)Y��-�m����fѳZ�'��W��&8�IR�}F�L�kۗ�w���ôe�ؔ�n��A���q���ꛈ<V�:��s��x���hq M��g:r���oF�/�	Ar&u�O���z�O4l���Հ��XJ��)읭���( %�wJ���q�+~�J�(�o����=�,\��i�y`ϭ�L����`\NDm�qRȖB�ߊd�B+��C�ǉ�90��/�|�i�&x�d����u��@ZToF�`mVv>����2�?ԪO��yh�Ka՗���>�<}nV<	"��Tf����]���oK��b��`��z����U.���=c���lX�/â��菂ې4Ũ�֝��'��#Z��Lh��*�J\��8�o}$�uz��N�-�P.��Cj0���� ��Dۈ�q}.��ѫ���'"�6��ٹY�Ԯ�r���U,J/�6YA�	�cⴣ�x�����\ЩK����^��vi-7��-<� ��u�����XQ�)�]`�
o��k�3��Y�������g�:���O\��D\����>QO{<ǆ�d���A�|�O�`\
�8t����pz7���Y���8%��-�V�㵥������4���'���T�<��Ӥ����/`oG�ig3N�X`���
mE�Q��1
0��[�,cБa\�"��ߥ'�C0e�|����A����@��(Fu��jAE�֌��QLK�]Fc�+%�`P�Z�?��(��d_F����!�@�VS^��b�2Ȁ҅���y��)�CuN��L��I���~`B�؈�^�<��V��Y
KRN�~y.�0�h���h^�3���O��O�Eߎ�O����1��$�7�hݍw�:��%i����-]ʯ��=����PѲ3nba�UG�z G?�7rv�8����n�}�/�JO�l�m7<0�ގ�Ef�W ���7@�ܺ�nG,S������B�8���^A��uVf	�xaZ��@ٶ�lf+ג���6|67Zߡr��!���ׯ�m��Ew���t��f�q��^/fw�#XA��m?Ȱ�ѫ�-I�.E���0�\������{X�)�iz�!����?���6X�&��j�<�ƀ z�W�����p���3交<�4���U0�'�.]�;/��Ҝ�d�(�w�DoP_3����IᗙkO{a`$t�U~�ذ�2��i���^�%�M��/
S���	_</���{�Q���Y���a�!���/�ĭG&>���6�{�Rx�D�:����y�/ɘ�1�L�vLe�(��z��?jC���v!d\@G�>�2��Z���v�(�r�޳��6���w���#]�0��!�Y�=W�#P׍M@�JA�]��E`@��#�*:���^�bI���t��s��BSs�.8t(�gU���ϗ=��:ŵ�ֹ�>���ٖi�^������]�?Dġ\�{i\���Pe�Y]��sAQ*�W�@fޭ�qt���u��/��Y6���4|�i���%C�F���L^O4gң�/�.U�te*`����l��H���h�3��Q�e��r�8uA�����.����*�\�Q9)����#��D�8H�o��i����S���
\`����ux�=�MݤgU�������q����U��?���)�k�Q�� ��'�r�ndR �qP*(��5�!H�0i��#1y���G��)D:=�U���R0�j�����I��BӠ�T��I=��r ��\���i��?`��ႄ��P�_�2��Vz��5��p1Q5�;7���7�M����ӷ���<���aCU�U����d�������?��I�*(m~`TS,��@��Z���aZ���s���R�c`(��qCF�C �L�[��m�̸��z=h��O��v`�Gm�)[:W��Ab�,��,��)%'U��K��g5��u����R���1��H�\OR��+�����4,ѧ2��ݺC� ����GO�`+���;��H�y
��O�Ȱp�h��68[�D����AL�OQ�+	���osK9�c�hF����L�������?0!W~}D��OI����um�b�Rˡ�ej|;MrS��`����jQ���
����() �؊45z����w!��N�oۿ<�q�_)#��D��1��ǡ�_Ў�9bK8��6c=NORYC��x2���yWω� ����@�꼩�K�5�v$�PNq�RX�������$m%Ʋ����C#��4B$�sVw�0��z�e{6�1>����M����sQj�Ǜ��q��*����c��̋0%�M�hoMr���֌��v�t8�m�u(^�޳��:�Ԫn?�8˦!؜���	d���������bb���nO��7�njY4q��o}�(��:_�h^�=��K������}\ۓ��8��|%��u��O��Bo��9A1�j}
+S>b�,�3g+�h���b@n5E���\�w��,���0�����%Kk�x�m���Y09q��	$P[�9�?&x?1r��~��Ǚ��s�ZE�m˨����D���P�ﺫb%_*?�mȇr�R�ކ2��'��^��L!�0�KV�`��"i�ƽ�������].�^��o�����E!@}��>�4F���̞����Bh����
ĥIQ�~&�>%��!g18�T`R����!�5b~�4��Sj��g#�\���+���aE&��Cւ�(5��k�ʾn����n�ӵ�'��3�)'�ýbZ����`X�)=B�|�!��{����#�q��� �H�S��!����S���� ?��s�W�(@M��3L���'1X3v �f5"zCcJ��Ѵ���ކ�Ʋ�o�<���|���E�צ�ɡ��W�ω���4�͎1��>����@tA�5��Tq�r�`\8��%�m�s�!���zC���8��V<��6]���/rl'����B�4�6��2��x��bO[4Z��|>�uY�c�#���S�x������y�Jt�\�Ѻ�z��LN�m���ܠ&��Ũ�,I�k�������T���d��l�K��E�ku�L�q4x��JG�y��>{��ྜb�1��M��/��@x>��ע��1����cn���0���iە��j�Gn���i�[ʶ4i���)�x��=�N<�jŊ��^����Ye��\2��2�ٔ�#w�ZQjn������������S~�&��F�"���@��/�NN��s�n���R{A���!�#���x�qCS�CG��C���H��Q^�o�<o��^ȵř���^;^�I�Y�J
���K�ɼ��F��I�Ǎ�O�.MF�[~i���+NI��>�~�����W<�>s˿�nd�m���d �ܢ��/�{�ڂ�[_��`ÈRh�
vI6e�
6�wG�&��pĹ���{���$�u�cSԄܓ	^�-��>ב{o�C�	�{���l��E=���7��M����w�׀��s�>^tjr�Ec�A,���^Q���C{��!�"A���� p��f��X�.��m�4����G�N]��ux���
O�^W�XTj��wО�D$A^~8��¸�`�^o.O;�ۚ7yhi��:�7x�i�;'�wrw������MY�؟����:��WH�pW+���~$�҇���]e�뢐���A><��5UqYђ��w�=��F��|�`&�
P�q�]�:���A��]젍�4qTs��j��9w\dV�*��><ph��U�"�*���ܢ��'����i��F���Ww*�PΏs"�I�&?I�?D������
�e�#rt�sպmR��w�/l:���z�x#:��	H�!O(]͑�����M��PP]��J��g��@$\}�E��0�Yn� |�`v�^:ȣ*�IЯ��JV�����h1;�QgD9����}���f�k6�p>��'(�mlH�j�0�O c����یG�����q3�>�|��t^��e!�ߍҁ���d&�Q�
�(����qе���w.�+0�"����SVäR�_J�+��� �2��	�sp���T���Ь
Q�� �}-��f�o�"
p(Kʕۭ�;Y�ӫf�m���@*G�1�Ù�D��ߊ3J� ���K1�$�nO�\6�fo�:�KC��@�sk���ЭBJӍ8Zy���r��ţ9�*>�]������n��V憿׺����z&���2��n���$���E&kT�.6�f\Tw>�=�6�ϧpV)��d�WjO��E�W���}5��ٷoE�,���ӬZ�!MA����@ӫ��۳��V�v�ĈG����^��ɻq�2r`�x�T�������JʐO7!�d]��my�fw�ak\ء�jj����tK�����W���$0 �.�k}�GggV�`a�U�C�VRN�U��;K>���[Q~�ۥ����0�����vk�ə�Ft��t�u�x�"�7�8�9��<��Q�|���5�aP����� �),c[���X���0Ǔ�-f��:cϭ��[`0`^�X:9ѷw���3AS;���H�e�P'�ܨ%m�@yR�/�ncDr�G(-�s��`�] LI���И�3�����^���MӝA���R���֯A���� Y��y;$�̈�����+��	&����ȜIQ�}�<�|n)��$��g��[��m���6�W�_C�o�[r]�2�kS7���$*�����Tԡ�B��+<�T��V�T�=,�wb� A"j���]�����Wz���&�[!߭^0�I��;-���~�+B�[c,�Z:2�����>���Xx��YHFyO��)�X^�U��us!�P��p�@�<��F��\��HY�ϫG���,�-���ʉ��}W3O��ނ5fv�Y���)9!'� @M{в�7�A"+�o�5�@�P-��=��OkX#˺�2s�j}`ȣ|��EL����Qݞ
��AI��o��Ӑ�~� ���и��o�Wg��".L�i�M���yhZ
1Y)����K��wd�V�=3�m�����������U���LM8�ݛ*�S ���P�ƹ�j�]`O8R���|�\X�|G!>�	��ߔw���o�A����Z�X�6 I�������쎰pV�mc�$3o���v�@�X`6��]��ܒ�.m�}'��5L)�bT!�7����|JfMd�'
92nՔ~Z1�U��KwWk�'���5�n/�|�Qk]����;�@ �ۮM'�T�)��8�& o�%kܛF��5M�!}���8h�Z�ڶ����Ĝ�ס�UXÞ����z�[)�m�Z��ۖU �GHB��i/�d�4�LW�F���Yĵ�	�5�t���O��z6���/��d|TQ梣�뾵���?�r$_!B��Dv��仿ߐ�C�:5΍E\�E�h$l2���t�݂ ��NT)��b����e�v�J�N�T�Z9������[�!�E�`ڿ�-{n�	ꎁ\���) �����d�de6��g�n��U��[E�mPL*�6|[P\���zEi?�p���OX��$��?Hf������"fW�Xdq�8������f�UC,X��M�}�r���w�K')�ֻ?�h�5ÖF�'!����Y�V���wk�Е)Bd����{��D4��a(�p��"qW�'Z���H5N�V�>N��w��FG��T7��;/�������3m�b��b��f�-��'ނ����_ŹK��1��EE���Y��t�������K�$�o&o�����i�R��.�c"�p���&?<����z�K| ��r.��r�ϛ,1~����%�v+k!�F}|��e�4(���h�'P\�zg�&�'�&W������*��u���*�R���ɇG$�ޝ��M+����ŷ洑A�p)�G�!*�F�0�%�9�W�t�6��`#>�s�䃖��?��F��ٚ]t�.D�^&��@�j�k��Ht߃����L6�v�(s�J�-�k��a#6��4����p�+2d�*�h�h�,v-��a�j}hq �M��̵G�"?%fk4���z�;�O�&���]�;�V���,x��(T�I,z2����?Ӕ����.k�����3�6-!���ZU��3t�f��L�$&Ay�D�Rz#�Ő����Ga�F�	eI�$�����,�[<��j�!3p%=ī�%a�{F2��=�}c�SV��Ѯ�{�S1���*�Y�S"
I���lB�� Q��#d�0���MU��V��cl�k� ҁj������2VHd�]| ������5��x�ÍD��G��_����ai�G5��箎A��5I�������@�cƜ�킯�y](����<�5͕�`H_ՙ����-R�kC:qm���L�ˣ���@*�4�z��i.�q�S@�r o�a� �Q�]�Cb�o6 }_�� 	��8���!�Lm��g����NZ�����7'ʴ"��3/t��t�eĨ���q�F��'i���,�a$5�F����,�1l�Ѓ��J�D�d-�8*�����є���@;������s�'aع_��_�G�VM�Z	���L��2-���G�il�ؼ��T/����7�H�8@ԃyѯ曄��z>#Y��Zw�W�~�ٳ��)i/�J����R���ļyb�g����]�}��� �~�g��MbXk'uW��(_ ��J�4q��i�n�٥N��	lc�fE���a�<&8YGFʨ�Z�3�̳����o�S�Y�GF�D7������l��2!���\Vu�i,�Ǟ�Ѿ�\������2��mEmKS���<�UK�ɋ���d8��J��iD]�t�f|���I�����~b":|�,�L�)��x+�I󙖞6 Ò�/~1��ܭ��־�WʟTt ���è��um���p��V	�n���s��&L.��eIA�قg{;�SE}~���i�����/�sl�#0�,�Q=����^* 1�����yP1���Ȇ�X�K�؈BH-]W��WV��W�2�x���f���V7!Ƭ�y����b`��n�O�ㄙ�^����%3'������Md��\ռ�ҪRC�����/%O���X������06[��Q\��D�x�y��&�[4\���!Ͱٳ���������/�MAhO�m�U"3����N�O��r��HS6�c���/U]�Ytp~��.�;a�tj�>�kެ~.��N���5ze`���R�h���׶�ԓ�[
pf��D�)�Y�~�B4dmD�c�����G.a	��1a�c�#�������ǒX2��E�e�'	�dzz�|MQ���ݸ�u�ق�� 9_�j�\��������;[��E��9�)eF�Z0���IM#i�z�%�f7vm_e�l`�U���wׯ)�mdG�/_��d/\2�&��M�>'Ҏ=�qTf  �LT��L8H<�!��ڐE׉�O����n�P�a��t3���_)+�Q-<��.{��UZ�z������+W.0�K��p9\¯�� m�-�/��7�+�E۱�!?�����y0kI�ڧ��j����{����qP;h��	g xp�.>˚n�l�ߒ�D(���8S> ��0?�;R�#��� ���@�c(l�g�?��� (k�W'x������)>I\�K>h�''Z2�o���ܽ�5�4_��HK�H�w[I	s�tL���[ɓ7�$I�w�T���ײ�a[JF-�߃5��Ԯ-��\��Sm��o`�|�8��D�O��$W�����%\y�O�o�Q|j15(��0#C� D�E$�7���A���^S3:�w�,��Y8��;@*aK1ݍ�"���6;Z��kq	�d��CO�	����ã�5#���L- n�;�x^��<.�DA�r��"&���&�j�;\n`�5b��@���� |�����_;ޘ������td�lU	�侓��Y�O	J���P8{H?���B#��_
���bZ����⎳DsK�`Ŧ�}кKd�7 \�x�g��������I��h?���-��
��DMAA�:Q�+g,������j:�Ń~��j��存	k�%Sr��߻��v�ʸ�\z.<��r���t���Cu�
�9=�~R�b��'?��8~���ï1�:�;��|�����η���MF)|[��S�� e�X`, ���v�#9��.���W ��
 �)8���s�("�Ȇ����`n*������30KdUl�N�p�U�i��R�I`�z)0O{��sA��f��H�8Rm)R��%RG��
�mm&Ȳ~W��c�p0�h������������2�H�aS|7�,wD��)"�ֻ�Gkl\����K�qH�%L�!�$�Q�R��B�C�bU-��z����
�A�u��.)����gn�/ d.h���Nm���j����Nগ�ӌ~.Dx�7=�ۋ�Ҽr���%oԴ���x6)����w<�m�9��[e��g�x�o�[QwJ�0��.�7�S���O�O�|^ ����y�t��6H�)n�JV�i��'΍e2���3 |�U�$	���D@�������4ȭ�Ҩc��K�l3�(��M�Md-s�6�浰��Xd�������s�Q�jw�g��y���Ȳ�2�<>��!�~���ymy2�o8O�$���Nb��j+�(JY��֝�z6+��Vſ Tܦd������Df4��0M�Fg��4ON�7�i�zH�ҷ��:���-�so=ė-}idǬJg�	=a�f��>`G�ie����)����#{����@5|�?�H�;���a�0'��7�-S�K� 6K!GbQ�\PԬ=��&�Ʀa��c��,Pn΋��/@�y�bF�o�o���	�����kh� U7��禊y��lԐʫ�6��$������3���N�iFu6�h�n4muh��q���(�Hg�gLk"�N�E�r����Q��3���$���)��O�G%cԓ�'F[�?� �t�L�U,�����Vr�u"����L��5���$]pT���A����w�>�����B7�?Q����m=��>�����l}Ɇ��םԁ直���7U�Ƙ�&�}˔Y�����Ad=w�"V�*��:;a7$<��eyIG�4c��Dw{��,	��*ě�L�r�C1���@����!Zw���25�^�r�LT�pC�f4�#��A)��;��U
4�t�-�F�ti�(��L�5�a��c���2�P��j���ӢfR��q?�R�.���ݯ2Z�R��$��T��)�n�.�/G�+�KW��[�B'����ݝG��bt�V\hy�^U�����pT���cY�����Y����N�)>ф� �(�Iw9��/�q�.׏5<1�U~6c�;��]�co�0�k!�1��ar���C̡Z�7B��_S8�J�7W� �q�������V���F�5̈fe�5�W��Q���f�~/9=W�fqeZ�в����.�9�>�)�����] X�����a8aE;�� �N�|�<��u���,V���*$���m�p.I���vݶ�؛B;���z�ʉ:e�Jn���7�V_}Q�13�����z��� lI)�P��h-
�O��T���7H���� �ӿe$��͘ӏC�L.ɻ�b�|y��2A�u�%�L��%\��s�;�:%�k������W{�O��>Ќu%Ɓ�(_�K�u�@V�NWR�t�f�a�]�ivN�Ґ3�ޫ�e"��~r
&WC��Q����g��I�������3�g�*\��M��[���e`/#���%D�����Υ��L˦<ɋ�v�$�2����V�8['&��Q��B
�+>u�6S�@=D[��^l�4��>=d���,!&/tV���xG�]Š� ���	J}�'_��QEi�v��2nbe����#ػP�X�;T^~u���+���h|��w�`KH?��K� �yU�ә2�N���B��RF���QP#��W8!���I�Q�Rx'�C��˹|h�PRϊ{R��\��F�Kmub�}��ׄ���^�P��-*ې�p�������j�nI��a�S"�N�tW�cQ�?[��S��*e�Q�)ⴂ>��\�&v�luY�9�<�Qۼm����A"]C(g։�$(z�ܺ��Wv�X�y���8�,q;�d��6���1D�߶4����`x��yiG^���̝ms[%�ZG������F����^�v�u�[����3�~����[�aL[:u@�lj�Xd��\''���D�^Z{<ѹ�V�F&�|�O��Ö�r�3�6�A�e���r�'i�4%P��*�rZ�9O�����#~�1���a��j�[�W�_��v�#%���
L<�t��	1Aa�8�u@�r��6u���YIo�P���5���ŖX���)��\�B�pqFw��n�sm�ȹ�ta=��A@Qd1C���G|��p�`5)Y��2��堛��)�B	�9���&��v�=�L�;�_��ܽ1`�x�u�͛�I�;���>_�T���Қo�善d	�Z����k�A�X�����.�r�s��nd�0+��@�kp*� "g�:�?����ێ���-)��5b5l3�?��^9,vU\����n�� ����%��(P{a�»l�5.��Q;F�?�����Dt�čJ씥]ȉ����qqG�R1���}-7�z�L��������������W&��J̔�Ő��eRؘ�0������!�p�5s�Q���-�,�k:��[�/����ZnzU�W�̊q�]��&��*�E� �H��2���n��������P�Ȟ'�� S�`w��7������l:�q!�I{�_e'�2�f��N�8�c����)mv<��]������Uޯ�A��w���<e���?�+�86,u5=�J=b$������z� �T��Z�ҏ�>k�����*̰2j�踣+Dj:U�KL&�����`���-��`.�hŮ�� ��ԫ[�iB�~�ri���#V I8�*�/O���ɧ爽[&��RiDX����R9�򁆩`K��I�V�{�E`��}�aj��m�m�K��-�6w?�ˬl����;�c婂�d�J��ʽ�4�4�I���z{_�Zjm��"����9�JuJ��v�P�#
�=�c���gtJj���_�l�:XN 	����A��gY��?��c���,i���>�O�(�/gs*{C&��zfi�fo��+�B~Ú����ͣ��79i�9C�ʹ�M�KQ�S�l(��������Yq�*��ڲ1x�&�6T���J�[M��ؐ^�\-�Yh+j�հ��_1���u�;��E�b�dS�
3B,��q��sa�;�g�������x��a��+��T���'T�}�Q�H�^�a�����˧���\�,��)��l�Qj�ڴ8���8�31q�A\���Tp�6�NG�y��D�z���h��~�����r���^�`�s�܈���3G��쵞�D��a"N���Z��B�q��M	4�F]o~���K��_�[�';V[�oŬ���H��ƭ˒4�sё<�N:U0��R��T+Y��J�p^��9��o����������<ġ��+0�Az+�g������V�����n;�8�� ���t����s���iح?�G*:��JQ�X'c�èD.:��Ƅ�C�#N�����.On6.�&�u�a��׿���U����܊�ٕ�l�)]�YE�M�t�@
�V��z\�w^{�/�8�<�\�%���n�_�b�����/�zB,�|i���P{+�I�+ZjAvr�W@�,����jqb�)-�2������_����1$��D�y&�
�9�֤{�M��,c��C_ʘQF���H���&�Mmݙ~4�;��O0_
!���rK�JCX������4�9s��\���I㈫���e=�z�L��ɭ��A��h�����7���c<Zƀ��a�"��˾�����>pk7��V���^����R���@�qQ��7^���J-^G֔��ܝ���R�hE1�����̉0��Ꟗ2�`l�tFր�k�Ws�r�1P��us�6׺����}�LI��ӒY���|��+�뻋��jZ�cγ����L��Pw���đ��6��s�tzr4�F(0*4���Pp�ʦ�����,C��vJQ@E_�)o���s<�� 0�Y�\(ȯW��v03t�f��`ɮ����xt����a��-���LcN\��`6_V�.��}��UpЙ�R�m�@jN0w9���mPfT*�,���E}`�����ϯ���n�	�B����{,�j�����>S�����1�?Y�zr�{D^ho��Ɠ��6�K���?l~�f�Z��T!.���3� �#�T�K��P��	��Z�ƪg����j9#n˽�x��]s�:^}[��MQ�'T育1Y��s#R�M�i(�3�Ա�2ٳӮ���.a��UB)ǌ�|>G��(W�	t%���l1y��La]�~p_CſF�z�pi�ɑ�{�B@��w(.2�@^��
M-���BEv1����m1m��䫼��n8�z�[��Ѻ���oޏl�M3'>�nzΨٱ`���������;�-8�4c���V����zTg՘&.ݗH�ud_�9k]z�Y,��=ӝB[���g�X6��x�{�I��U4�u��q*�×����"2���(��`����&����) \獒2$��%��ׄ��-����k]y]�V���!���m��L��,��q��W���������=����Lpl��6��;�l�b��A@�+�,u��u���H���7TD�����	��~��c#�p��A�⎠>sOV�����B�$}S�B�i�	L�W����[;EajF�m#�غ"pV�f� �q��C k���$.���:)��#3f��YH�$�۩�o�q�oW!��欂��P�:֘�78
1�&�E�x�,�
�O�z�P���A_������ʜ"�fˌCs�|a����"jD� ���hS}[uu>3�cz%:��.���VE�cP�,���	�ܲ��N1�xT��0"�����ȅ>hZͷc2^�>+8��I��pD�/`"�ԉ� ޓ�h����c�8��4_s�����`������֙��ekK������7YP�Mx�7:���v��#�	R��Cp��l]�V}A$�>:�\
F�M�[�Xk�fH �8�nW8Y�Y��]bf}p���_�kxs�۾;V�'�ع�Ji����O�E���^e�v=�C�*��]#�+y�C�}�	�[�if#_e�.�rf���D/[ggJ��\�O�z/+d*���T����k��Dy�c"k���aQ��^HO"�ģno�pDH��������8�3��O���_����pK��{�~�G.bW�]��.!����������������$��h�+Y�L��|Ԣ�9bBil����JE��	�:*&����"�������Ψ�6��n��99{n{�,^�.��F�|b���~���f��J�wj��y�y��{�P��ц�7�Y|���O^�-�����O����O�l<r��:f�c-����iy��������~� ����պΠ����R3@�������}h���L��1���7�&t��\�yN�=�q���i~�`;�v�t��[ ]-q&�Y�����(@�K,%i����v����)n��(7Hb�"�N��/�~c'V{�X>��>�n��N�gԂd�yVx�������ծɩ|J���
�,uxS�:_֥$�����GG	k{�KS��������j�����W��tFqf	���> B�?f�^���e��0��o^�Y�d�#��#�!�8򖌜'Θ����]:�z��כN��dr��\(�l�k]��|1�?�IH]��"�vB:�\0w+�m�Q��I��/�r��²ECB��@�9��������i;����D���֭�0���Ӑf��i[f�~�}��=�.��(ΰ�܉���A:�\90h����
	�Cn!]%�-�7e]�7���cL
�@~�W`��y�� t�Ga��*�o �t�������U�#�����ߑ�ˤ� }N�i
[�X(A��F�
��i˔�+�������/�*]����QY�i������]=ଵ���?y��9O�gzѤFaK>��-:�y��=�.��2i
�����)۱��û�/��%�ͽ��g�1M�Z�C��,���n<��n��BU����-�	�24Ga9H��W{��82|X�D��_�wHu5eO~�<຤E��~#ǲ}Z4C��tq���^��k¸�\+�I�y�/�4}B2/��@�Fh
�T7BA⨎AP�{�ՔG/ݿ E>�<��4�D3+í�(�ݠ��|ҫ�����2��R������w�I:7[!Mw�q���@΃��y��P�Y
F���S"�cz[����l��`�!n'�ЅbB�"���޵���8 1�x�n��5~/:@��b�q6�7���8j�I��6j��3��bfC�"�7�I��͡�6�ȱ	��{\�����a���q����q$�w��v���ߌm$^⺾?����kr��V�s��-F/w��ZV	ٙm�e����>�dv;�=�;-|em�ŢQ-��tiRM�k��l��f@�<��M�����э���|^��l#�L�\4����%����5Yf�
��U�d�@)!/�Bw�؁��&5�	�3]s�ڹy=��� Q��R3w���E�R����>+��`��M�3`7gtĭ�%���l|we�zX��$�Ej���XWj?^���e�z|d�D~I����w@s��	���x�ԭ  1��m��8�[;��O��)�K��c�q@�N+/ZS�N��f3���{�,�bW1�s,�Q��@��T��r�gxR�{����PPf U�H4z?���EMF�3OcK�N�]��+
 O�G���{����K-��S�p�<�t?㩤4��(,	.!)j�ӈi���
ժ��X���Y�UFa���I�#�ց�i��}r�iC���g<�2���a�K�շj��%y�F.��S��&���逶��ю�;�
E#f��n;/:�И�@a3_8�i3��/ν����gr�K��;J�+C1�a�?�����H~���h����Y�
V���Z��b���F�<���$(d mq�4@O=�O�E�?�I���I���t�~�-�&�K���<�V7��A�R�/<_z�Y�L�)@`R�[��/��,"[�i�uC�n;A��w��餼2� Z�``סm�2_'�H-F��Osvs0K��- cd��҉j���'��Sr��9�>��ޅ��+��0.�+�����/��/	6ۉ��ן�_o�|bO��9�˃�S�T�PPf����su�'��zY�2��m���Vr��Ax�^�O,3B괸�qA��@���Tؽm �w�z���t�sߒh�!��c�M�m��
BӘ�I�8Z��-����4���ҁn6|_�`�Cj1'�LK>� ���j`�ɭ�� V=|N ��4֎��'��|�XH�Y�60��R��6�}��:�1��^�*�S�k{l�0�U�;]��#��'�d��z���3Ow!-�/2BA��l����w��tC&<����c�4b���	v#�������P�y0� (q�n�8��޲�/w���S���Uף���Eo�#��/����9���5���&�`��2f�6�d��z^��hP���B��E���x��`�z�l-�B�f�Y2*3��-�+��ѐ7�`�z	��Y�ܔ�!�ֱ�w*�b���Wk��-�ᵗ�S��m�0���w�7�ɬ��T�Ē�AN�;t=��Q�<�Ж��{��`�Z�C|u�B��z�m�7���v\x=?e��El�[���c//\�K����H��r�ٽJ]ǴG�a6Z+�����&��1�p̘�����p����.�����"Mm1�_��/�˫~��G}�?����.^J�~+a�*��>�<��pt�fd����궐���;��8a;8π6)=u�*�-�\{�t����^�Y��`c,�~����u�yY�W!��9�n������q;\[�O߯O�?�� 
�,q��%i���K�T����a�pw��[��	�D�r�f�CRmm>�4��2�^�&������ϱ���o��=�"{rZ7;[YE����R����&�ľ�Cp��m���_�I��Ϣ���$2ͻ��3P�A��k�����~��O��7o@�Dw:��"MP7u�P��G������G(����_��\�ֶᖀ���e]���T�a��T�N+��ռ���ee˸U�:�a*�ָ�G�aFT1w=��� ��-�H�TS�?���C��ð�>l�w��Zk2�oKkQ[3�I��~�Q5k��@h
%��4�Vii���'�Eݔʆib��Kx֑0��x�̺�Hg�J��E����x͈z��_��x�y?/��P��O	��ޅI�<����q�Ow�����r�����"�����x�r[�8״��*o��|t:�i��<��9�/a�.E���.$�a���=>�(�����mA�:��|���zGʅ�Q:vˠ^�����0�I�x�ԖH0f3�'�.�cbC����j�mŸ�画[�y=R~R3��;Fo�6k�k����0)��h�w�SHa\����PB��v�k{4�ǖԣY�J�]5J?Ji��}'�ۏ���w7�)��+��yF�N����j�U<͘}U����\E�A�L���Đ_����u�����F�G�.���Qᵊ'\jK�3�q��s���B�������!̏SX;�-@0�ղ�Eӫx9�	��������3#�ޞ�
�����>�я�K���
 =���^A����,����z�٫VƈI���X:�7pȗ������t��=��9��F@t�u��$K�s/�������A-�V��'n}w�:��c�Ďn���S��M�@n�8n��8��.d?0i]ۃ��
b/C?��X¢�hڵ�+�*|1��4?��y�)��̗Q�M�,�_�h�����t�c7pA��N�/�&R`�z�:F�i�ã��鷱�x��q0B�`MQ��������������������H* ��5��Ҏ}l>�}��ww��1��x��B����G$���R_�_�N�/5O^�a��Id♖9N&$�xw���רw�}�b�x[*{0�*�Y��� �J;p� �d�.�6�fLX�����h�s�7�O�Wo�O<�E	/Ė3��ްB���.tQ{.ɗ�2Y��Bˏb^*6+���4�����!v���v%��k��5b�19ю9���_�8E�+�VЂ��J�k& �<\�
�"���-���p���cĞ��E"-��54�>��Xw �Mڣ;zr���i�g-]o��|.`�m|��
�9�A�,��zAE�CO������/$��!�G��J;b&��ǲ��2�SҘ�6$�Ph�����o �c��c?O�'�Z����L��}��x6i��a�� �oL�9�Ez̧J��fxx8�����Ě:�$��-�g�$�mbE�`�`z]��0T2���%�k<��W	��|���]�;#w��Ju		��*U�Ûб�� �V)�G_g�cz*��D�i;�r7��Y��O�>�gr%�I�Qי1c����]����ByzҦ�U�Ȍ� ��+��t����4�t�1��2�!���P�y�����A0-�J��s��4����c�V�F���⨈\u��KPG%�� l�ÝDdoN��h��6{w%{j���5�4`=�)�p��q0�<�9��O��&F�fN�QH���9%M�_��͛�C��0=,�:�ͨl�y�B�n�_��| ߗ���m�Q�Z7^O�=�w�P-QAp�����Sm�?4�2��	�MW 5:>�[�2�����[���/u�,��*+de�-��*{��훈�0��}T���-��t�)ā���d���D9�N<Z{G�\�ky�ظݙ��j�e�1xw��M$x|d�8���y.���l-��R�!n9;�δ����,}��t��<�8����|���6-H-�-��x��/:�L`�6�6��\Lj�F�ɟ��Uk:^�\gI&�qrE_��?/���F���g���I[��L���]����P�g���)�h=)5���$�&�K�Y��kq�F'}�v@w!���n�VB�������ذ�3q��RҬG��]�<\>���A�G�;�&����"�g�ΏZ[h�mO��!�0 բNчH��S�.���~Y%�E��p�r�
S?Q"%xU��Q�L06�g��s��j��xN�ql���t�
!����,y����3o�F]T]Q7͢8S�����D�V�,O#\΀@M$,`T6]�d?2�����{J��S����M^	���C+��"�H#f�[m̡v19��q��/�S���g��*V@�P��R7�/��v:�N�;�`�T8
2�� p���@� �Öo.%&X�#9p�<(���������c�f�L������@���T���y�W��,���=���i�v��b�n~ �ͯ�y�-���꙾�]9�I ��2s6i�ȓEd�6����Ƚ�p�rf� ��1:��"��
�hѪs�m(���:�m��-�B��n�z�Ɏ���[��g�CCU��w����l qĈgf��A�
_	�<D�]<���Hf�B6�)  �4F5�M�|1�ȅe�`����$� �g^�!I/Mr'��Ν��kT�6�;M^�Pn�$��:���F��i������f��P���]�B����i��.�T2�(C@�]Xv8Q�}C�q�O�o[N⌮�yQ�����3��&5r�"��6F�<��i�.�]>�9��niIcX���OW=`��,hG<O��v���q�K�s<���H���_e��Y���pg9ס��"�����¡C��d�ڬ��������#�8=���c*ޏ��)7}��,<y��ޔ�v{Z#<T_`�P2��	@��g�hVG�� �Mc�β�k~{�4[0�V��_��5:oy�0��7QP�I��*�r;�B6]�����
��on%�vI��9Lri%r�\ ӡ��nz���Us��H?�1�>�ࠨ����_���1TcS�(��-�ɸF��&�/���bRӯ����R��t�¨"�B�Χ�W�(q��v���!���m3����\y��V�ge���@1"+Í:��׃n�Y��to����k`�$vg��e� 
����֛ �Ѷx�S��WM�R�g}��rRm�Akll�ҿ�;|Pgk��tҌ~Vxx�e�!�#&��FZ<Cs�9HR�W5[l�
հ���#�]ה4f¦&��_q��+�]*� ۦτ�R�0ug�dG��fk�V�<HC����(�KoGȸQ<GAo��>��\9�@ =͡���wQ
��Y�[�>A�HYp��.fp���e�d���i
>�-b_�z���s�1����o�iE����7l���*��/�@o���_�l��nLn*y(����YZ�k���?o�BG�C�p�k�sS�P�8���k�XCk��xK� Uy���&�D�����l��T�Z{��g��lJM|��<��ē�Svr�>�5芲s���/��H��aY����╛�DE�j�@EF��,�cV{�U΃*���|i�_u��]$|Ь<*��U���+٨a�$��Z��
D�c\)�V�_�J4IFBÝ=ʓ���\s�漦,����u�k�%z���7�.Q�vRT�	P�[���_��JX�	��������C���S�����DX�e�OX�T��*ҙ>�����3��A`�^���B�~L�.�Ŕ�'���f��k;"�ʍ��=_�k5���t=⾇b��p�+k��2��X��	N��T?��`����t͓�O�8��*�C�^;���A�X����I#�X�Q�E�
�'k�ýq����d��GyH�A��A,0{޳1h:��`�9���v}�Q��d������?� ,�h��᚛���Ld���d#0-|�l���8(Ǜ#ⵣzrNI��!"bX��u��9v�'+��C8���w:�����R