��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��@�yU�ߢ�7�k�U�U@�FAh��D���S��T��.��8��8X��l+ H�YHN���DS�0i�>#bs3h]�^�w�(Np���1��q8EV-��Xi�]S�M����OJ�8���owmQY�l=���h��^N�I;����MS����*c�	�}ͨ��p����w�+��&�(��*�LN��Ԣ�GE~@>���1�Tj�.��G�jcc`���WY�%>��x9G�M}�����Y�K�<�BU��q����Y�~8��)+�fpH�QU��8ԠW@�K
��x��x�6u�2apz�c~iZ�־�
I�:���{>��+Nu�Ak`� ��b����7l��ګKՃ��ؼi�fIJ@�v��|_�,�$<]�9#��8O�f�0O5Pɒީȱ���b�ﲕЋ��e���}v#����M�az�R�Q�|B/3#��`�]^,o���XY����]yr����vaD���ƀ󶲜
uK�v��NNbi/�:r�v ���"��%��
�THOY������̝aD^;�+����ݍ謱�k�3�U��f B��sF�uV���-��1r��7���Mk�-S]t���si���,M�^�/ƫ}ު�`g_�H?X�$��Ym�f�zĀ�I*�O����t__-:�"���ry��ƙ�Go�G)=�,�#�C�@'g"k�5��/]����!��PFJq�vK��4/��i�Fl�p��j�*P�NUڒ?�@p�%�
��t�%s�$&��Ò�S�%�n��P�W�+N[9�B"`p��w���Vzt��W���!e z.hS�"Y�!�qr��0���ːq;#�3��R��h
�c'��v�	L�]�~����2�!0���yI}��r�r��}y,�ۈ�âFq+BO���k,Ƨ;e�y7�ɪ;0 Z�z`ѫ��~i�6;Rǆ/�N�TB63�Q�����\,�j���5q�5��M�Iy��c��=jh�������D+|���>���f�J���<��$6��f2a�p�$���rY��Eb&Y�T�[)J��f���ـ�N�� ���#�����q�Wzdh7���W�Ć��2P<Gх �_�������w��U��م�e�����[_=��(hIh�Rި��6%~|��3���Ƽ��T�{�!����6Daͷ�D�ƕn{N�΁�p�~�̗��/�(��D���gD�Q?Բ8m����!��3�*xNur�%.t[��_h��v�kC��Ϣ���I�Ǝ[D�$�8�v,�P��C]1� ��S��T����0ݤ�l-A�Z�ݮ/]h�0�S�����E�rjq��Q�b@��n���6��܂�%5��
N*�9�8�����䟑v�D}v'�gr,����e���Z9��nu[K�{'���Pw�vb��� �{�GA.�&w!���u�<��ߣ�{����ޥ��)V;���������b��Au	�W���# ��J~
BU?�Tk\�r)\���zE	T��J��G�p[��T��ڤ~�A�$��H��4V�y��|N�;����̪�;�Si�X�*a&��GHtM� �������1���Xv�8~�2I��IҚđqGt���}�D��M�?� �]��wQ�(3�xS��'��V��REV�k��V��h?k,vU��XZ��V��Nx�Yӥ	KGx��/ ?�PS��O�	�V���t�����m�v��0Qy8WX�x��1�g2ض_��$�&�1^Eu�_]k�E���YG�|����C�ʙ�
�x�Tj�pV���v�.m�O@�<�xblM�F²�����c6_3U��9x�;c���Y���e� �f]��S�Ң�Rӊ��B7�c��e��/�wv76�Y�	dN���;)���
N�W:E�9g��U`�4]�����>0���%-��A,��h1)���Opx�
�w�C��MS�m���5�럵�Q�[��Vc ��V"���ej�e���Pꘫ�␓��߲�$� ��X Q-��.��!az��s%��J$�DF�{�+�]Ok�������/��;��� ��t������o0-ߑ'n@��mS����{�m�UI�/³EAN0nNz%l��g�S��a)~8�ܼI���gɥ���Qvޅ�FI6� �������<���#{(��]RL[LY�i��H}ޢ�ϵ��R����Q��^Й��MC�g2؉�ӔR+��C^�U�,k�(�p���3��+N����cC0��Ț�; T�f��$����24 V<����j��j��v���{j�L5_�ew�\�"
-��Sц��S�'$᱒ܔ�q�+P�z	$fcmrk�>�Qyf:R���F�GyĐ�O=�=���E�x�Bn�R�Z=�ܨ%w��O��o�?1؊��&E��_S�p.�������JI�؅�V�	��bx0��^<'��Ķ>Q�p���ۉ��'�ƹ�,����v��y�0�A�o�X�9�^��,��9&D���� JC�V��\|��RS��ηώ��4�:h���<�x�M��4#94����j��=�%�!����º�,�Qx���9�Do�L���)��w�P�{��T��dc>�=�+���i�gՙ�
a'm���Wz�����q%2����*�yL!ZCH40�g"3���1 jK���P`0_�O65BU��4����ǥL��g=��C�[KV�����_n�O u �]�+m0M�k�Ⱦ��(��瓄�p~����w�@!8������	X�k3�H�������s���������<,���FFc3(���%2�-Xp^����J�E��b�_��G�x��L�R`��
���WF4�������d��̴�_=��djZ�'$��kc��b�^��2���w�6���<O�<��oæ����M��dECNXa����/JX�!��ʀ��Ub��������+����%=����cz��$��[Vr�������7�c[䖿�8�i[6x�y ��:�kU��&?s#�_P����`��L�\������&KT ø��8�a��L�u����N*�$�0��O�N��%������}�$�G�>l�6���$˿z,d5F�p�8}���O�[��mß9�n�*N�w�k#>��b��>�s�?��a.�z�4�h
����e�B~�?�	%��^V�����3w��'�)�S����p5���+ǹ6��.C��3	`X#q�@F|̈X��� �K
�:��>P�q���vr4yV\EHS��Ԥ��K��X)��>�Ttx�o(1f}#a�`�4��*x*���o�Q�����FF/!�YYuT�b�&�&(K�|�~#��Ajİ�T��L=��v,���p�X��bw���$b>*�9Y��@n�.qby��̼Jz���v�./>�$w���;�;D����.h�pK�m⇱ͮ�)c����˛i�JTBCk�6r|oD����,/�N��9<�_�⟕B���>o������w�UpًX������Uf�H��:H�(��Pu�~v�mڶ�4�q���$���v���9�i��H����ٱ�dlF�3�6��>�ZD���vI��
�� �N�:>z�>if���젧]0�`�tey�I�4"���C�*����c�@��)M����Ț�(����sW�����[��"���^�8�a���7V�L��lYx�������?ǅ&,�Or㬁{(	������wdF�O��zD���*��l��뽏�<�>?l�2���ΰU�K0V����k���9_����Yqu�A��_2��o<�A�����ŰΚf�4��z�%�����HƜ��4EMp���Q,���q�1��Gr�5D�j(҄�����({�7_���(|�)���$�$�#FhM�|T`��	��;r���̹�H�ܩ�h��U��W��71��rE(#�?Q� ��b��wp*�wP�B5X�"R�S�|	K���1�0�qv���ǾbBL������#
6��&�;��󜆡����Ƈ �]�������>a�]�!���KS��/f����9��e��&-"Fd���d���"�_α���M�A?��+!k#��F],` �(�;�ľ�p�хS�����B����ԩ>�?E�Ȭ���KL�M��4�+l/N{�ߣa�R�����J3ƢO���o��1�@�˟e����=�E�60�F��[x5�N������Kyo'T��_�4;TëTcY�a��v8��ٜ��w�%�­�@A^7�"����ny������|�l7c�j�oj�����䵂Q��zB>� Fg���zHӊ!�l��XN����'z��aC[K@W�_J��3|�!�����)�\�b�Q��[y-)�Rp���&��J�Y�/�!7�d>3���.u����u9s��`#w,*�[l�����Hl�OП�Q@�:N�[����/׋��*���nT�6v����zN�����8���X�4$j��\u�f��qx;�ʞ���Y����7��9�������"���dX��Y.�{gs�wy��Ƕ?,�fq��i�(����-�x�c[�Q��)$�{���`��RGC#ʸ+�hb�����D�W~ /�U��[���0��:=�w$�|�(�+&��Znդs�0�
^C���I�8G��(/��&JT=\�	��H��r96�N(y���5ʼ<�׏lr����=�����<����_j��R9�ױ�/ƙk��h�14۽~��P,�m<�kX� �GM��nk����HZ�m<[_vW�e)?}'������3�]\�ۤ8wU�7��٧�l6 5\������L|c�{�m����e� �����1�߭�"�*��V�
 �_��n�}s�� ��P���F���M2b���pL���D�msר�s�)�:E�R��o�FI#&S�&�OdY�6���ĳqАl]X�&�b�@5LM��mXc��@�"��B���r
*�=���4[�n���^��F+������D.��a����H����g��y�����,/K��0a�`R���5�2�
ʧ�L��8ܘ��9��Gv0꒿��)�&-�{���o��]�
��L��Pf|�<�?��yp�n�A1��4؇�͓�53���HpXӗ;��7~�â����e�,�=�A���'6p�E{�ʛV�o��4I��rF�m��v�@�.	��!6�����auEL\Y�n
�?uZ6�Gau��^2�e1��]�~��2�鯍C٤�ԐD(r�W��v%5�K�|TicD�<}o���������V�т�Q�ӫ�����Pu��ɸWN��.!��>�K'�_�)��]�sx(�G6��bP\���=L�4D$��fg5j��������K�Yia�& nZ��.�
N�.�}�b9��)�o83�����`jַK8��A�����I5�.��epD~�0��G���&>G�-��,�z:_Gl���u�!�Ѕz(CL��r�4�,�:)V2�#��ޢ�_WE�8HY	a��>y@�#ӑI�sV}�p��N�����%f$�T��1��7�Tk�b�v��DK�w0�pah�~�5D�Lݯ���� A|<�8kZ����-�3��������h&9D��_H�>���ޙ�Qu��(>��cbsR�c������=W.yFp	2�-H�XU�ș�����_E��
;�~��ᆁ��u ;~��L#��j*�!��$�e� �s���܇ak�j%d��ݝ�Q��|�g-�'��Ab�{��M��s]� +�1�����r��c����Qi�B����VI�v�~�?���uv���{�j*'X�&��-����ï]�gPiB�Y)� Q
�Vd fd�e�

ҁܨ>ɂ�?�g[,!�nt��+B-�Xe1���ʔ��a��k�'ŔϟX�CB0�$�8�����m$�t��{�����p2?���v.(�6
d�b��V�*�A�|ԧ:ˆpJ���֫X�L�6�u{��h��R���#�bb@6�m|�t`�ǒ�BQq@yT�}����A����)��h
gc�#���2� �v����?�v#L1;�Z�tɋ{�S��A�UN�x���X�0Ǟ�c���Ƚ�1����ۄf��_~�y)� �~�"]��*I[ n�2�_�y��?ʕd^��j��s��(���^�򱖗T��M�]T�M���8/��kv.J�E'��g�o��$��م�֊`}���5�'9L�O9ˮRʐT���P�<�^���Ӣ�	Գt&p�����t�gBW���!�`:8��Лn�AQ�����Z�ӌ��F�-T��X:���=�:^ײ�/���\r��[���e׷�?�p�9�&��T�ݗ�	�����a������F2��?���5J-X ��W[�bվ"`���Ha�s3�v,B�2��d6o��G�C/vܛ;��Vh��U�W�kOL����$�`X�C )�6i(��֚Uܒ����S=uc~sYQZ��t������[���^�D�7�J�X ���UE�����Ν�;<�>��$��=iA�Sz�S�ZG�C 
#�4�=E���ie=���:k��)q����o��u�L���W�$j OF2�� �h��'x��
ιm�|��	)�4�'����g�,��YP�Uy5`�]k{���
�ė��!=X�������1/��=J�pC�x$,v�`U�����upEr�hJI�F�Y�dK����n^�+��Zó�4�ol ��d��$l�A���{�+u��^�PT��p/�Q����;`�mg�恻_�S����E�>2(�;3ᴆ������������B�]���-Od�R ��;�U�פ,���x�W^ql$�FA�:̍O�՛��M>�
O���P8<���՜T�"��A����e�2L���F㛎H�����6���/^�#��X��A>��+�?�X���B����0�!wNS��ͧ� aUxt�{sĨ��bM�h����2Ԝ��BVO�����^����J���G`[
 `'^�oE�k�"g��J�� ?����BV��RU�Vx=�O�Z2�,Y+5H�d��.������k�䅶VC�Ѡ�.y�ED���+��C
Bӟ����d���B�}��x�c�w��w�$�n;�.wTjm��
V)�>WK�c�]AA�d�; |�OK<��ChWE�F����T4Ʃ��4��H}å�����\��8��D����������5� �w5��إ۶W�${�r�u��Y3�*�"��4sA'SI] �ZO6����A(���9�P2|�p�<{�M
[Y�g2���6$������Q��/���>�RK5�#L��[�Tj�Gܙ�FQ"�	r��qb�B�2f5�.E&������A���,\������#�TV:G�%*.���x�O���pK����@�##Wg��gp��)_��Q�j��9v�_gVx_�x�T!pz���f�c�l�hUo�B�/
A���OdQ[l`G�×-�%s��<�ًS�:���i���Q�9����8ϒ�t��8^x�<IF�������ub�-�eR����N���A�6/E�}u� &�j����'��
z.�y?/N2�?1Q�[?�3ms������r����f�̘@���q������f{�ߨ����k�P��o�ΰF�Q�mي��ֈb����g��N�tD��4�yH^��B�����'��ᩫ�[�0f��Ȼ�!�@��e���?����Yhmp�F���'�	^ip��'^��2��.��O��OR_��S������8S���u�y(�۷3ݵ��dYP���	�����^	Ƹ�.Z�R��x�������!�Ywj��[k��ޑ��R�mJHYh2� .uD,�t$�j�ܧ�U�>�'(-:G<`��u9W��0�����_�?� 99�k]��h���L@��雘�&R�Z�����Q�����6<�M�U�MB��3����)u=��Zv�N�-k�D����.-fn��RL5z���P#��|���U���/CU�Je���K��f����qV#�<f-�MƦ�.e����S� Д�6�p/�σ��y���^��Uл�m��NTa� �qC�ҕ�
�F�!]9D}��f���$;xu��E�����f��)T/�S=�_ä́����A�r��T�O�A�x"�=�h~�ZF�:K�I�[H:a�2"��i�|$@/�y���o�J=��.�;vO�yK!C"\��ݔ��AP�s��]�[y7+�	����0�y�-��z6-[6���'��Uq���>��������9�d�d��\�����j,�Q ������o"�Ǧ���"R�qJը(;�3tb���o��'a�_�Ծ&���8�i�kV����Z^��	���n�l�c��,�D 1�&&�6���E|�p�}�"��E�%�� �(�����0S���|i��ҒO��U//ނ	:�*�Rn���=�z*��2O�s��óq;z]�,|��������2��
��b�\^�G�Ү�҅lr�����(�E`l��x��@n�B.��x���U�E-��\Ch��Ș��eۙw�i2�Cf��V���\��r��j�0�_�2ѱT
�\�%��T Zk��w���
k�e�&�����u��:��m?��eR�r�!��PD��ǘӵ��3�l��E;�E��e��]���A	��]��c�YD�0Xw����m���d��d�t�tL,��{�H���;;acG�����V#0��c�	5�_N��p5�	BR&�%L8�:>��Yj�����B��ۋ$2[H�z��)j6"bY~�?�t�|y�}	r���l�O��q�|�4Z��ؖ���Gce�$�"���K�w$����U+��(��c�~��0�#�8ME����/]4jDB�Aۈ�d�2���^��#10�l8G������=j��"�|ᔽ�#
e����K%5�vs� :��?R�U�!䒻8�.Ăөi�l1kx���lՈ��j�˨��ϖ�����$d�zbRox��7��3b�c�e��~.~r~�;�5����m	`����^��\o�Ao���.)� �8@��'��A(# t�{�%���\�dO-��I��D,�-�
F�����rlL��¼*��^�ATj��Lt�FGo��e=Q��c��u�����AK@� Bsv���=�s_V��0ڛD����Z�y����-@&����b�ϓ[Ľ�jy���f��n���	Z�K������Q�3@�ξk�d4��y-��&>T���ة�XF�����t��o/��W����9к�eh����Hc��8X>:8.��o�s�ţ�X(`����������BB&R��.m�Q~{���s5c�;�W��E�WC%V,��t!EbpSh���l[Y���DGһ����mx����*�=�'��WHw�I��0�2ض��F�X�w�V�
ܦ]8�Իq��O?pO'�cG��D̐
�ec��㞲,]�Qy^�����c�x�-
���,��͑��R��1n��U5�7w4��4��� �f}vo��B��"�ƴ�呁3�)�p�摓�B �I����������t����ҨxI���/[ff��2�K����8}��-\S��m�c������"꽗SL%[3�h>�-+�[��V�B1i�tf��)�w���Võ��u���	�K�U�e�ֵ,3���Ñ�c@����U|q����-V}MB��G�+JR�	��+:�(����&������tV=
�9�R��L�8P�(����;wVLEJ{���h�)^|�� �5	�ߣخ���B��:��A�=V���Sb�`{����zN̞���{I�Z�xO�<T,�!m�3I�2���;G�Ot$�\Ԉʥ�8T@�,�j�H/
X�h��9ή�.��n�h�{�.�S���;�!���1�N���β��]��U��u��7cʪu�?�)�B��z�պ7���J* o$os�K@����s�o#X�m1G}Yq��N;Y!����C��>�hO5-�����"(Gľh���U�`R�5&Z�b%�9n���P65*�40���YGӇ�����S��;t�҈� ��u�������Yپ+�g����}q�'u��u�'��~�4΂;� DLY\�	�8o�/c�����6��m�(�����)#��E%�"-����~�pA
�� ���y���$�\p?}��KV3 O�M��$#��zȋs4��;�8w]E�{+�$ӷ�1D�|;I��(�5S=[�߈�N�i8@*%��@�? ;Q��0�џ����i��'*����"D�^������)UG,���C�A��hw�}���&U��l�̧�$."�"@G(:�v�x$5�8�������rC�!;�d4�?�{�+xηGN��6�w����-�?��c�2C��Mv�4�<�"\]��EZ��q[���t�7'D�<)m��j%�S:K�E�ش�a�r�(��k��k(=�mp�m��&3F�|��a� ����I!hS�ΔZ���B��D�9q1�>��_������*m�(D�9t/�C��|h��D��"_l$M$Ai�����~s����.�M6���h����g+���l�78+�	��S$2W�;��4�4!_-��#o�uX��~�=P-%�]{�G�ebK��փ�K�݆�w�O�]Nd<6+֞{��R��!�Lc�ӱP�*���zH�?�,�����L�� �p��? m�:D)`@� 2�f3�uld��
�^ց֚�T��}�Q�ߞU卓��"��'qި7g^Ù2�-S����^u������6����ݯ��0���o�H��Q7N5�٠q������,�V��)9uH�5{݇M�b����+���!�^>8������S~i�Q��(�ܖ�𼍐MMBm������T�_B�%�PMg�2^C��T"P�'� ���!H��d;C,|�`���@3ڟ�I��I�M�ý\��萧�*D�����,�)-����v��G�TCu1����"�H��[ 	���_у#"���&��;�	41������ݮ�C|WY�-�)Ј$��Y�7Y*�B�}UJ���:���$F�������.+˜��b���t���A /�ھQc��4�|Y��]���7 +59"�>L<WS�@��kRt�<�AD3�١�+B2�teҸo�Ǵ j� @��U�۩�����w�P7�������M���M���X��^}�:�f5���������PU���\*=��� Kp
F�J�u�r�b����0���_,�S���Iv^���<�}��9���H�q�YʆsY	 N8a�֗t��`]�!���$H���A�+�x�;�*��7J�����^v���d�IU�}�s��%���%E��r�����ɻ�C2�x����C��D�������̸�2vg�h>���0�X�td{��ҷX�j�2���@��XU�����(��A����z�~Jo��i�{����} 