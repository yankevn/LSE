��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��z�B4j�$}��yk�,�e�;�t�.t>��x9u�������'�,��mUN��_��3�����_I�?�~MW�������w\Ti|�ݣD�G�m���M�jw���[/=,"��6dGbm��%o���t��e4ɉ�"��u1�{9�����0:�í�)�)Y�Rc�� ���9W#�D2��g`�*d��ͱv�����G¨6�A(ƅ�F �azMO�:�?gg��R�B_ko[�m?�'��YP�XR@ʣ���]q]����}'lze�X{��_w((7����� �pm<�.H$� ��Ə&��AR�ǹ)s6^Q�(3\�����ȉ���*4~�N�:0/���D 
.�,�m}ӥw4)Tui�R|�,�z3p��OqQ����E-]��`�Y��;�����{���%0��A��t�^D�'�o�P87eI��]s3��犲��� ���}N�1Sݵ	H�H�1��A}· 0@�����9��������?f:�`�^�mB��+���V9�L7�ЌȜJ��l2��M��)��F�T���Nt�)���5K��q��KW�<��xW���e&U�s�90����3V�r���/Ƿ�����̍]4`I���^G)�.��,h��r����z����8�����ո��B�V(�Y��5��� l|�0�^��Ս�HLۛkة�(���[Hx��aȐ�i�,��WZe�c�cj<�4��;mPf��/�]��C���:S���f=�E)��"h!��?N��ꋔ�q�����㡌`8$A��=��p]�H���bJ�rwn­�q�n�ϊ�$��:𰊟�9i=�	AW�]wj<�V9�Aї��s|h�KI��z��G�(��<JK�S��e9��\�E��9��!�F�%j���Z6�no5�aN��{Mݪ���v�'�����ܲ1D9��t��mk�T�T���r��V%���QyMs�����$�65�iZ�� �\u��o'�����O��w�������C�@�� �j��r�3E�BM���(�	f��֣]�4�,�b�=j ���<ꆄ��Ć����y�{�vlT�Ί՜�mU)r�����S=��f��>�!���軽+2Sᓯ���|g�F�F��;���d�~��(z�ts�%P��A�X�:�7NT��c���y��P^e��:�e���'3%����h`�� ��/c����@nDþ����9,	���"f����9���@P�Q=J�=$t�(ގ��;�t������_��9��j&����o�k�Z��9���]n��p��#�>�,u.���*������G)YC��7>�v;P�EgC�<��(Vˏl��9/�Br�h6踷p��4����S��wb�]�<s�����K;k�h��#
�Y]ǚFU	�
eC�R��jX���,�mH�rtV�7��+ո�`M��3�A9�v'zZ\�LFKh|S��{AhN��Zl7��mi�b��!�ߝ ���##�Ӧ7�vR4�`ny19[���vN������b���)���qE'4��{k�j�.��u�����ܡN<�M#�V�E��!��(n-@�!�E���7����'&J���݄r�v\�&Z�4dc��شE ���:Oy�荡������
��5�Y���|���b3�47���'�
G.�l���5���8���%x6P�I&B�&���n�h-�9*��\ ��^Yg�k/*-t��n�	l��ASڈn���J�~G�]�l�����{:x9��h� IM�3�TC��܆
��+F�w�,-e��R���6=�
�W�|�4����SR��Y/��L3̻��!k�D:#���q��z�O��U��_�}z���h����0���Vs9V�1����I����_)��Z��Y���8{
ȭP��	�s�������{���-0��F�G�e��r�oI�%:�g�����1�B3� \z��9*ś� ������y�'L�ȭ�-,փ<|�[l�cE˒�g=�^��^���R��UHS���n���i���9Q��%�?��(����M�:�+�.��T1�������f}��1�e%p?��፼�o����s^�t��=Q�ӟ��:���FQ �R��)F�!/�2�>;��[
"*�+2�R=	�hv��%A���<7C�`g�t�O�%~�F3���	��@3M2㳾�ml�AC_����h��.��Je��!I�N�:�P��w8	펠?D �7���>���cP��W�VF̜X����8k
]�'Y�O/��$m8�+_�Rk�+$~^���.��8�S3�[�^;��ȧFz�1��+I��Ze�L-y�QJ(}D~.o&����z�e�2�7�P`XR��=��ʇ��e_}�t�Բ���@�ތ0hWQ-ЅM��B�� ŏ�N�o#��Ie�s6:tp6+*k�;��-�->v���zM8��mW&M�|�C�(]�$��8��u� ��Mk-?�	�nȿ�|�MK�����Ie�v���B\'���<��T:�E�!��$�pt��5��>�!2h�����o��	e!��akP�GP�����p�
n�̵
-wܫ{ZO`v�4����7:kD��t+����E�p���w��� 0�~�|�����u���K��ԧ���|���rUB���9T�~:O�Z�E�����{����H�:�& ��w�����5���g�9�.��(V�dT��������}d�d5�2��39���� �,7�R�:3U��ƒ���1�Z���Ib�L��%A�H�:��8I /���v��p�@���4�>G����M��FK�J�ܯV���ƶ\�R�����o�$���s�W5۩���v��7y\	hι�xr�W����)f8kN;O�$7;���i��ױ��{"����_V'��
h������0EH8JU	�|�o���6�Lc�ͭF�wsk��im�e�)��E.�C,+���kr����(��)0�r7�i�����4-�"��"t�w��WǬ1<h_\-- N�(��IPD�s���(������ҩ�T%�E@�����B�ZK�:Y�f�щ�`�Q��1aᣙ��@�L�4�^0���Z����J��-0��&=�bN�V=ר��Ͼ����l���Cj�M�r�b�9H[
�������A7LK���m�wנH�{G��)gq�<��6i��H͎M���/`
��RO��ļ�/?%���� ��seRN�o:��LW4�����,܈ pbJ`��j��QoYْ��Qd�Y0	w%�s÷p�\�i�+O�����j���q1e�/�����?�ln'��H	��(W�+�I|<!���S?
R���I)�W�*$���?	ʗ�Qz��O�R��ɭ$L0Z�~ۜ���15�q����S�M1h'_�[�c���%At��^�PY҈hE�Ǒx�w`���C����������(�N�=/���zyJ�0�YzO��c��v�y 8��It��+�6��<SX�� c@j<=�f?�r��O^��	�-B�g�	h��C�r8gOφȶ��9x	T��Q*l��O�9Λ��m�d�]�6K��~���=���8c��s]��w�o�� �L	�Z�t�98�+�� u��1�qrn��m{��{')�k�x
����m8�ab^]U�D@�u��Ì���^�ym��"T�k���k-�'9NO�#/Hܟ�*��T�ǔGb�x¡�mTZ��0���+Y9��3?���O���^��Lt���=�S9�D�t��؀A���\B6���(�����9p;��גq;5���2�|y�m�3�4��J0-����p��wBE-wf^p#$���� �!��Gc�ZL3���Zwl�X��ۅ^^N�J��9eݬE��q��1q�t1��cQ[K�{7|�Te���؈�ٟQ���f�/�1����5T�ԇ�?���x�(>�h�?h�@�$a�QH�Cu|�E]�v��1ݽ�M�;Pw�0�[S�ZNy�7��!r]�#�����H�~Q���DX)��L��-0���K	��+�M`~��ѕF��5+)�[ឱ��������xU4���\!_�����=���Eܪ-u�����oJ�e��]
l�|�j^��r�1��N**`�"Ɉ�	2���;�4��:��
���bpP��,� .�_�)c��Y�W;F�]s�Q��!�0�����8��M1^��:O��ݛO�p޷�GVSA����ۦVNȲxu�Aa �TR�ƣ��}�(�X=�yd�r���)�N��V�~�� ��+Gٚ�͎����X��ص��xK����9j3�̘U��XG�<t�C
e��� ���@Ls��9�Jߏ��qRg8]t�79'�sB긷|�p'�UIb�Ud5T&�ū��}��f���59��R�Y�@�%���d�/�lt>#o��G��<��A�f�0	�}�nP�����Ҥ;��Y�g�"�>35�I���Qt��ɵ�1J��K��[.���|� |Pq�l��$4&k˾��(u����y}�奮*`K�@�ú�I���&�j��Զ� %$��v�U*&�.���bRn��8��F�+%|�&ag�biց��ܲ�z&~�'�G��� 7�k��i��7L�!-u�W�3�����m�2�%�A����$';��=l����M-\]�g�ط�l�R�py�|��L�v�̭ �����-ɪ�>+e�&�%1Ƈ0��)�&�U~��������;���e�Ib�y[I����c3)���ҩ��7 &�)�C�6Jj�`�Y{�q�A�Pqca�6=���#/BA �� �{ȑ;c�ֳ6�#Q>O����ъ�W��1�%���ڎ�cA{n1E���J�G����{>n�넜SfC�[�~�����Ov�� �l�2!��P6)2������@q[x`4W%��j.�#�8<��H'11
�1m��n�a��H�֪�W^�u�y4��q(���k�V��^�ݪ�]j˫�p�NE��s|����ĭ�̪,�	@��5�Ȣ�?�<C�J��z1X�r<�S����s����B�O�Z�� �P���v�� n;�{�U���zb��C32��~c�<F�*'�Y[Ib�n����gc��\\84��΀/9��#S��R,{�H��R�����X�ǥ�WL���5�a�u�5B޻K�!�Nq��p�J��)=��wh,:r4�nr�m9K���[�?�y����> f�,��,��(2OD��߉n���S�6��*��p��d��B����n�gH��Nu�1 �n�l����B�v�P4����cg򍸆J�l��Q���h0�/�E��{��bs#;��'�6�ǡ�e:�p����� ��g�<�8���$�d�N.��|��λ#;�E
�T!�-!�j���K"�<� �xE>0c�1jך�������LTA�@�n=:����R(��si�{���[��x�w�P�� �Y��\�8QE#2Yu��߁�㨅ŷXg�ߜx��Eլ��P�~�H�pg,~7My�?�QT}�c�/�i7��bNy�fדp�q�P[�2O����3�߄�=r�W���Z��?SRN��i�j<��� �Y ����.m�"��1!���B�σ�.����@" �
�DwC�8�M���)g��T%�;��IO��$�t.T؎e���ٻ��?���Y!�.��:�f�s�<Gg�EN�ꈖ&kfslSzuQ�r���U��70-+#�9 ��9vY���^��qz�Z{}ogT�Wnc�i_eN��$V�,Ѹ�$O�͕��{P�B}���;59�6fϋܙ)�Ǒ����/���c�>�V)JV�(���G��A\+�aZ�u������)�l�E��� VY���r$`�YA����d)�6�Nɸ�Y�>��:�	��� ��������l<gg��"DY3W�"�+��>-�9���r��Z���;�E��i���GS�KL[��}�� ��-�a����0��8mǯ�Z
��aVr��
$�>�,E�?H_���lA!�g^��j�U�$�_�譋�����$�d"K?ܕ�˖|v���R����z��)��>;����he���9z��#�L-�'��閠<�4�*�c��g.�fc1��\q˃�P�`�F�p�w���(	u���I��F�D���1��pˤ��e� ����WC����aSYʌ��9}��m�A����N���tЈ�&��35\x�1Y���9�[�󞰣��QjC0��"c�P%�Ea*<A�kBX�N1�I�Df������죃��scIpF�h��<.�݂e"���(�嗛 ����䥫�˙D���M�C���ox�І�0K�q%�Cd_�$��ѯ�7J]hsb�N��R3��v�Еu&ͧ� X$o��#e�����7=g��m�_
�>�E?;�/g�?k��Df!D�O|�A��q��R��}��j,6��4ds��4�t�쌆@���S��n�$yaO�+	S�f]ɕN&�TV�T�������
�5KNyw���
��@J�\	�};�N|��U��IdY۩͌2�+��=�q2��f�"0d����^:ڛp^�s9� �IsB�t���z �y\(��;4Q��Tj�o`]�ڠ�[�����؜��6fΚ�6P1l�L
Q�B���w*_3�ER=�[veD�>2I*]l)�o�L�>��vv�-r�X����P�����:��M|.�s�}�B��'C�c��e��ze��P�?�s�ÆC��M��`@���TIz�y�k2�%���"�y���(�&b���t@�W#�i�x�N����eJl���Յ-ma /��<���1�J0�e��o�\����,�U��5�X�$��[�e�Ŝ���W�Ur�M6J�Jp��`Y��1���l'�@f=p���3s(��#Sm^2<�Y	v�C/Z=HeK�����S�P���ˤ �����LZ��=�;�<eoN��VC�L��ҍ��%H�\3t�}o�?����!�m�g����w�J��l�h^�^�Ū6���
��;T����mS�� �B����՞�R5W����:g�u��}��(���O#��Oҭ�y�-K�ئ���	�Luk�VY'9��9� ���� +�����|�[%Ժ=y#<�6:�Ƌ�Z��M�j\ap����TO�L;cq�c��z"�p�TS�J�-��9�~hH81@2���b������}ݍ�cl�.H���u���n����S:sc0H᫥S�T����R~�CZ�}��{�ܺ ή�d|�tVQ��P�WVc����_|�≱<+�{���8q��	���EZ_"�A��σ%S4QV:�&�F���%��N+c��%��ڹ팗����="z���������;��Zgd���:�$�A(��Ȱ��-L[f��X��a^bgnc�HΙI|�.��$��;p�S�Ѹ�Fp����V�0?�q~�Ƣeb:�^c�/��֖~8��q,�B�&�|�~�g	���)y亇� �)"��i���W����_ R���Ux�9��9�)�b��W�0K.T�τ��VI&��@$��ׯQٰ5��,�AT��6������ݠ����k���M�VJ��cl?�7��T�H)]��d��Q����6.[�|Q��J���8B+~p�IS_����KV�r��"�k֚1u �-�V���MD���Ӈ���Z�oys�N!נ:�\Ǘ���^�5���=�f���*�~
��]`�#v���:I 
��":h�B�^�f���IxSw2%��Ի����}��*X����-sR(Y�f����^zg5�#v�O�-4t���?�3D�S2��C���ၯލI}*e�NpX?�]�\k��3D�;%9ƺr5�z�����n2M��O�(�a�4�Ww��7���ӆ2L|1�%m��?MYF��1�|��9��c�%�O9"v��o̝s�8�tJ��x�:��[�)�1��	�3��~H��h3���V���-=���MRy;��A(�m��,�S*��A�,�Fi�gd�j�;�@�����׀´�Z��l  �j��V�-N=��e��q�zn��,��� ��%�uq�̝95�V��v���TF�F�c�{���A�k��ҷG	*�U�/oع�����[ ��S��2n��=$�{��2�ѕv��q߲�b����-{�C	d�eh�f ����X�	ض\E��%ת�"���CI5��V�CC8�{��ɷCe6���%p�S<�z�>�gv߼A�Ks]�8У|���Yp{�P�/�F��mcRr͆h�h�ѫ�'�i�3�M/�e
u�Z	A��;N��2���_�5f
��~|~)���c�r�`��p�o3��"�I>�O�G��L�=��[���H&��إmd3!2Nq��s����~�R��3�KR�X���.ʋ'[!6�ί� �G�����|����n�~M�E���_�VX�c*ܮ�w�v�ܝVv���c��W5ؚ\������=}���5���{���\奶) �J[�Z���u�w��k��z^�b ��%{��V��!��߃�Ӧ0k���s�Sj�[/m�e���W�c���w����/�J�\4疜uI&Av�����!w�����=%�oM�6�B��S��giO�m�a�p��Yo;'\����H@0]C ,���HM���X��K ��W�ږg3;-h��5����=�<UzO%��4�*�焇f'_:È��]apY��{��户��2
�f����}==�����PH�lg�{A���_���cT;Ш�6�+F�����\)F#�5a�d?_5ݹ��ΙͶ���ww��2�>�g���L�V6���0eW�n���3G ���=9�%G�A��p�;����ф�,�{w�@Q��Rˑ�<!����#g��!�ɐ�Ѭk�r�Z�����EK�yN��g��Ցl!ּyf���a}�7��-��e�;�!tXc�#��6�� ���=ܚ.�Wڡ�F�ؓ/�
Yd>4D\�N��p(Q��ŗ��8^�'�a�����a5i���?yef�򆟲6�^L����0�C�t����if�fu	��12_����-�AB*`j�_���t6��]��?�Lnk��7�+�\^J��=1@��P�|�š�=� ���������u���sKzU����D�+ㅥ 0�l�y��m��ˈ�8���x-��T����9�%�p��F?7���{̦�_k��GQm:�&�o�˗��a����o�o�"b-�td0�5��y��p����g�o��`�	�jl�>�}7U	��$j��ѫM���[�I�����зpvV|v��S��� ��t8�
X"Nv��G�(A�W����΃!�����[��;��!�O����(��V� Wxch��$�?��R��<��_�ݕd#��J�����b��� (�̅�8
M>�Mη�ɍ0�}�#;�w wYuk�-�d%�ʞO�$��<'޻�}H�HV h	���&����s�s ���d5;{[
����]�VF�������B��g���YC�P�H�C���ݓQo�:��!&���N��I�Z
y�3�ڡ��S	0� |;�f��X����G��A3�S�{�C����!V��bL-,Z�������J�ƽ.K��+�l�ñ�n�l0�!�������M����/��8�`��#d"��k|EC����RmLC�ϴ:�.�R:����ϥ�{��A	kwB_A�Z��
�.��_�X�?�#J�2y 2Fo�vFP��a����ּt�ɭȡ�E�ח�3w�3�,���&R��zh��#�*�b�<Jt<���(� b9�̾���m;�:Ȱ�p��J��r��aR7�F����ă>B7w�_1ZJ'�z�[�XUv���<脌B����Гšq�6�z�X��)2�����F�KN�ۤ88��Iqwtp��l�[���L�Q�{GIw�tr����n)Դ�݁���u����R�������t%������N��"�~y^�z[���G��<�sԕ����|H�B���m��@���|���r�QA5N	��
o����ۇ1��G,0�ٌfw�˧5�Ϧ��T� ���cD�?6(J��M�H��iт9���{.�vTuM-9�.>�+J�Z�Hb�]~�##�c�ϣ��~
L���p�͍�prX�ăY��]�D��Ó=���3�����Z�e�='����&v #��һt�qᝦ��KB�қz�p���NP��Т#���YW�ѽ}&2x��`��x�f�6�K�%8��Y*�Ɔ��}�j�X֡CHx/'7_�dkNT��ND]���t��`rT ����9��oM�"�H��c�����QѠ�,��+¥0(������]��\bl}�Y�:Db4���8�")p/�d��߲֩�%�ݞ�L�~U�"2wF.�b�:C�
�$�vw49�z�c����JF��t���ߡ����o�~��2�)4� � �9�>�gC	��4��3��"����U�o��I.z8֨0���F*��6�zB5ǝ\�F^�?��F�K�a���͚ᒀ�8+��숦������>n�XL����1�<j������WЖ5�&�����Xj?բ�wkS%��a6�m�{�4�,�l����䲐OAw���5�ʍ�Ɉ�(�@@�EMB"�|���n��$4g��Y��^�$c}P*�7�v83�޻�ŞO��nqa�zni\�A�?�A���{���!j| m�����N8Y�P4'ОZT�퇼|�{^�6U�c�Q��H�PjI����Kp��T�|b�W�����-)��G�����`�Ƚ��[$�ݎR��N���flm�?�aN��p/%=Y������'^c�M�"{'����%+�E�f8*�'�үbjǝ�e�4����2ti�?_��?��(�y��
쭗?w�!Ⱥm5@�chLy����G���wO򌢳E/t)�{H��n兌�*e��GC�@$Ll��V7���7X�~w�onU�&�*4�u_(w50 �(�)����eeW�I�M���?JP�]�:K���@�;&O�H��3I�챇�0$۫�����
�c�L�W(jʌ ��e� �]���a@T//�a�q���"2���ypv��"��?���:�%M�`
2/���14-59��vr[K�*Z<x�	���ϸ�#
�����z"(���k$�=��ܢ[E� ����4��Lk�Ȱ��x.�Y�;k�kˊ��qO�>g`ȅ%7�Ny��l�_�Ӭ�^��	�"��#�]I��\W(��m�[��˵�{�^��ru��d �$I:�Z��lv�y�s���������ե�C^r�T�Nb����\K�!�x���&�3z��2|���nî
v�0��fA�hl�0�F�{c�)h`���֔���y+oZ"vX�(�_MǔݹƔ�ǟb$�2���ƻ��>d~F��H�-�2�*� M�;�(��$�F�C��P�+�� �N�FN�5?�~ܷ��w���l���l�8F��u�fׂpea�jw�A����<]q���ڡX�A?:W�
҃}b��۪�˭�̥'�rgb>���
Z�Sn.,�ɹ���/Ȭo-�i|w��>�>aF��6DG,����i.]�u��Sɩ*���Ȗ�jCS}R��u�r*�a�������h�>v�]H��N�k!�9�EŒ�]��jĳ��C�"t!�#>.�c���(S��?�./�PԞ���I/���͹Y�-"�n�� m�@Q#?f/$�kzc�_����47 f+E��� ?��m�֋�����l:7�@nj9�⚚ g��t�F�/7͸-��"���̌�hH6Uc����~g�L��:~%p�\���7�-�HNe�k6¡��d.�����l隝���.���uy�T͉�7%����&���@������,R}V��َ��~�ب=���"�LE����0P-k�>�� 6�9�&1{����b��˕��ēۋ#h���V�<䋀�=!Yt���}Rei辊���$��x�0�\�͸�"��ᗥ#nA����pV��'�߸[�+_,#�ƕ�4J���#HM�nF�9$��;d�K�CJ���_t3�ױZ��`?�̔�a|t��&���i9L �J;��ɫ*�|����պT$-�%���6%���3�T �xo�^ u�쿘@f�Up����w �2Q�E_	��d�숥�N0.�i��P�/��f�k���M�ΞlL�2ݓg� ��a�-&���0��i�+wu�M���c�A]I�vQq
�i��j�ѹ@��/���c#ߴP��հu\�)_�ڠ>U��-GO�Z(/+�YTc��tQx�w"�1¿�F|�>�~o����67�-�����9X�ˢ�	Rk����I�횢L����hf��R�a�_���~j���ze���)��(4���mK��7$	&��.�|Y�bY�U��е!���DL`@g�"F���=�y��ǃxl�#}e�:\r���YP��#�����zU�t�?����3� RS�>��nL��0�\����� I��4���^D��:P�][�}F����QTbl�ȸz��p�1�Q��Z���K	k{�q�aeQ�� 6��y'�L"��)gb����i��!B)�L���10����0Vᱯ��5����g�M_k�]�F�\B�;�:h�V�ᵙ8���d�'�bٟ��ô��M���7!>��tA�ް����NЄ�UNQ��!8�W�,#��N�W �S���*��@���Tk�ȶS�k$��.}1�$j�=�s�qK�b�ڦ&2Ź�Ѵ�9q$c����nd%	��ӵ��Ͽ :�kd����V�<�ݧ!�T��c�7㰇���;'�(anX�F��_x8�L���O��׆��Ʊ�8� ���f�&�i�A�#d�Q�� �Q�YUBA�*j�ωr��4�8�v�8k�_����\�����a`�=C_K&Ƕ0."#��$®���$&�ے�>|� �J�IU��5K|��p�L)S� ��-���;[m3��TS��K�
!_Rf�q�/��Ȋ!3��zAJ�����d�IӨ�sK��p�jG�̞H���ԛv�R�m�{:���˅C���.�H����8����R�ơV�\���XJ�"��en�fq�m�榭w���z?8Gg,��~��y���h	�h;&��������gp�Pe4#'m4�!x=��sQ@�VDN���F��pr��I$sB��h��txn<�?����xޡNQ���~�u��� ���"�0(��{?*�Ã@�S�X//��r�%�L/e���+�m^��sw��	(������p����+*��
C�OoǶ��:3ښ ~v�*�3<c]"��I�1|��ilrZy�2QWn����ϻV6~����O�slW�z`Sߗe0��_C{s��R�𓙱���*ޓQ>�.��CB�,M��i��[-�!��_�[!��� 68�H�hL��#�}�[�Z)�J/1�e��f�p|�CL�]�#�E�]�΀F�.�S��sb�)}�j-�����N,��fD�|����8;�*����5:�.Ѹnky$SV�.�χ�r/Y�����D�/�mj�h*�>f�۬���`J�>zqV����j����"�W����UW���: `�|�$�//�Gb��F'ƵJ�o�>ܧP�!v�o$!d���ƈN_
��g��(4�A��4.���G�n�rr�M�F��hS�u#���Q�I���DWh����\J��:(  ��%7�9^��'K�N�	��@G&�NZ)P;��)�q���u����H��A���D�]�-r��`�w`�x#%�Dc��5v��9��4���]�����򉂣��&8U�F�_Z۔>J�)/,���y��ؘ	G�oc�fjnu3��z�l۝�Y�B	��K5&}ցu&��$�qEĥ���'���?�H\�{�ͤ9ȩ��l\�z7B��7���l��(�t�֖���|�v}mЫ�L���c��{�Z�pGS��^釺%��~�+-f���y�9|�ꫂ_���OL�e�9�S��,u���J��ᒰ��ĉ�mT�jt%x�&�~�9�O k�˗ȑ�=?��ը�D������" �}G�$yqm�����|�\��s��q0����5�:�y.�t��ޠ��2wTEe3	��|Dv�d/r�|T�K����0��[��ڱ�sq|�,g`O��w���D�:חy��&qw;yS�gޱ�L�����N�\������#XLb�a��� �*CWwF������q�[��Q��L��H�Rj�UKϿuv5�^��]�Ίf�]�PݡK����Et�.{8s��3�o�림��uw��e���O+����"Nd��0t��2���Iy����:S���o��j)�
k�_K�Z�`�O� I�:|��	�$p��\�}���M)�rL���P���^��>���	��:��u|��v�9W_�
��)�r�ɖ�4Dj�ۋ�j�˻���`K�bř.T�4[ �_��w�Nx�$����sn+�H�L���k[P4_x:bB/��׵;B�ߚ���j_QU�n׍�q�k�}�2�=�̫j��\��eV�Q��5��L�⚘|N�K-UO���+�|v1k�T~��r�^$#�=)��fo���^h�XO��WG<�I����;��st���B�P��k3�ܔ!��Y��݌���U]U�I�����>dA&������LDm<�\��'��c��!�b���>�ZF�w�	�)��6ӺA�2R���	�Ekݧ3=--1p�rr4}�R3�6��r��V:���pr�8�2IJ�D�V�6����)qLTP��`��F�Dei���ƻ�Q�jVZ��]�Y��x�t�2TeZf�(xT׫�9���Ń���F��"4%y���	z�g�DT/C_�'��5>�v3��qA�疫�<R�������u���~#*ݼ�"�&y��>SNoꗨ�)�pS�QN�.zE?�LO/E���2������(�*��7��kd �J��xyf)$�~�]�.(S�&!�휻��l�P:�oDRi"�W�Xл;��+��������~.��yN�n�^��f"�Kw]J;$ks����~�Y��lW��(�_�I�A4����&��3n��Z��Cb�w��X�D
�8�B������݄�B��^��j��-�a�*����Q���v´�~ӟ0Vϸ�f�ִb5�]�)�W�q���؜�6zߏ�'E�n=th�!uO�51�\z��+BA�7A�Q�b�P�I����?'|�������)�p%K���5�2�� �C��$���]D�F����O�g�s��'t>�C���������$�X� �!���E	.�YC��|�tBiX1#;��ۯ��he�Y�:Go���>���z�����J�-�3��M����j�@nCs%����'t��,���1r����Ѐ��G��� �9��7����Nڟ�
g��9֊<��}}��P,�.b���n=��A�MRsUi?���9��c-����N��C��F.��y�\�Lc�&��i�m��(dT{T�D{q����6�z@r��͛n7���%E)Q ���R� ieR.�s*���g�F�H!���qAy�{;��5����/�ybtP΂f`z�'����I¤���>\�%3��|0"��Xܠo��}�*EPE����	�1FZ��2��˅��Ӹp5*pU����U�҂�.ĔqDl�ҽw�q�������_��npyV����^x@�q����ȿ}���p��S髮�G�
���g�ܱ8�t�+�ϭA���1�L�FPv�s<�9�g�V�a?L{ ��cQ�f5������$z>J7����րs�$���8��?j}�{�l�"��,Q�	��A�5���v1R~�������j���_I��Hm�.$���XU�X��:)�j�,&��Y=�NH:9t����)���B��������5j�ezR9Q��p)�Ѳ�e?d ����򝬲��,-�ə�滐^R��3���z+�ᑣ�*ڤ.��~[sߋh7K���g)?���D)�oI��V�+��d�ţ��TǾ �|q
'z@mKz,ŧ�����nw>3Hb[�3�D���o?�H-���*5]��q�"�B�>�0-p,ᵔ��հ�ӗ=�¨n��5��I#��������:��|�a�"s�GD/f(�ӆy��z���"��Uh�áa��Ncp��TSU��������TKV�� ���Xp�B��6��N]�0CiN.x�6ЖW��S�ŏ'1aF@�����D����={7f�h� I�a�r�$��c��Zij�n�	�#�%ϐg/i�r�袊G�O]�^⏞OTM������}_:�ό􆗘��Pσܿf3��p1�ֲ^`.X�tZ���@0e��:.i!&�-4�� 5�z(��=�:E<����nc�.���DM�w˞��G��?B]w���۳�����)�wW�%�q�N�gP�;ɰ[ _[��ɦ0KT�S��.h��ں�,CZ��i�k����������	�(+����/JKɇ��V�jr*88Q/ӕ��&7��-W�s�w� ����%��!�:�<%c�W\_c(��2����H_��cB5���b�8ց���)��I�o�'b ��IdIN�����_8���%��7�9Ef�p�E%R�0s����C��#c�E0�l�F���²O�Y���_����h��$q�k:��C����@�x�ڨt-Y���u�BԨV��埌�[3Ty]��cBrZ�28�f6oi�-�m����� ��Đ��x��널�P�Pz,3�園1 ��I�Q��m��& �6~�>Paփ�p伤D�w���%B� ����7��1:��ڀ����ss6��,�a�:���C�H?�@� �ST����`��� Rq�c��� �Z�'�`d1��{t���ʖ���P�����6<KE��¨�w��I/0m�NRi,�����U�T��tI��ccw��PV]��e��P�E�	��iS�����I��L��E���r��h"*RK ��L��	��� !KB�	*�M���r�5lv ������A{�����jXܾ�S�ڢq��A	W����c��Q^-EE���vu�1���ǵo�H�X�w�"R�0�wax�ǫ�mr��;��+�j�˦v�����(9���ڄ�㟞�Y�Y��������6#���7��.{,Ͽ�q�Np�w�|��_.
�;X��:��M�HH ��@�7G~�����;5���rW��S����w�!)d׀e�%����h�{2>k6�w����v$5�����N��9�kPf���<�_�
W�!}�pG��w����5*!��̺2:�������G�	5CGfq0
�?et�.��J��a1�:ƫ@ѥ_�B)A|"�/83e2������p�,�*�� �)1��R,�~(]f�/�� ��|�#T�v�Kwl�f�l����q	��Kz�����t�w����MC�#@Ǥ?������+��ށ�{�ͫt��<v��a�2k������O���ve�R�^�D�㧿��3ֱ�P�-�^ӂN�����p/��d���m���?��<����zʷoOƇ�[P�0�Q��}��l��І�VQ𗪛W���ح��h�!c�k5G�Yab���UD<��,��+�|� � &�F?�햖�*�K�Ҩ��J*�c(lWX/��)7Бe7����؜���4�|l�{������8�#o	���������9˽�y��'�\;��yȓ����6�X����_?�L�RH���1U�$P�N�eE���7���5�0f��qj�I���H���-����k�s���s6՞�wE��-z�� ����*��qЛQj�hZK����Z:�!{;�s�x?O��"�$�q��'4���;��gف+S�������!"&W�1�+��ۙ��������υ�(���D��A�+NT6g�GL�_�7ɰ?,�}��8�N�0|hI`����Q�gwPi�<{hYM����nS�O�R>˿{c�f.�+C�׏���[E�6\9��?Y�S���猸8����y��έ]@u`���IL��%�%��$J���6m����,�/���/�4:�t��leaD��Q��')�ꀄ��ڴ��I��X��U�g]&���M^�>����G5�G��[(u�����;��������wMj�6���|�riZ���l���	����.��w��uPU�2�k*��s�~r3���h�gզ6w�e� ˡ?�P�.�_5?%nkUd�50dK�_���G%�0ҟh7�y��@|rhO�	�����Q~���s(�v9�|�3U����zl>H�K��u5b������A�H ��	��' J���.�����]�4�'�=� ����-�ؕ��E�o�UԈv7���#���E|N	�`7��c��guf)!}ġm�6�`Z�"![�+�m�S]�!%��>\e��N���l�+��l҃;��#(7�7Sd�����*c[��?�~�m+m����&Ae/5�7tI�:��{�/+"��ʮ���^���4]G<
z%�b����1��p/�a�c�z�G=I�X ��w��4���x�6��!�#j��޼0��9����`$�������e�O��]����5g�k�ڥܫ$t��>��,�Z�B~��!�i�#4����F�ya�f���-ߊ?#�bߠ$U:O��2߻���:�D%<]��� o9(#��4x�(��s>JG;�M���;�'LX�P�X�_�ɊN~6kZ���<��6y!k��\Q1�pG$(���{¶�47���
�kڲ��lP���:F��Z������h�,�w���*�8�k���.~q����z��3w���.��XL�*�:��l4}!r`Q��p�͎�n�A��o@���] Gk�V�S!U�"�3�6~�П�*J���@Ȗ���J<�	,P ������{$�G������Q_�I�ɝ3)��ʳ�R<-��*'ٽ`���<��<T�=��&9��������C��������L[���M#��}������7�j��t���y��S��!W�UqF/d�%�U=a�ւD��+���7�>0�&��G#v��}
 _E�l��:��>�C����ؼ�=_g@�祷J��wsө|I�f��t�Q�M���6�y/�C;n��R���e�Jo]���6M�Ơ�}��a��I<@��0���߲U�= �<�,�C���	�rh��&�KC0�#F��k�=1�>!i���� GC�����K'���Np�h�����Z���f�>ɮ�!�
�_u�?P��r��'E���C7Q��p�*Z���q����ZKN��:uկ��BI�;d�5����@�Sjq��U�=�	�����>��d�Z  $����f���/�4K�b��Ȧ���KN� ��X!��B��h�t�CX8���LO�lm��8�[ڎ/o��擃_�P���p��j�R�0pCV+4#:�)����-��-m؍�rz�Έ9-?!��\�'vg���@0�xMT2P}�dEn�u4F��cu1�G��lEȲ��s4���-d�M-A{�m����������*q�n�S�Z��� ���7����ƤC��~2����^P��m-��
�m�E�w��@[o��?I���/ s`~3g���i���g|Vxߎ�N79�wzߦ�!l�x�ˡ���P��/�#\EӴ�&R"�ic��q`��%����O����=i���M�`U�N�o�rNd6F�c�$l����7�з��g���e��SM�eP���Ɠ=y�]��<XTx��@k�;���n�Uސ}��?f����x�Wmc�2A��a+�%��#NgW��v��ͅU��!�]��ifTw�������~É��{���})�w�(�cPq����3ŝDW�D]��7G���RŁc_�]�X�S�u�[+����pwF�ʟ��B��kTa�u��=�����������8���%۱���&��Qh����S�;	`�����X�XFW�����8��'>�VSq��ޟ��;�F����6�����J5Ҫ9*GF5�[t䲯Z�}��0�;X�MZ��-���ҼzW-;[��^~J�=0�sG���!������\=|S��U"�u�KDW����7dG.����h� ��]Rj��j��h�L��g�������DI0)V4��ٝ4dO�`��<4��,�2:�rF[т�{�����§�M�Ƙ"�ci��7r�-�r�q��eX�r�%�(��aj��7s=����G����}QX���y�����s9��Τ,�F�'/�&)0�*��۠��24X���T�*$�]]$�.��̧m�����L��9�tm:	��ܳ��ՁTvA��0:��'�#�Y}�$ԏ�!U5�	���Q��(o/xa|K	�CF%'/��YcRQ����j�D����g���6 }omh�C1��ȸ�]
:.|�մĢ��ܒx#e��yl��n[#w�H���f"33����Z�X�F��r��z����,�����H:�S��소���1����8i|ω�+%Ŵ�2n2������\Ab[�+@��l14.q	ϔ��b�~"�=Y�㳟	���ɸg3p����^k�=	_V��-2λOM_�V-Ϊ���G�uw��lFs�p��M}�{֣9�dW�����'�Rcύ��[����<�k�/�&\:��%�U�X�s�ī��B�}h�\�d,� ^�z�ac��I0p�� �zL 
�A��4��*��]���g�G��8~܉M��뒬��>��⇼'p�m�`�

'���O6�(��|&Mh��.?L�#��7%C��_�5���@%.�s&��'G�e�Gl�r�j�a{N��}��9]֦3~�]'sk��gW`>�EZ"�>��������b
[����7X�0�Vzs��֍��`?��,�����s���僙44^Y�`�ery��vE�n�!��4�V�x\��ka�ȵZ����C� ���ǵ*`��)'�J�Uܟ�Ư3g�X�%ꛎ:hl�Z��s�2}P�wڦ�i0�c�Su�aT�m��:�&��8��4�����XY �Rj�ek�&��R&M(��{`�S�dp�0n��;@?ߊƦ�I^'-�Z����r_"TV���/Yyś�h88�Ҋ-��/�g�k��
F��O���|����๊+GjK���A�;>��.Az�uyyTt��ҟ���lY�i��[��]�PX�w��>A�Bol��E[��X��=Y?��R-r�J3�35�h���E�a]ۂn�%����M��I�j0ؚ�W1U�d"|7��%�����d�8���V��"�ެy�\�硭Tu+ER3D�IT���T�2�b>���a�	Zt�Zg���Z�J�F�@�4|����Ҙ�19��aQK�#���o`�\�	�j͍֧(�{����;��7�K���rBY�圯R�މ�����h�p��*���	���l	��-|\��q�m��T�0����4]B�HȦ� s�[ù�5������[Lb�ܐ@.�ղ��ɖQ�� ٧F�������o^�w��{3>c�ŵ����C�uA���}��jEh�Y���/K��^�T��!L�#���2��y��n�P�O��7��La�3_xm�i�1d���$�x`� \�����k���$�����c���%���9�k�Ç�x/�5�.q]�/a��6� ��rV��/�()�V�U��sK��컖�&R3?�$+���"�ߒ�n��΃�y�v�N�kɪ�{�Y�B$���Z��DG:�T��1YX�ݻ�o��i���$A�$�:���=y�7lm��&����u��8/zY�%|�ȊJ��=��]J����sߌJq~7Cn�:���2��][יO�Ӧ"]OU:��� ��O� &��Ka�׾]Cͽ_��`���q���R`'^��o՝g�>R���=��'D3����^�:���Ʉ�Ǯlk�Ei��������-�/��V��qW36��g'��6z���:#{u�}!�F�u��UY�vN��+�bZ��~_-]��C=��4d��G��1�!_J�}o^����"U#�������J�����<J���^#*���8�2�A�m<�Xe���qɕ��&�ZL>X�����\�90 E5�[��94��ٔzx�Pu]J�d��}\o���h�>7���G�~�
D�S*-�/��ɩtf͛+�P����aIW�If���h	r�x�[�@F����0�ζXU<� �O�1h��~Dֽ�������)��J�Cĥf�ŗw���Q��m��$�j�?�B���]���Q��R`}��{ncX�t|	�mO��"ew{�I4��;���� �AK;���Y�7�oX�q���:�J.����G~:���
�-����z.k"��z�^5HB�����jޙ�\���/;���uY	)b�LGi�����cC[W���<����}Z$���T6��f����Z3o|�Bq�!U�jM��)'������X���9�T���ח���(���{m�J*Fp��9��D�qƆ�a(%;��er��g���Q��j�E��Q5`�M�-���]��녀����M��p��5 �6Ln2�l��L�ڻ��̨
��=���?�
�$��G�/5�U���Jd�0ꦌz�տ�UR/�_�	Lw�[��[�Z�p��>��	:�J~����>5^�1vЊ��92ٗ2J�t�7��NPL5�K��{���k�x��o��'��F���s���$i���ԁn<��E�f���;{�z�kJ21+�FaOV�M.W[A%a���e�|�=Z�������2)�4a-�F�/�0������fH���Z� ]u�`�������!���Ju5n���XsU���""m2f1��p�]�͙M��\�/��EYY[��#���1>����g��a���|G!�0��M��5�??��<Q~d���z��z��Nͅآ���մ�y+d��*d�88˱����́_4'���٦�m�Rm�k����A�^�0�b���w�s��7�e�d^Ӕ�VΌF�[a�˘h2f�{h�ȦU��j,Њr8_;ɪ���Mޠ
��u~�fcʢ�EMD�{��m:���0ª�ػ��hD~���"}X�}|�[����ͭ�������=3��9tD
O��
��$ى��=���+���3D8�;Y�E��jj�L����:B�u��Bѭd��;R޽���1u	4'�f�<[����2ѱ�
��Q�I�S����n=����x\[�Y6C���q�5+�6��ǒ�� ��� ֲO,���ZOO�w���-�3j0�ic,�9hm������XH.��BY�&.�.ʐPg.ۛfyW�]p����}:Ϊli�'�(Qr*����O�OO^#�?��]�����n��Y	wL��^�����o�,E���[��tD��W@kb����Ь>�ނ�1wW��hTy�0�/��1�	{K|��K���t��>j�N��	��A����Ւ�?���&��&�B�m�Vq9;E�D��D��4QPO�X�V'���ڶ���B�x�
֊Ne��D-'�~\{h^\�3�;{����?P��&|hb�����n37�!>x������f@��A�m�d\GMa��聳b�z�쒤Uޢ���~�ݵ�u�ނ���!�=V���=�fP������|R5��h��j��l�?�Z��g���f-n�W�*��2Dh�`�fww��s�/�5��x�Z�~���66ŵ�(̐Z�gw��m�������0
[8��y���Y��>��z�Y+�b1��4����c��Ou9mBa�>������`?䫝M�cQ�V���"G)�F����&��cls#�p����z���6�S�3K���g�GF��,e��!:����1��K��7J� ~�S�ӟS	�����w�.�}�3��p	�A�$��s���֚W笡Ջ��)vb>?��?���:�5쵿��C��i�θ��=t���Xm��ٕ�6������*����1���7Gۀ��X����8���\�$:���f��Ñ7Qb��Fr#f��Jj=PtJ֖U�a�x� �����"�|Wlɨ��);�i��z�&�E��n����+b��c��%T��ʅQv�t+	�j4ux_�ʸO\�11�ԧY}���y�\(��s�Ϳ[V�Sպ���s��-,%I%������ka�~{��� �5��}���	?�5�.�l�5�'�5��j�����j�Vn��X���G���iǖ% N@�-g0C�[������z��t:�/r}�uL�g�������鮓.҄s%��k+�'���z�N��	�,`�ۍ��Yv������[j��M��,17����_��7�~ak��#��fr��`1�I�Č]�j�l��?����z�B��L��;w���Ǚ.WjC�M�]��{�l��3�G]�r����JU|�� ���0�C��ĩ�G@�{u�J&��tN|�'�yr!a��A\D>?�b��<,kC@
"e�Fm����i� !�4w���x�=����V��m�����Qy�,;���J�CC�f��:�3r`�p`�Z�|WH�N�������"�ć<:h���(�B�\�{���c�l\�ȘW�o.�����>��ZP��w��04�rN���VdS�+�}�Y�˲�[� ��$�w ���hN�#�dЩ����<�z�!�a��W��wbRe'g�_1S58�?	�7Q,91Z��1K�y��q������S�d����#R�[&(��+蟔�v�L���Sg`���Զ���1�S�L,����W[v7m?�B��Y�!F904�M�[I�
t����)��ii�J�Zi>b�-��{?[�^�rX�"��w�f|��B���Ѥ�BS�G��f2�|K�T�6�d�0B6��rfɍ	�k`��I*�§+WR�����N��FĶ+G4t��ԃp�xV�BO��P��wp瞧Ft�T.�0��u�*�A�A��y�w�����R�%�����s��2��sW� �]��n�H��WCy I��!����m:;>�_�Qεq�HL��ű%�S�a���r	��G
��n�h�?�-h�s��[�'��j#�!țǡbn���� �~n��Sر���ߜ��,J�8�Ih{��QÆ%lO��B,bC�����4$L}��^.�Ԧ��z)=yU������!��F�Ր
�=5.3��;`"���-���8V3�F���-��wY�-�X��`�˘�h@{ׁlG�A�g�0 U��0�ȵ��H����iO��
O��O�k�x4��������+��	܂��h��N k���Q�ث�D��Rÿ�J3B��!v�-�1:�4lr�� \c��О�ЏE�
L��b�w��`�Tɺ��R_A��^5d����G�����a�6�YHEq����5L������>�Ja�k0:��T�J�y��d���W3���i�t��G����X��0����XݪV�r�z̉�$d"�H"�/�p9t$�P�ﺴ�ß��(x�8\��4�)p!�1������R󇇹ʄ�,�Y;�u����]��s�l�\hŷ��L�m%d�6����mwPO�+T4��RPU-��O(K't� W+E@C'0�bԝ��\�>����/�B��{mA�$���^��F[�-kGm��A+�NlV�%=�.�$�J�Ii�Q�f�g[�y���;���_�ME�؝�F��������j\���\��L
�y��*���:F"0�H�h�f�W�'��q`p�3� �y�C������W�I��0]�&&�C4F)ʐنyL_5I�J�ڏ��G�&3i���p�W��C{��O�Sס�՞�X	�c@@���>�	l.^-r�WVda<p�)ˎQ�Uo4C7�y����x��t��?��|\��r�ɰ���8�;h� /6[�����b���O/�.P$2J�_}����+�]X{�wxW]ɣ\�kK���Zs� k�rw���{Y��S��Zcd	F���=0���<�(�IW�!�|e1;�M�DAG���\J�$��>�)TRE~��31�"ɕ.&�N�f����,�����e���#+�����;���)�ֲ���
�j!� �7�9j�F���0�^���������u��?ߧ+u/>S[��1E���=��Х�ص���.-V�ABP�\`�w�E�,�����k������I���bB� T�ft=�?�i�L�f u�Q+Ku��Rn�Ȝ��\H�(��45A)��[�A$n��y���1Qp��.5�j��@��웡�l����G5Af��\��E�ں�ǘbX���*� ��[�{�.���y���=�NU��U0�� ��4��<c����ĀZnr;���f%sI�14��`D|�����r�Z�D��U�ߜ���kң�jdW�Յ��Y�h�d����\**���m٥��h)�u�pui,����|����S�M#�N�Ε���z�Jd�J.�̚���f�>�:���+�S�<�ѝi�`蹄��F+�b��P��Z��l�J��/��~�uj�B!e�~S�B�#3��$(��0ERX�4H2DW�%Ǳ^Ŝ�`?2+\��~1�����w_MQ�@4m5��t���/�Ix*{A�0Gʮ�������F�����M�_��SQ��^U�s&	T��ړ.~w�����R���^Յ���}����TQ�q,�G���Kx����;h $� �Ⱥ>c�=�gU@=s]��_�D����&�I��V�ۨ�8��7쪆jw:SpGL\NB�� �/��:���V�Z�؊j�jg�
h�����f&0���N5^̭�=�zN�Wd�!��+�Qv���n�,_�ΐ;���vϟy����)��)ӂ3���Xㄥ?�R��O���h.)��J��Y�-���v�[[�]�P�c�Gs�G=��E�m"�}�&��Y܊m�ۥ�/�hϟ���*1ϋ���|���e���3F��zyr��<�Ƞԭ�zd[�ESK���rYۜ�Dn}մ�zU�0�����S�IY,�A����1tm��D+9�\�G����~:�)bh�iu�9s�E���`c�����AA"'�:�I[��|��v�+�kX��p�\:�e���(�˚){-v0lq<�	���X�jl�28����0����_��E���,
�(x���j��rE嫬�"*=��GA�uit��C��CV��m�yS��x��Njꋆ�/(0o��v쬗�B��G�+��-��{Q�g�əQ�AG�	���~y�/�2�K��k���\�,D�َ�/g�Y it¹.8:���66�Q��S��R#�9210�^#�7����re�<�Y��H�����Sj���s�>�#�V���x�Ln��7}�	�'+��?>��̀��o����<K��ku��V�¨}]<�0
 �0~D޻v��s�O�;����n-���QŦV�߆�>u0��G���7�h�y�{%.h��(n�c�!��K�ۡ���r�]�u�U�����#���#���qz��ش��A��n5�dU���X����#�/��n��ßЁ]�_���� 0uQ�j���ə��\�����]���q��Ay��>��}�;e���DXp(�a3����ʱ��PE��ca��a�kp��D9���"m/�?<����)�cZ5o��h�����8��_`�sy���i����2�G���"�D�z+4�8�a�eW6$�Ղ->=64PY�<O%�6H Jp������ĸ6)4��Z���p���Eч�tC�b�Br���:���{
���&��!Ŀ�#�b�b��Dw=f j9 h��v8eqX�I��z@H�6fJ"!��E�Ңcbd�U�C?\(ťl%1��)ߛ 1잠�;�tW���A�'���eeE2{C��,&���HF��[(7VuL��gF͜t��~�ҋ~I�8�9��
��Y�1B����Fw,xCv��Qʜ��eV.959#�����yxI��5��ѱ�x�`G�yB�,pJ��9HH)f3㦱�D�<�7Q�|�J��\�9��?f5�S��ٓy����t{ي�{�](�xsEct?ۧK�2zל��\at�폈G�g�ѝaT���I�T������K�����15/Xo؁��������ƴe��x��x&W�&�:��[�O�i϶~P��}~'&�E�W��
�q[{�V��ö�G}7�:Ѫ.�g^V^���N���a��QJ>�~i�KY�L������i[��;�J���[8C�,?rqh�{���"ԖHI('�q�7e]�q�����۷���b$l�Y<
c���~��uK$C��p��&� �Û�"c>$�ZT��F������a:͟�Bt�- �D��,����T^,4�������Y0k2��Gϻ]�j��5��Uc��K�~�)7zhjr��:�&��T���J�!~]�r�[Y����O�Sݖo/�j�g��;��7���C�k�����@�^�������3N16���v�s�c����iâ[0�!�5~Z6.B���0?%��7�Ȥ�7]UkR���a�ĲD��W%9�vF�|V���{�w���j��$��UjiT�[P�p��Y�h/rO�,����\�ّ���^��3� 4҈��KE(����7fPV��5��_��ҭ��%ڍ^�D��������$���8�e3}!ste��t?��d���|�Vi���P�S��A��	Hi �>؁GOY�F�M.�NNp.}�s��*~)��i@(��kP"ت��=��w��a���?�Q���/� ���}�����$�Y�S�کO��j`
�k�Ȣ�uE�Z6I�W��v��^�gU�s)!�a�,MS������`+�Ca��5�G��˾zmV��/(����1|�اE���iO��:Q�6��Ӵ�> �Qw�oا��%��G�U�&�UU���`��:RLSZ���I�V�@���5�6qf\��<1�R�{���@�\�mp0�Җ#� ��`�*�.ݷ��@`� `����>]�'�s{QKԃ��I���%�;���9��xi�qob���j���q��Bs^;�r��3뙤�Hi�y'�(�5�������G�<>��[K�B� �{���u���@�?_#&"u�k����@���F�:�]#%�[�Bp�pŲg�c�	#��F�hܟa��	��,f�1�5e����5W�:����[ �c@rpSP�cF�8N���\�+�X�qi���x�`�������&.�d|������B��<�7���*�Xi��+Ǽh�3VS]���b�޹g���t��gW�'\j�.�H��r��9���r�X��9šXȷ ���e.`�'c\�	�%!׏(�����:+q�_qi������<E�C��Wʛ�-��A��OA�B���z�´^�c���^l���D�]�F�;C�S�↞yE�������=��*�Ct���gK��f���E�	�uG�l�y�NY2Gx����O�4�2>�V�y�n����n�d-�DU�a#}4��*S:[��)g�+����C��Jk8�����ة�%����{n ��G,��!u���#�u�$i�a�L2T�״łu';	̈́�����;t�g�#1������q옐5f�(*����E��*GB�R��T�v���H75�Ű0��tY��^��W<~�����|)k�x10`!�9-x��!`���M���#��ɏ��W��l��J�on�ȣ	3��4L\�
y�C�q���<��І���~����܋��W ���3�J���`XOݎΘ%�80�pwm|r�S����(�ǝ��9$Dܺ;{�)ўq6U��HrP�J(aPJ]h
�a3n� ��N0>����
��"���k�4������8*��V��/ژH��á;͢�\Dm�bq�^���4�.��C!��@���s�S���4��T0�̖��7�]�W~<t��ݘ.�\�}��7�,%�����@��'���#՞qB|�;�b"��a��ڝ+6���/>]��� 8CC�KU�ׅ�rEqz\&�N�<����"���*�o�D�k���_q��f�;J��l*y�1v~
q���XK_pr��������6&c;EX�K�{�J;�.���S�B�O۝��I�!@����xcz��������ၗ"P9v+k���:8�[�p�Z;(����9bs�WlW`E���u���5�[��"��zP�A��W�fҟ5W�7)��@�Ϯ���˓"h	8)��:�2�y�3��/�OȲ���^ѕ;��gc��C-�K���(�~mp<�{&6�YF�8�Ŗ]݇[�L����AKJ2
�r��d*nݑ���;h_U�:�	�(�X�/�+��9ά����S[`~k;��3���%��r#�K�=��%��@&���Ss��%}��H��r���'�'��oV�1�]ޖ�[2�iB�(sW�<8���Nb�G�E]�DKt�k���96w?�sC�3�����+�j`�v�ֹ4�D�1GuY��:���
��x1?�Ƿc�d�x1j G���P0 284����;�$��Vȿ {+�(��p9ԋ�
T[�-B�[(�qZ�s�QZ�!�\9�z�5D�����`m30���=�z�?^(w�'[�z����D�Cs�u��uNh���K�.��8���<v�Qi�c8Z

2kj���x�֒G�1�)�B�R�4�Pj�4���5О��YA��y�*B�l:��*���0w�@��ve@y�TB�����ɷ�T!�V�d�i�u�G��a�ұK�C6��d2�E�.�y����B��#�Aj:�x��e����7�i���z�@�M���#����G�+���l��$܇��4e]ע�,\p�
=��A�j/��U��=p�o!�ܘBj���;�Ej�B���a����ň��w�X |y�����M�W1)A�R��*(]��8o�a�=�PM�< �sM���c��[p�z��ߛ�#<�Gj�.p�eT����B�H�^��7G�`�4=���u+㾰�Z����Y៎�Ug��xB$�B/=ٱ_e-�tӑ�?le�I9
H�>~�M*���a��_�5n�)JD�.��Y���@B���S�op��BvydDA��+�_�/�BN�n�_eΐ�Un ��O�~�dT���h��4�"g�WۊaZ���)mK����ic�ʬ��HM?���R�!��+�q��D��:Ko��\�����r�2e����Z��BO����KҚaxQ�`�)�U/[���Q�XmRυFh�X�W�V3M��q��D� �gvU0m)��� 訏���Ě�����=W�R�g%��s�_3D���������̏�[�t����Ⱦy	C������9�o��tx�(%h�c!P�?_�|E���=UV���?��߷��a�*�&��@a��,X��;���$ID�χ�ᐶs����y"��l��0�-�1y��1Z�|��0x�)�����P���Ĝ`�H�z�"D���6�:��
���/lF;8��q�e�Er�q�f�ľŬuw�9��0D����luv��4C�;����(�ʟ��Z���dݟ~1-��/�r:O��Q��n��=2�0��,_W6�mE��e�^��^�H&�v5Y-��Y8�/��f��Wnl�]0�A޼pC!��:����L
�7���Q���|ڑ!�s����J�%�~�Etq%c�%�(�{�D~T#��M�nb��?E�[��ͷSh��O���1�?�Z��ă�r;Qk4�/b �{}Wg�3������z7�?��$�]3a<Y�J��,��*�r�a����O���8gEtBLʩ���,��+FD���<�j�Q��~k��h�G����2c�=�o9W���(4Tgw�QM}��7q����R�HW��NLc�(=�7���� �N]]���lf޶=q0���c�������wH��{�i�c� �xM��◇}�3�xƗ-S�<Ä�K�@���R�� u�
�nO��1�uҕd^M�)p���]���a��c�O�	�TZט�3)�~�'E�����U��%H
*� �z��:�[QXݸX����R�0ۖ��<>a� [}����g�����"R���VԬ��\}���KAʮ�n�]h��<���׵y�FT�YҪ��ϵ��K��"=fe�9M���@؇A�?bZ}ROD��3��g�h�,�L:y5{H�C6�f�~B�+m�*��;��o,���6Z�ܖz4 o_e��]9�����Z<Y6o�ng��@��ۀ�����>�{�S8���-�_�j��8�+_�Cg?�g3�5{=	l+GC��X�_��9,�6��Ч��_�~����>
��@R�B�n͉(v�=G.n�PCRG9g�̺
�,�+�@ϧ��Jq'&Dw��$��$
%�m��$�V��j�c���l5�|��g-�"մ��\JҦ�sh ��*P�70Zv�MD�����s�ܹ���T���w _�س���.�L��	�u��ƅ�W���1@����W̱���aF���v�AV���y���ud�3��x>�Rg��_Cg�g���2%q��)���ɦ��̀X�X�,���'=�ɸ_W�@Qc�$�9��c��)�.�>3�t�V����Y��4>+<���C�������b�Q�����t�'��s���a�fI�b�Yv�Ѱ�I�."����K�)��<�h���@�)����tɼ���T���:HW�/-����+\��_c����&n <=t);̱���t_�*��kT֛ΖR2�B9	P�|�Eկu�TBq��%�{A/D�&f�)������!�A�8&�$k	�\�1�E��a������1d�1��o���כ����C'4DhC�s���l����ئ
pG�T��0ſ����o�p~����;� ��=R)��l.[���l�փ��Ok�n�ŋ��j>�!����!{n��^��a�%�
(���a�/��1���>z��ǉ{Ű�n�е� ��xc��P_�`j�%�|��$�u��Yz�nX�H&mk| $1X���P;�d��� �B�����L�t_��%m����(��䰢���ZEy�b��Z_
�Ε�����G���&zd�Nb[�{'!A�"�~r�*�����J�|#ux�K�{���C=�#�É1Ӆ�J�т�}��0N�g�8t���=�����GS��]��@V���)���݆��Q�E�ʲ���_���� �Y�Ӹ��8��<�N|4�th��W�"jx�����=K��������<9�9'���لn˸��V�"���M?H��D}��w���ܻÂ��f��R�4��0@�|�|6e�*{\���L�?���NGOЅ�l��G����b���Bn�)��']pX�����ѭ<f�����%�P���� Eq,SZ�2���TAqQ$Z�`G��$���?���쯉>��e,���f&D�<J�N�v�E8�e-�O
��0��x6I+hWH�� '�4I���^xeE��M�k�M����E|X	�\dOv�CS�Gh7q����?x�-
�u�w��y�t�ҵ�
"	��!����w�o��O����� ��D�y$nW���
w�TC�V�ySX���	;�Bcc���E��ç	~��q��/��7�u�o�M/����78�����e�D %���|�I_�f��6�f(+��NK5���nSsA[����PM{阴�/�|�~���k���E�ͫp@̜�|��H�{�� jo�M�M ��9Y 	fН�N�z �N���hu�D(_�:�CZҙ΍��m��jY������=d���oA%��u���|.�qJT����GV��>��`ş+��i�$�������1v*Qfm��1ݽo�Zu�����g��#����At�����$?]  L�-	g}���_��a
�!�9�`�W�m��Y�̚3���B��l�Gt��̇�VZ����t`�����J����p�9k���ͽ0����`X&o�(b�{�V^U�i�����音�|�����b�����ބK��v������r�O4�c<S��Ĺ��m7��3���l�ܐ���Qt?���5޲=���������4}���NKw�~WWڞ���}������'�,�8��.ѧ��"1���SeFp��qm��I7*���:Ԏ1�[����Ս�x�m�MQ�8��4�M��N-��,��V\�LF��E�տH�L�$��E)������
ɂj���(�u�.����e\P����?�B�����?y6��&����S�?�������Ʉ
����-�-Oo�E������h_�#i��K��g1	�5}�|![�Ww#�"��z,2Cd*{�/^���n�wޱ./% �z���?�I��%Q>�b�޷���q�AˁY4�!���euYǼ.�ܶ�Jg�L�z� ��z��Y�=�i �绹3��J�����9ьN$�`��
���I��<ke�e3�܄��p��u5�^)��P����a��� �~sԃ$F���F[?�/[��jLW��	 �I�Зc�a(�j�j��+�C3E�8�?l3e��/$����x.@T]WH��5�V���mb_z�x���	{6	�!"�d�~^��3��c8���X�����a����S$(E��s�O:xb>"�i��I�Q3yo�C�]�#yy̝��V�����<8�Q;��I�>Wo$�B�@>{�.�B�=-E��>b��=v�A��W�H�5e��PvTk]��N�V]?���>4%�P�O�+�$ݬ��q �<��k*^�=�v6 �����6*e�4��˪�YU�s�_�$�rZ6��n��99rR�n������< ��k?�)zE����:��$3)�蔧C���':��BU��wpS�|<�OQak��KǻuvAۖ>c}���N^���bH��=�U�]���S�kJ���J��E±���	-��6�)�:��������V�'~�;ٗh�0��/���zX�p_�8�z��SRwQ`���9�d���n]3x�番�����:)/t�yu��_
�))��֨M8�(�e3��h.@Fv8`�{�m��Do���M�qf2)�D'��&E�1�9�M��i+�����2i�	td�����p]�j�vj˩Gg�g���"5�&����D���f�#8�R��*���41o���8��뎽w��];���T�`� ��h�O��@J��@�*�*�C4��3�wP$�
$9Ra�͞f�qM�������Yս��;�L^��X�lL��]���i�����J�aקk!�?3�՘�ԝbf�*�⁧���{qN��i���0�Rr�ra��[���5d�Gi��������(� [ITB7�[��e��n�� A8w�!�C�`z���rP_m=ekJ�@�<�	�đ�ɷժ� ������'��&8>�i����[���Wf�Д��W-'��KB����|�s�m8m�O�A�ɟ`8H�chV��f�����Qa*x�r�E�sK���c�Xir��^�����g�F�m��1S��v E��9���w��Mھ�=�teBQ���_4ϰzI�0�!Y�lV�a��c%n���X��>��V`�8�TN=�º
a������sR �BsB�)�-u�:3�R�������M�s>>H(x[ϽX�4̕����{�c}P�%2^�5+]�tG�G�f|�8�"y0�%��aT
l/�X$�8�*�p�JFn<4ʟ�4\�LKm5l���S��O�@�0�v(��#�\��w�'�2a�S�?���J	�S0�i�����&��Էs�Ǆj�7�K�S�[�t�P^�>R���)��,�5���T�3VaK"�9)���^��h/�q�]�P�I�ug_/���x��X��cN��Ek0���G��m�7��V|L4��F��##Vb��sTd(�o�fiv�b9��Mּ	U���:�w��AX����Ԉ\bB�G�CA�c%RIQ<��y�_��ʕ�������i���=F���*�Fw�!����6T�r(�#�1i�l1������ʫ)��^�T������ٽP��!ܒ��W�U:�����P�wf@�3��YIH�]���Yź��
�Ϟ+�I1�q�N�Pu��i�UE�CS��D㕻���U������oa	R�	Zw�V� F˙�y�gk�bֈ	�6��O3�LX#�<{�o�s��5W�w@��f��C2}y��(�z��I~�wL�~�i�t�/�ѵ�6�mg��qI5���ƿ٠3\&��Yr���`g�e��j2>��o��hP��8��l�@�TM퀅������p�E��)g�?I��;芽V����2Xç�*9�Y���7?2 �CU~j�����$��zƛ�1���^����4u�7�.�E�2�ܑz����P*WN�3�NJFP�Ʒ�%���W���OvK9��jI��xE$��?�3fV�ud�\gVi�W"F}���]���&��D�֌��İ�R���&<6�,��������bH��{�0��R-r>��_�e]����TJ�%zǛ�`�����6y�6�5���~�t�;��;I�+({�Tk�{�F����Յ�Z�}��[𽘷�`L9OA�:c����]��5�M�2�٘߅b��﷦ۛ��Qџ\��ܼi�g�'�
�h�)��G�#��o��cUuv�l��n���F0,�^��~ ���"�&'*�4���)�t6�GμE�'*����1�l{���VH�=��v��i�(j���\*�5��5ӎ&����AC����S*�כ���! Gr�X0G�O%��U��>|밴��Ete9��h�q'��s�@^�&�tј3"�A�	��	'yͫ�57��/f�9����0t��w��:�f(1���5�N��(s�D�ڙ��&a��D��kN���|�"�D�I�����!���%�B ��1���N�V.ORz�D0'��1�D�	��p������<\�2�:v��2�� `˔��ԖK&{?���3�q��z��CIg���]2)�]�����#=T�41X�{7$�r���lR6ڬW�p�d?"HG���	ګRV�8��N�6��d��k�eo�j��,�[��I��:`��i����\�cR��!s�V�̺�oIzmߢu�B@ Nl}c�52M$���cS�P�DW�Z2��}
�K�!���fb3��A-���_!�����U�����}�Z�O����Ȏ��U�Q��AHj$�sj��"{�SsJ
�豀��ɬ��q�G��˴�[bg �.�Ҏ#�ة<�f��ǌ�Ȱ�����D�R$%l8+�������w+N�R~�0`�M�� �m�,XJq����w'�?j\ �@:8���ğ��� ��tQ�����աA��WY�
����q�t��ԶAHe���⸬���K�նs6����Uɩ��v)������Ş��;t�۫���c����?R�,4Z'�^X���#2�wT/�o�\�ۮ0������K�t͖c)���A������I߾��h�������p:/��!RF���T�>gDLA�0���C�����0����_��($�H��"���!��N��!�Tul��c�*ŭ0������e<F���K�_� y��:�.-�u#�>�E.��y�.|Y&�.�J��cb�o��^I��g��sK^�I�|���RK�"�ɂK�a���+|��hM����(��W{�/��ZV�9�q��U�#i�MF�H��n�v��L���$���o�j�d��Ҝё�
����ơ�Hiٛ�o����ӯ����+5��{j=;&7uvJB$��U]�[[�S�X������Ӏ���X�K{���h����t�>������w�.h�m�J��A��{Z��Ht1#!�>�}��f-8���?��++!j[�Y��(u�J��l�W��G�F=��1��z3%1��`���R�ٵbG�`�:�Ō�c�������DS:Ad��}�6�G�Ͼ�"o�N��'�%W�+��4�2H[�nU�����Beٚ����G��������Ֆ5��!h4��8]vo�}`����OE���_R��-�����#�Zy2 r�T:����&��.��[��Ze��Nb��Vk�%�ӿvS�+U��,b%GՕ��,�i�.�{#٣R��j��7L+��!�������<�ra��"��y�ؠ� �E�ԠvX���cժn{!�~]�3U�B�mf�;TP9g���(ݰs�5N�����s��M*�W��B���ph}F�/��X<�
��è���D�om����˴v�qϫvk��#�Sl�w9���xls�5݃�'�Tmn"ɠ3�b��^|e�2��2���Tס'z!�*��=��Hq��)qG��G���s�pnT�I���؟0��0�1/�gō�{�!��.�)fW"��}���`��ܗX9�,|�$q�\�~`��rR2ν���Z�k��5���z�̾nj��!p'�'���!��.EQ���3���>#�k�{��Gs�����jtd{s�?�K54�׺qe�+!���ԏ5��8`�ө����'1k0	-��eh�>c�ϭ�_���ڃ��M����J���m��M�W?��Ap��d0�#�i����Ł��u�Y�P��w&]�L\b��RT�ſ�g:t��T�U�?��}�BQ`��uF$8\7UH�>���]N���S��"m�v��K9|�������$6�t�a�d`$%>k���I�s��t�Jl���
u
��<���z!7��-��"�oY�Z���������u*K�v�ڿ?6/����nu�ᗂ��Y�N� �{1�U=h�4\;\�F���fl���WR�ה>�P�S��(�[�K֍rZ��7g�0��ԹPO�q�~H)�����x�q�c�Ta 3�졽JUchտ� <�w����g�6&�	'.�c-jY�q[��a�O����?��1�׵1��"U~������.`�*�]y���r@��A8��rfS{Q��c
�d3��B$����[Ռ�����۪�1- Ƴ�>�uJ���|j��0���B�0�`��D`X7���<{<Ԛm^��x/T�j�/n"��h���������7�*���^��Y�dQ	2�=�u���mNFӼhAl�GE�$O� ɚ���*��6t�(�(�{4B_⹒�#�����./%����3kd|���#�]M�O����򹿂R�<�Oը�S����O��;�����a�"%�(Jz�t����h=L�F�v������������Á�O�>C��H�m�xZ´�o\8;,7T�����_࿓D��=��ك5��7�����H�_��s8���U����Op=�6g��\Z7OCW��g��j��r�j¹5�Uc�\0�"ڝQ-���ep8)���r1�(�>�x�9D:�9(ܸ�0�H���f66bW�g�!�¥M��gq�ˡq� ,����@�-7�lx�R�Knw��I=��nI��y�v�H�����RAtz�er��I۞�܊z�IIq%�[[+�+  � �����F֓I��eA;�)dA�6S��P������H	��sQ��FFZn}-r�������m�E�b�Vk�?U�ģg�y��D�:E�(.��ߊ�q�*�L�H��~�u�37���s�22�C���B��*�qn������]�w������1iA�
H�p��d*��|�������R<�=�s��Q�)�]��� ����aȪ��R4��x���{gt7U>�`}04vcE����oE��@��3T��#	{����Q�2�U�/v�Y�iQ͠U�nvXr��6���j�����8�>���3�	��h$ڷ[�%}��4��X�Ȳh���;F��rP�~ƞ�a�*ֵH��ׂ��ͥ�z��(���Wy��[G�}����B>�|#�X<��I��n��pw�.�>�^rN(�k��z���)����9U0QTg*W2s6�t�4�����$�4�%�؛i����(��0wH�����q�&,-�-�7)�GJ� ��Lp�]����r���($�i���5�Cd]��;pX/^]�J{}p�s����p�=����T>q�����0��x��5Q�̝(<ۤeR����&aI�%D�k����V�ǁI_�-�+$��y����߹D1p��JR��{,�\<
�<]�48�LR[Pqu�c@yx��3�KwH�8�\��_��6|�ױm��ݎ>�P�B��1����Y�ij�`��Z>�34,ϋ�}lP @]����lזEg�Q�F����p[0�״F���\}��j$�eu��v�=����5]%��9Ϲ��ZҸ��8E���@iU��Ց�Q���]��@s5*^-�H:t�;�~%���0���N�=s^|�b��"� $Ͽtg�[���ɺf���{���v�$��Ѷ�׊ߌ��`XK�u!Jt:�N�9*��wvE��W5�]R�_�����:�~�%�'�)���A��S�-��f� V��w�s��]\KB'T#��1[�=3;z��7xi(P� �2�/J�\m�/_�����C��jH�+�7��$B W�ab�d�<�8|{�vj�;9a.�_�K�dB�Y��! ��,�$<D�[�he�p�����ӟ����3�@����k=�@��(�a?#I�g���9Z&����L׷��q��$� wY�b6ve�c醙q��_0�>�B�S�<Bx����L�y������h�--�p>:m��a�,l�1���lz��9��^��Ɠ�i o1>����6n&�()��g�S�-9�N�2�i�j$Y/_���L�y�^����G	0��B����\^��w���,C��zk_K+��+�y��P�'M�1kwI��	_Ȅ]��sY��k]n���g���W�%O�(���M<"?�V ���AA�U��/fCL�^{����� �j�|i,�K�u��͑0����}q�E�Z�L�g�T�@��t1 ����֤��T�u_#��t�t��<�6�A]��PӲ�����T�-��T������pi�:,5�x�V7�<��n��?�^_LC��ίh;�}��M��;�K��*���?���+�0�@Ǿ��������_<��0�5���լ!Q}�'�ͳ/��{���p�ءsv���u����䧹��B����Ԏ�s1�h\��%&t����ZEXMO�g��3�V֜�M'������XCjF�*�W��!r߸��m�lNT5Ba�PG.Yj)'|p�����)A����I`e ko� {\�qڠ�(d"U���&
�� 
����	�!S-dKc�� ���{�|$�tv�ҕ2e�� |rS���m��YvG�`t�"?NA_p+XD�hH4Z�n���c�u��n�c�O�s[��0�x���b���^��6k�*
�D���*s0������25���ܡaڻ��+�87��+�ko��݆�V75uT��
V17R��MEV~Pe��Rj�N�\��]�+$(7���р٩�br�;3�Rξ7cH:<d�k(��H�_��+ٖD��L�s�M��Ycd��=�.���	�D$n�܀ ~w���Ʀ�H��
:]O��jp{��	��G�?�?(���6�6�ǈgw�l	IZ�K��uΨR�1b�/�ۚr�U�����
��b�֨g}�]~` x\�O�A5=�)�� n�ܯsw��I&1��`w���S� 8d�V�(�
���ت���!��陊e���<�|�Bj�0�bXo�oGlV��Ԛ��p��wz�Ȁ<ߘ�!k�"�\!E�hq�M�4IY����gy������qlaB����g���q-�Xv1#�?�Lk��0�E��p7�.[����x�����N�~�N�p�i
�\E��%�/�"�,�Vä�T��������d�c��%yB���r�P��''��_�G,��[�Vkm�k��p�t�3fM��{r�|.�b���0����R��������Tew2�*H��\���E����NE*j�������z��w���/�{��*���w�* >x/W�c�	�l�{��o����|�I#�z[��o�Ҡ���ۦ���چݗ.u]��f�/�nٓ�~��T&bߕ
"ܿ�����; ����nEe6�<���D�j��ˣ1���h��N�;�A0�R`X��YHl֭�5ה�݋�2s�'�������Ta_~�Z������Z\���)lL�Kp(Lţkh�g�� �TL�Ft[u߳�����5����ڋ] �8��(Z���_baK ��[��!e�W�uv����O�p�6��>UGf�q���.M�����=u��p��B��1ޏ�f�v+e�3�|]�e�����/��PBl�W�^�	����	<�Z�(b\��4��~߭/�4���D�����������]M�������;��&�Uх��1���wsy��K��L�i��I�ۧ���778��R�B/���P���{��	�b�0r�h�}Wmv��
r)H_ǻM�)�ӥN��{�7���N���'ի(��󈔾�gEq�����s
#��zvy7*�^�e�(G�qg6�q��qo ��?r0��a\�6�����	�6�b"=jĉm���R̿8��<��^" dEu��i"��>-A��S���O i�a~�\�=����)�c�(�P:#�m�6t�{���������'^���yB2�"GC����q��N���B6�b����*���Զ�X��*�S&��A�*��x����quj���H��'2HYSdù���mA��P��4N��Ep��cO�V��*��
�͊�Ƨ>�d�Tܴćٳ/����?+���/R�D�a��H=���������RJK��p ݻ��ȧC��r�39W���J8��*x,��c�╬��$�GL�V/�`GY���G������x���|
���߰+�b9����B)��c�
�{�9#�S*�FO)}�Q��P���h�Qs���CT�ݖ���Z�0�ez.ѓp/��#��w���*֣�C�j�UD\xRb5_��r�������k�A'rH������i�Z1j�~%�xP��آ�"t�R��E��4�M(@Gst���We�*�٪���7��Q�u�OQʳ�2+�"����2�fE�qy�U	?+�ˮw� q8Q"K�C�y9�Ĳ���zu:�Z��t�A�NJ�+Ԏ���:d�k����Q���1�#8�XY:���p�@�U���Z����ؼ�[�M��)d���Ps�`P�"{�xl�!�ڔa�����=� ���d~��X2�O�KC,������Ȃ�Y�k�j�0�~����U�(\����(f±�h�����/�C�*��y!��B
kO ��n��d�\�H�I1�,6���K_*�a�w�-ƭ�G�\͡��W$dd��ci��Vb9%Dˢk����15�/k)F����Q8��tG�
�c[��c�'� 35��+��Μ�A���p���B���-1^�X����J��M��^�t���w'4;�5��������.(�2
�m�A^���^����S�Qt�!";�]	�?&-�z�����7�V�N8����="�(��p�m�L��Q�:�QGvS�QQ=�i�V|��!�d��%d���8�O�F5v8`�e�AN4�����#F
1���| ᘂ�fQ�ߍS���T^�@K��
�,w��-��8�i!V�>_�\��ԏ�e]62�&���9�C-�Vey�Ӽ�L����:�	G=?�?2������&����M��h�go�0��a���0�@D���x"?�v��;ߢ�Zq^�<��]�$N���8�2b��q�aTkG���		�@���|�:���G���U�����\�:���s7bwAx�Ձ��
%��ѱ�wo����A�S*w#�V����[�h��|9��ߺ�=�G�%����o�<"d%�z��ЩQ���VY/���:�v�T�,FcH�[�l(�k�@����7����?/���q�u1VX��&`����HC`Z����a���*G�1�MKﴞV�-�J�����˹���hm"�ҙ��$o�<c0�=Q�W�3���Fi��,08� �zz=Euu���\7nlc����41��yؼ�Eǔ�xk��Ns\��������7�$��P�E<t�LZ>Lkd�a�~��j,΍#�2����TՕ�9'�L"t����0�3 ��;\��?n�=ƌ�W�Y��F��̪U�]qSP���z�m���2Gm���;�/�=���&���1� E�=g�Yˆ�!��Jt��N�A�F�jꃪ�������g�Ԡ w��ڻ���QT�t����<��/�Vx�M�k�d���ΰ�1A�ЃR�Q����q�/�ҹ��,��-|_�7K�����V7�m[���v�РP�'�s��`]�����©*��n�N��A�n2��X�K*	����n��9I����2�L+����d�G5�>�;X+[s*"���Kiwd:��t����hIܸ��S%��+H���S�[L�ٻ�nS=L��<"���r����X�/( �(^�,ԻS��T-&���rj 	hr��ԫ�+os�<�G����W��?My��h��Ȍ ��m�ō�v�b؆-�Ο�D��ah��`2���w����7�;p��"S�/�&BI�3��WZ�d�ƃ�a���X�ڟ�^�2ء,�q��=�KHBT�n�$�Ұ�\Zw+�wHr�I��"?Y]��i������}ڕ0���!����D�"-v�Y��?z�_1���#�4�L���u��T�O�E>?�uF��W������#�P�Z��BZ���)$T�3$�@K��n�*7@��w��c���Ʋ=��s��V�x|D�}*���q�#�����9u��i=���+�1v���f�滘��2ܥ��/9b;2q�0�0zN4�g�{*��BWY�n-c(�>��  ���^)�~��ӻ?�f}������wɍ�	yM%��L���l�M���Rg��q��mm@z���ؔ�QQq��r�V(�n�P'�A�xldCu޿3%��ш�d (����[;��������D�kB	�by�̎.�2Gq�2L@�R'���u��4V-��6f🀇��N-}x�5U�߼ �x^G6�c�챴h�F(4ۉ�����=߫N��3��r�HWG���R@ck.���>�ۂ�.#��@\�n�4%�2?Z�A���'�5��ےx�b#��Fk�O���BX���~X�!qX_*���?�V�'Ȁ� �Cr+�G^ٳ�`�Sd�x�}Q0x�i+���7�\;6��N�.t���:R1%.������m�~	4��%B��W���V�U����~��H�iBLBm�VE���vx��>8O3�T�'�X��k,��Q4m߶���у@+��{�ق���mUGU{��������eq�բ�.MT�i2\\��W���&��d;�,`;��Ќ����f�R��c�.���X��F�G8�o�g~Y#deR
!w�������H�?�Z�e�I!(�_��#n{�%ԂH{={"!pw��:�j�\]nA?�]RoV�hl�m^Ҫ����@/�� x�w7
��8k� b`b;�Q�:�e6�0QOP���+���0�[CL'W������x�-jT2�X���$�<"dΝY�!���O�%KD�Q�`MC���;���+A%�	pRE;L�������D!��E�'$�G�n��V�R�����|�92"8����+�<V���^t�Ğ���W��٨�;X�=9g4H 7��c���	N�B�����)]��
('��~Ed��l�p�)5��%���1��8z��rD&b���1�eл��Nq-��A6�:֝ww���֬gs/U�Q
t�Ӭ�����	A���l؟��|ߋ����`���e۵��Xg����t��Pg�h?l�dF��WFsI��Vf�,Nd_S->���>L�þ@^��@4a/ւ�G&$)�9b� ~edw`D5|�8��`����kM������t�#��8�}��s���9��oL��kz�m��kfl�4z)ã}i�Z��+-�l���9 ��F�Tsz�' �\�.�c�l��-Ėfrz-mV(�҃/�ά٫^�?/�;_D�Z�m̀�|{V�kL�Xa	ʋ XJ�*�@�4� P0�B�z�S�K}@}�������η)�{e6j�We��M�گ"m�1=�`��DU;E��������Tn��ۄ����e��)	d�4蓢�2NV�1p׆#h�)
��?�𢁫O�[�k'EV��g'�D-����#��k6-t�
��~6��5�k�΋�ޤɴD]�����G�SF�w�PG�ہ�?u ���?�d��X9"�:t�ۅJ��Q������oKfA�5<��O�+�%���5�y�t����E�B��Ix@0���ݑ_2rVF�ߺ�n3��}��2{�5�N^�J�4eH�@.���4s�%���Z��x@:���A�I��r�P�����,ZT�i�?=m�45DI'�8� s�]�����m��m��@J�x+8�.�tG�E-�ݩhE=q���$����d�7r퉹����b1�'m�*<�����s{��l(��L6I�F@#XK��XJ�+5��f��+잼2]d
ˢ�J���u���/��� �&�'��1���E\t���x���w�S��z�����. �=�f�<��t�e�>�����IB�t.8��IF�N��^ݝ+լ�u/������44�6���4�š��C���R��i+�KP��p�{j.QA�A���)vљ��eXJI��L��n7��@��=��a�8�3�9�;{*rC�-�.E �~z9��?ǿ�W�n(T��<�X7�b�F��������������(�[BNU+ęЧ�R��,�0��ѕ����V�:���!�;8��Q#G�6�7!u2y�h��ڲkQ�y����K|(�b>0��8���F|"0�ui[��#wJsW���i���"2��=ed�n%�r�Xlw�O�xô�5�SKCd�J�9Pą��|u۪�\���\���@����x׽�܉}�F�C�x����P��R9c�m���ʌ�^Rͅڵ�HZ����]����(B��ܽ��VS;m�������I&��|�z�{�^[I�� <B(�5�F̺��&��o�����S���S0�x����ʃb���	�@��Q˭��bԸI{4s� j�l �!��di��� �&�pgV%�����N� �>����R��L�U�p��uW���m�(���~j�,��MoVO��^X��"\l��.�"����ʜD�%��K�׵[m��D�c��l��3���w�p�Ut���Ζ8,J=������!g?����o����@���K���K�K:����C��>���%����(>�R�J���;����`��%��XW�������Қ���ơPb>:��s��e�_��3\9�9���Ɔ'��'yG-E9b�#Hâ�+��I��N�q�H&���˸$LK�D�ہ`�+�둁H�Yc���f��dg��y�SH�C��XF�J�'��d�����8���x��g.�r�����%ipY�8U-9���u�._��D8�qFK�
�f/�=�p���.����{�`>Ss��D7?&o����J9�QI�|�C�j��%爦��y���L�J�"
��MW�NQ1�� q�ƥ��fhn�rx��<4�\(>C�7T�ݜ�
��z�q��d+Ȅ�cʁ�3����z��ӨX*��n)�"I<*���!qC:�5g��OJ�=A&I5{M����\Y�Ij����F{��:R���޼1=�×�/�[dMu8��&��F�_:�O��!�X��'����fBO9��:!���fv��Y)5
�`�1|���ȋ�	�5��0X��C���r����obD0?�)-c87���fu^x���E�`��߭��,ѻ�A��>���˨������ ��$�ࢤx��L��jc��
p[d�C��
�Ɖ1�d�*ww]Bb�1$�vaoh�s0�e������#bL�k���?�-�:^�7h7ǘ��bW~Rm%�jҍ{Q�} ��u�(-zʯ��a�m���(�ZD$Z�F��+N_���pό��Qi�s�x��R�A�=gK/�E��V5FE��c��ݝ X+�/��i}���c�J^��Q%8�F���
�Hǥ��D���:�?M`z���݁��@f�.��5>�IN)'�Z�0�F5_s��O�k<G�h$|Y��oR[j*�Bo������0��Z����5��;!"�h�f{.��xHH��\#� �A�F���f�%�O���p`WxGDq��p�D΀(s�u�A��sTEf1��X ��%�)uq�:�������,��P��^��F���Y�yx�㊕ųܮ�tRe���®��0�S\���k���z�6Pq�E/\襙�^����ȯ��|3!��h4�V����t�]������*��$]۩:�Or�'-Y<�F�8�C��#5C�m�hҌ0A����?m�N����onކ��O��t��-����ǝ��͠�������:9�N����}���R��#��mKN���H�~I�{�{�_�'i4fwrf,//�@-^�1��7���z{�X(�1(������������մ\�6��n ˧�iO|{���H�@�ƮԮ�CjD��@=ſ	����{m/�m�jL��,hZzءx,�Bp	�',����ϱX+]\)�|44��+ê7�|�0�V���r#���6F�,6e�s�������5�.@��?�Dvsp]�hV1��%'�V�d�I�c]B������/�y����Z�jͣ�� �# Xj9����a��q�E��ŗ'�k9.E*9�`o\��ܮ�,���#�2,����lϊ�w���#��f��f��1 G����V��Fd,rYo��Nh��T�)]"rp�	�_0�wG�Z�`Vͺ�i�"1	ߪ���ir�q�i5�\�u`������+T��>Ay,ph-R�\~���>�I������}]w�犋o�z��RF���\ƿ����V�=%h;�Gi��?���~�T���T��+��Wj�:�;ޤ�z�޶�4Ķ�P�!h�T6V�c�xO�@.�C���v����L3����k��r���O�l��D�&2��x�6QɃ?�������O��	]��e��a��Ԧ]��b7*yl�+�KoD���4�0�Y"�,n�8`�.�ǯkK`90lQR�І�����7X�'^��U���&e��Mh�x��3���'�|}b������O�lR�e�c�5�&u�����S��R�6�n�� ��*4>��9ϣ�����6�Y�]�5��7�O	!�V}8Ujur��M��M2<
���6\��~l���`�87��WW,�1M���Z��FKS�	L���!S��[U��"�uZ���I��.�4=�}�g�T�.@��0�T�hms�H��Z=)�1D*����Ļ鹥
uq�Vf��E���{�2uq���ŝ�5?���b�s�
�b��;E3:߰���@F87�W�� �����K�O��@�JTЎ֌(�6�J&x�����7J�ء>�x���-B'aQ�����8�r�g��ks�T�W���1��C��BD(v�a֐=2^��R9�B� ��dۃzW|���?$u��3P��C��[ҧi��Wz$�E]뒇�� E	7�Y`����^���tUyӊ���8�R?1�\9�P;p��k�"���xwo=]V��z�LtN)��j�^4� �ӊ8��)(�Qa����
9��3���U@���������� @��jpo�fp��7�/��?�Pg�t����?bq�2I3�t�T%lF	,�D�)�3I����������X:{�tN[*�ʑ.�>H;��K�
sV9V�1���oNan�
��Pۥ/#Q"��&�iQ�l�R$ur��u���ܛ����I{��S�~� ��'����g� UT�K�X�/s/�,�2F�J���78`8��P0e��������������'h���6��\K~��ɞQ{�������u���¶�%���M�N�M��'��$�ǿ���*����,��}C�To^��j����w���o	Eb����+a#J	F�m�*"QlnJ��ե��`�t�n�O�
�QG��d=�%Gm܌Y�x;�*U�/ߥ��vD�,���
�{%Ë���$��s���kv|�!�F�_yp�˳��`�[�ݝЬ�����$'z���TZ&H��O�|O�X���t�
�<�������+5Eiѩ�QOB+�ׂI��!�3��esߠ��;���WQ�y�D��]�U>���`<(�>� �@qNC2��I�,n,>)�U�uoT7�%��H�պ�U���*�oE�~g�q=��~04���'���l_^�?�[�WP�օ#^��wz1I�s��dO�� ���#��]Y E}x�/Ki��1j�[����ϱ��������:QMҊS��%�X��b�G-Z*y�C5�+Q��7yi�(�e�.,���{Y2�#� R�	�W~����CBV5j�!���z>���a±GV=0*�o�6^u"���� ��?6��s#�P�hE���eld��h�o�M����uNކ��IGp��;�|'C�̉����4��)o,	�\�M�;�mer���8�);>{u}��-+��`NV0K) 	���NX�fC�zr�,�"e��Y��'0�_��y����k1eI<6�zy��͋1�Ĩ�ܘ�L��j^�ϗ�EŔzI����'s�������@�7�4PkD1�������I�b�$?�74��F��l��e����͗�1�It {�=�g���bn��=��g�M �N�B�6�y�܆�+����.�����8���_qz�3$8�{�E5G������S�.����Ґ�[X�����\�����3K&��� ֣F7�8���P+�� j3�o-�WH�&�n�=���Qw`�F��PJ'W��/�~�6����鿟�zR�~sr���W��7�}6h��:Ie��Ƕ�p���-�Lj0#c{�^{P__��49��jϝ����,#��V)D }'ܲ�pg�e{,� 2Â]�([�`�~�b�Ջ�s5�����1�P6sr�_���=�v��F�xm�uX������%��HP���*91����]������	�=j���z��O�'I�5�A�] �^fGO��\٣��9E�+�h(�������҆国}��$e�J�is�&v����"ǳ8.^ec#I��67�Q� �^)��|F]���br�-I����.Y{i h�Yâ8��l&bZAt�Z�����*G�<����(�|v}v�H�3I�$j�c����N��f�����X���	�ܿ���a5������$�R֊܇-�\�)��ш�5_���qe��yR�[����+�!\��0��:��{�0^Ö�]A���6ו P0.�m�<��{^�/TV؇,-� �92��UP��0��D`օ����Q�HH�-2r��:�M*�E�/o��\�->�~{�n�)�Z+�=��l 0g�����?)�����:^S�Y\b�05�u8���̍������a��wc�-��;���W��O�=�he�Y����N�9�YCo�(��#�H�m�1$�W��B�s-�2D-�'�H��V�<�2�C���G�Jɱ��ݫ�S��Q&����PV�R�p s����L�����v^1�����"I�r�?))@�rc������'3~�qt�u�-�;����1mt�h�/-jN����xb�)FP�D앦e�M�1���=FT�$ ��m��Me������Hx�Sz$D/C���e�LTP�&^��E`�oQ:O��q������S(į�����e�w�����N�?�4��&���q����C�!��%�V^�mPwS����M������:��n)��W�W�Nm�^�#1jd?E�.`�i�3(N��K��:P	j��M��u0��o �C�U7A���:��4����o+��=�@�z) ï��b-��f��-#�����F���Vi���L:l�To�kZE<3M\b	�F4c�p�:��G�-��"�u5$�p��j�_|�[{��/k��0�PP$_8�-/�L���^��7�]L_TI������ޔ4��1N�nna8Ȥ	��e��L�<H�K�ؿ
����(�I�4�Tn��n~��v��������(�EM�,w�4�V�2n�r!�t�@��7}��	�|���
m�v�ǲ�k'��k#"׀��y*ݵ[��<T�][@��H/�H�Q&)�����+3�_�ƻ���k��,�`H�*o��Q��bj����� a��r�D'�D�I��L�L�l�U��O{����Ua�$`rY�˚"٪���1::w_���. ��ݵD=-�4_IpPH��;��;�i������m�ra�
�*�v���dI�rw\m"L#�3�v2���ʄs����1�Oo�\)�u���|�Emn�^��
�0�ט���up�N͆��`-��q�+g�����%)5�6�g�T��\����c1��	T�5�̉���"��hmP0�T����H���T�����`�J�n��t,���Nޜ�yhp�NU��%Z>$�9ќ6�]��3-�
 ��X�	�,xb\=�?�>�R�D��D�g0�(	\0�4��_J����VcK^���;���g�G����Ez�Ow;�˞�(���ڌ?&�J�M�@��Zv�ហ��5y0 -4I�j:V�"�Xו5]o�ZC�S���gi�bÅ�Y�˧�LeC�� �����ٵd�SW*$�T��@�ϷO�ٜ?��fJgѩ�! 0)9Bw,$��}`����d�1A�	�p�1�L���nv37��T�#a�s�!6V�U7!��oW1����8rbZ�rZ�
���=��5[O�����s�pI�=A�붼�,^�N��[�}���������� �__�8�Y`#���v��0MԌ��-�9��%��گ2�p�:;Si}�?NM��L��	S��;|p���BM0%�*Q[O�uӀ���#��j�5�|Sxy�\&?E#����1�&����"L(�/�� C^A���Z�v��Mü���1{l]�Ȓ�ZN?��4��.H\�K����D�
��\`��ӭ�`�O4��\YZ����U��J������b4i~I��|��sѯ���ɇi�w�p���+t��_�����M+E�O�;E�����"})�#��8K��]�@~�P:�L_���^]�c쓔ܛJ��Rx �5I�Y���
��������h��|�X�B����Vo�W����� �tݣ�>]��O7>g�Z����̩��|�/(tV�j�l�\��y.�W�-8���ř�>W�2�<W�?���[A�ގ��DN~�i4",t��V�����TL=Nx�/kjC��r��_�{�#�!V/�@�P�p��D�=��Ԇt�VO��֟����ăK�4W�9�'�Op�������Q�F�rL��wa��(ҳ���pE2��R�X¤�"���vq��X����-���a/�:F��Pb���v��b뻇�H��"�e�k�u�B�Y��C�R ���'D�|{Ċ��4�埥a�Ha��+�
�;ǤC�L�sr�)gC()�td���j�n��� �skY����]vȐ�1Q�Pa6��q�[��!U�e��9M�������R~���3�I	,�<Sy��F٪?}Y(����E3�	M֌���m�wTWL��~t���R2 6�IDr��֟�U�~nk�A�Ӊ�g.u�@����LO�ڣTT��V�zY7��5���l����Z�P]�eF�^��YC�ݔ�of�hX��_�qJ���騽�Y���9�#���m��D�U
V0	��x�ʱmF@��S.n�o{�	�Xo}�+ �E��5|�il��R��"@Ͱ�~G�ױ��N�k"����$L�b+u;e֕mI<4�4�(����#�g|I�I�RBA,��)���ٺ��9�$�.�S��XMz�/��P�D�f׊:2�Rx��k�5#��יT-��T7/�\Z��� #�,��b^#��-�K�ރ#�]Fv�g���.f�Cf�������&(��D���U��of�y7��>S'Z9Q^�{q�0���m���>\��S|8�f�[/@o��z�l'ub�[ȣ0��Y���TG��(�F����^��e�clwfSj����N�ENX}�.e)T,b�X��F\u_p�<�g����aS)����p8n���S.���͹MRvD@�eu�w�!��7o�~-�@�����Ǜ�0P�?.�w���5(W<�lkEB��[l�<������Cر/��c*�+��23��7����*�ȵK���a�׎��E2�Mu^P�T\��<�>��Hw~��q�ϯ�sm�����淉S��Q��A4 a�^U@G�9��!>0q}�·�UP-ӏ�]���n+�����;�D�%i(����#���ɍ�Ҳ���Q®}�����xI��ǋ���{��|�8�m�_�++�J�b���v���"��Ip�Ϲ8�.��ʽ!�s���ՇkKrec�4�`(}�~��
��q�e�a��b~}[�oؤr%��^�4Ǉ��A���@�J���.��=.�vX���g�m�h��_�A�׎���VyW��Ⓑ�lNe��6�ە�`�C����<�NR�j��OҎGxW+3l���R��n�.�|z9�t�i�(�L�Qզ�Ы�惤���3�{?Ρ1�C�`�Cd���f�V|�
V����FYfG�=����f�l��{;�Ŕ~���<,4"a�S%�.'�-�eƶ�@����x��qѺ 5;���	�'	e��u�s%�)�[�y�b;A��, � �q�� �h%����@����}D0*!>i7&H�9ߑ*M8�+���W 2GI��v� 'j�i��)�K�
������jݔ��^�-�"[UЖ"C�9x�l�?m>�W"bs� W^�˟���5/��Ҡ,[%�(f@êW!�?�*D��5x��%�:uC!�l�Ǚs�N�,��=�@jٽ�+�X+ϖ�{�Z��q��Q�[�|c�4Y��=��'>��
�wZ�U�_�3*���[�f�!^��V�H���xh��L��Ԥ�.�K�Z�>Ǜ:���Rzdg�Jjq��z2]C}eb؅���瑲�U�ޭ;�
��$K��~�C�<+�k%G,��i�&�� %�1&��P��XEQS����L�ܑ��~���nɇ�%�^7׀�4ۻ�Q��Bɔ���B�4���C����������'�8n��i���f!�/pJs�2Pjk������!��>��A�6��
���p��?(قժ@u$i&D-��������}�9ql�WQ�N�+/_�u���}� rz�8!RL�ÄN7(��*��Q�/���d?�R�G#�3,B!7�ȯ��%>���!��h�ֱ��v���.��3�����%m�E~қ;�B� �z�R�#�=TM��� aĐ��f�F
y�}A d#�N-U��X)u�J��N�*y����
���It�;���-_�ƹ�l��ZuΓ��(���0�Gxt��Ot$z�!b�
:0#곳g:{lZ���!S�t��]�;߲6� тaL6V�Ap@z�R�5��	��L}�76X�hg\�x̲�����1�49ro>�|�E!��br��[������o�����^?�ߟP]>�j\ I��tW9��
�u2���24ѕ
<�tEH��79���N�z����cMMU����Mb,��~�����u*ՕMJ��ڄj0
����k��t����:�,J;0�XU��)���Thn�,1V�j%����+~|����E&�d��b�#Ze�e��'�0#�\I˓`�)�aܤ�n�����j:�u|���������؏���R�8���N�(}��X{Q����;���9 �J�I�rtq�~�h٥�`t�QE��:u<.�U������1��&9��G�'�D�zK,�Z�Ms�(Q9{+�0��g6�6n�\�c��F�FS������e��r�|`����ܩ��<�P����<�ְ3�E��YFvה��74u�����fM��[�|�k�f��/e����q/�t���u6
i;�*�������yî�]���l�����Kz������֑������ӄ�i���BX�ʳ��� [�(F���D-ՑMF��@���*/P
ԩjT��6�z,} :t�P�:s)��3_��b�'ʍ�`�GfZٓ�����Ras���ʵ"�*b���e�B~Vm4sk����F �1�nr�O�J�͈�������P�jiV�prR!�ل�9.������n	'�C���w���3��Sy4`�^]p��Z��Q��(ߔv�TL��P��W��ކ���f
s^w{c�6��Nz��(�)�Σ�����g ���|�^dxn'�Ϻ,�~�e,-_�аm����1������Ŧ��Ŕ�7�Ɍ)�� �U`g�m�S��V�����;Y�h�X�NN���O0����t�������1�;\��A�(|�ܷ�S:z面wXH�{��}�勓o+������W��Ω�d���j��P���8 �����|��,�Rv��:Ҥ���<v��<@����߯I,0�!Z��s�dM�9t�٤p�t�qv|�v����	�x��3v����} ;��R�ޣ��2��Vl����J�j:�׷��{�7���$#��͕+�0��ۏ�S�S�_è���U��70��9\��Z�o���Z���P��W���J��n��rAEy�&>��&Т|Sc�����c�W�2��C�q;$�u�B��s��Q����dֹ�@���v/��BR�1��C�]��V���� p~~*�#��-(~'��pB	X�2ד�cւ���-�n��t��
�a	���8,6(Z�U��\�-�/1A)ɤd��7���0S��P[���[vl�T��L�����^F;r�Rى�r!�$�ݴ`�dAؓ�Q5�u\����y�ګ
٘"�v��$���A�%4��N"��b'=f���u�� �oa�C;���<�	����!����t�|�,�jBַ�Ǭ�j�� �ʣ�aa"�z�C�۵U�^ڂ��cg�ٍ��i{����NY%�}��<�/�f� �G�N4�������"�_����N�㮳�M��Th��(���C�`E������ډ��ld���n�yy��K	�D��צ9��8xC$^�B�o�F
���U�����;k��)W0sQ�ʝh�]9j��VI�A�a?�������=��V�T�a��=����5P˷��op��F���Xu�%Y��*����H�:�f��Y��zH�7D���3g#$\��b��g���c�%����*D���U	���o����4KzBpa���:~Z8>%=�D�+�]���F�t��
��F*�f�*����Ԯ�rSR^I�{C/S=^P<��GQ)��Z��Ft�'�*�'��)��N�ᆚ��S֩�s�o�G��IQ���
Q�1���I���;��������Ь!g�9�-�R%w��u����x[	�6�{=}��>� 1@�â��g_�0\��Id�D=�~�A�*^��!� W3G��fI�]���m,c�ϱ0��˳���5R%�" B�v����W��֌��Kɵ-�KI��8��d87���Pv�Nu�ud�P@�X�RWT�bn�\ԥ�7t:놔��[Ym�$��F�X�*�-Gl�y��έBc�s��Sר��a2[��@�C�����s����h�p\\[%/d�ez�V��-�YA�e���{���#d$�S���I�*�U���賗Zh���lϣ�>ȼ,a�1�C��{�
�V,��'q??c�ū��	��$6L�V��R��;OE�����a9��\��;��OW�$8~T*��<��P�/,s�B�̮ �}���0�#x�U{�(�X��#lC�A�7��1��;��+[������� �Ww� �z���I���0�t���Z}���Ɠܺj���A��B��]D�ͯ�c[�|d���?���7R�!9�_��|��F��MV�Ǹ���F~cH^��G��]F��@���g��2�������\����dnֆ����v�"��v���0�L��
[Q�j��k�4md\ ����S4�d2�A�a�FB��k��'�}c��R��e� �ނ�{���<�����\j�L��H���
����6�6�a@��j`g̢�Xn��W�_�,�y�U$�am��MI����@�2�ņ��١���L�Ti�L�;�+����h��q�g>����݉��&di@����B� �#5����^;��A�(r���	�I��F��](�e3����Q���P���D9L�d��x͗�
W\.������I��d����
]	Zc#�֪QC����oڅ/��C^�������^hݧ�A?U��Z-�bl��B'k�"n���}Q���P��"�w,�,��r���苁��g������{�X�~3��~C�B���<�i�os^����Iiһ��;8S�oN����=m���[<�ќ˘��Ge�&%�<�Bcvz��~��BõI�ʯ*���J$�l;�C���~f��̵UA��yw	�q��Ҷ��!��O�m܏]������?�`tⳭ���zCqa~����#��4�h�U���G	�st\V`	v~��X�S�l��9-� �_�:��N[�#�(@`}�NH�-s8n'�K(t�m{�y\�9^�_F[�Ӛ޷gKkG=�ҌPl��n���'��T��\R5'��>�;��R�z��A��M�����S&;�95n8L6��A��c���~�XX��z/���[V��T�ߣ���kz���v�v��%�ſ�` H�b���W�8BE5<Y��Ϋ��w��B)�}|w��E�����E�,��:9	K���OxUGaC� ��6�.��;e��a����@�lt(�#z{�;���Ok|v"��l�g'@'��.G'��l��o�!�I�h�YŅ�牑>�I������M@��-^����0vaL�u׽3�,��gR�V��UA�;�8��H�8��M���G�r"(9��xI)#Vs�xو��A%�/Y�<I�r�{f���,�@D�e������`-�Y���>��D�´�:�0�iw:���1��ݙ�7�p�<�t��d���v���*<S��q�v{���Cl!�Y��WR�wD�=rGҷ�~�z�����ɀ�c�1fh%y�b�W<��&�g�6Q�� jȬ1hQ��u�����u$p%�/��X�c2�!|��/�U.�,�_j�e�I��v���Qc� �F��!������²��ܲݢ�|�]�4{D��>^>�א"KNd����D.�BX����Sum��j^��'���b2�(7$;����l|��Ȍ�%1�p� ��yl�Hs �âGﲘ���.�8�-����Y���"�l�u�,� ���]�A��Ӈ�,+�ڡ�Ly��[�nE:N����<0��<���ܱ������`��&/������i���g;����]A�'�n"C� �����ӻݩ)H�uB.#/�4��#ӆ͸	�����"�Fb~�\}��I��7i̍T(����e�
q~�n|�~�������/�d�"���r�N/���j7ܻ�
ƈi�^qh�?i��)5`�dɝ��>�xj��s�# �O�c�cW���u��b����[��}�66�}7@K�ha�<C1���A�,����3�7N�(��`s{e�d���E5n3E[[���	S�9 #*5���\��4,�YL9%���Vk���q��ǩ��N�����=BK&�`�XI뾡���P�&���I-Ž���L#��vem�N�{��t
-4\W��ݕ��k��
|�i˝d��ٗj�����rch���bg�׀�`UҌ�YR�%oX��6��"һNq��̸�P�C��z ��Ϩ�rcG�o�=٦�S�����힬�X%h�2�-4ݭ~�Ս���~|�؏�p]r�PR�b����(�:@��/≀40K`R��-�F������m��ΌĶ���c���6��L��ɩ����F�`�X/����ga-�g1�C_>����ꨬ1h��E�.�5�_�1�*�=�[�MA��Hw2]���BI>��;u�$C��;S����Cjf�`�F�����EJ�ʦ䋣��D��Z�&�Du��"��R�7'���ܤ|]`���c<z��"�[+��!��繶$.۪"�V�{w��Z�2xq�$W�/-�g�h�4.{�+����ێD�������]z� (Ը�K��GWl#�������_�L���	jHb���b�q�E�8��7�K��G���a٨.�>�31�=N��C��-�J�FE_U�le�NF8(�bj�7(�M��o!���!�'ԃ��r.-����$?C�q2�U�W{�B�vn�����MU�咣�h֋���Ҟ�:�)0��JE�3���}�}�˂�zⱬ�_o���H&"ϋJ��+��Q�����7}�D<~@������*Q2���𥳪l��/AJ&�ƟƊTi�.���~�uM���$�Y��bٙ�{JL���特�G�*j���XJ���{�l@���MC�F^l�<�+��N��>d�R��)`��$���5<3�Ā��R���
��,�����k$�D/����"�|��Weʝ9�.ׁ��iљ����j�Q�mC��%iE��G�
aq��\��#u���;�wt`���FO)�]�����D�Yg��F�Ѩ�W#�gSN6�߲�]�x�s�a���m���6�ӆ��?�׷b��7��׫�m��9������E����:�^c�?�G� Z6���Dz��d.�����5א��a�6�[b
��v"(���eݴB�Z7���������q�ٛfI��r�Q�@�jH���q�?�(�/|-Z�j(�b��t?�-z�z�c�UC&�$b�H��n�]N�r���� �Ѕ���R��k�&o=]�Ww����d�4�c�D���La�'�M�����R��f�g6�߻b@gȣbM��˿����8嫬�Y��0���Y��N���>1$ܲ�2h��"�i��N��D80�@���Ϸ�B,D3�VELN= e�{VS ���4���yo�qx���t��]�[֥v#��[�9Ҷ�b�a��뿤ţT��"�j��+�X�Iӭ�8�jɴ�Uɏ0i j�,���FdzX�J�1,�̐0��*'Ņ��X(���p�_\
��q�I�|���<{���AAhG�w�{�>��~���H�m��w^T��=�1ӊ������p!��W2�^q���Ne��O,ɘ炕ب�x*�x�Vw�����R�;m�2q3δ�L��O�k�lsdf������[O�4��H��b���x���[�R�R�sl r]0�O��j�J���h���;#x�S��X�Y?~��rÆ��p��z .�����_���9%*�%��>��S$?�S�$J��F�SF�'�?ꪆ��rrX���>ŖFˡK����\�?7��i�o(�hd?x@ ^��ޢ6ǓA��̦!�a��>a�T���C��<�%�NG$�m�>��&)f�?��uꐗ�rD`E��2%�#Rj�|��x/�z�B�y�IJ�8����"8�-�W,��ʃ�Cg���Q���B��6��gUK>�Hk_�6��"�/О<������-�"-���q�ږ��0���V�C�Daf1���F�=���V��^��T���߱�8v!�a��k�IR�V��_��!������ Շɼ�SW9�iQ'���[z��Wְ'z3 y5]Ӯ�toN��P�,Jx��H[�(e��{e��'q� eg��
&փ�U�ܘ�EP`��5��UI�D,���IG�n�4��ߋ���=��ի��	>I�����Ӕ��^����jGq��(��۰��K�+�^n�?Q3�lz�u��ll���G��&�<�ϡ�*�;���թ��l.�%CB�֩���`z��}Jw�:OMtg�7y��<uC-`1��B��ә�!l��[�~�d��=E8V~�Av=��ܕ����ާc�񈫪h4f�:j�L��j����ǃ5)Ƚ��G(��$�槧I~B���7�ؚ��j^��*����O�Yd���I�d��3[\�ؽ'q3�o�#����v��'3�zLI������oh8�qS��?Qҵ�P�:�|��-#���$�a7Ǎ��ף��d�)�n�yt�{2�JŪ�fa~0@Lш�LO�i��<D!nT��ﳗ�-�w��#�T��Y���"r����r�����0�����4�������t������oKH�����ѷ��hi��ӁG�v($��ס�E�[������o�:���I5#4�c�ɹ� �5/| �5霙Ly��ib��c��K�K�v�.AyjX/_I̺���a1�3�Jn	�����M>�*ه�*�/�C)�j��UܻХ�E"��]�/�V����M|��K�P�j������i<�����(t�n��? NUH�\Z|P����Bu�5{���]�wy���)\�� ����`ߦfÎ*�q��/�Ga�@����(vxG���ͬV��d�Z)=vuT�0|uC@)�AC�F�R�*��8�Rϻ>�)@$v/)^���1cW_���	�v<��Dfx���������83�L.Qm�A=�B�߇)�H�2�P"������'�ݢUc�ΐL��Lkq^)���1f)8��a����<_���M	����w\wR��k���۽�8��kK�z,]H�O*4�g%K��"%�S���#��!@=�B�É:��`���t�N�rM�A��'���cde���"�K~��7 ��a����|J�$�b>�����bi<ދ7"�~�L���c;	�!��[�=����`�3^~�B������6XX���^��'K{t���ؖ1�F�?�f᣼��RN~��fw=���*|���Q�J,~�+M����2����ϓ��P��1���*�1��dBg%�g���\ݰ��k��j�΃�]0���@jȖ�2�x��`5`������ۭ=�GN����ga^B�8��\�O�IHzg��s�:��8}B���J�"�ŹX��&˾�y�໿�[�5,�Xwm��X\���F}#ws�����L4���&�	e���"y�fKNt�Mc�NR�-(���ZEf2D�j�4.�L|�5�<�\hQ�[�Z�򈞨���ph����ǧ7��`W�ÿ�_=�DÔy/>K���J��ۜ��-�����.x��6����{���ma�ȗXܫ�~bK�Y�+A������f&���s��X��Afc�t{��b����M�8WE)cR����]��Mu�+��(�jqmXv[V'��Ko�b`97�4��F��X\�|Hi���C˕�م;������=��C7�#�l�5{M��Y�2kH'����Swh�N�c�)0~+0�D̰��lIo�b
�/�,��:�L��pD-rX�YL�jj&
lsq~ei�a����p�TǆJd���E�k'�����Z�J��I��ۆԼtV�`���!���0:p<I�֑9ܣ�a��h*j8j�]Hk�7�*W���&׫��v]�ڤ�)oQU��������[��X�v�J��9J$�o��}c�`L�Z�NX���*u�68�-[�%�-����LG�E3M^���m����J��}���jSc���KB�����3�*jE� ��)�[��M�;��r]��Mv�M�K������na�o�#�Ĺ�ѷ���q��n�O�Hc��v1x	�q���v �(�h� �N��Nx}��"��"e�@�2E��/��e��*�4`(pz��ُ8z����Dw�#}�����M'{�p��5���7*�Z{N�&x�wOi�Ѻ}��+���NX�X�F���u]"�nU�}�km簼=<6���Ү�h.͏��St��m3��F	���g����ۘPXst�~�l�R3�i�<B���ܴ�.����H�%��8*�v���y��^kgj���}���pڙ�R(�������A�ۚE�� -, ,�H��; ��s�4>�US��Е�ɧ�D���4��Eƥ���0��C:��na�"�5�@�b-$���IŽ,N���~,��pk'��?˰���6�'��YD��q�%�Z默&��L���=$� (�6�M͉�u���@_q �-^�h��c|�/��=B�$K�N3bi�>>�V�|��ǽ�a�$~#�:e���:K�t2��+�Z;⛔s��e0T�/��z��7�x$�`%�%���5���s�_�*	x\\��0��C:I�d� ȖL
X@��`��F��e��r�q5�b���
b0��u&J���'O�Ԣ������9[�8�eay�	N V?<�w
wB����;Ć�������L���a��Ū��ϳ�*Ht�U��/�&�YK�hf��AG +�f�m�P�?��`@��Ef`��kP���?8=�nj:V4X�ZܹT,�A?� ͊��K_�'�0��U-���A������_b�#|o����3���@���r�,�ŵ��q7��	����\5]9�>Jed*�t?����(ڼ��W���<{}�%9��,�.�mn�7W�F���r�*����eǔ�c2� ��܎��&�%	W�}5[x��bxz)�<����|h��Y����"ԐDR��9�e� ���
�����_�#PF4:�.�l�6��/�n����7���	<&��C�LuL("�1m��q�Z�zЎ/�� �)+A1�Y���v��
J�)�-֪�7��n�Q�U�Mw~�:�y�6a��fE���.7������e|����oH��lK�|� X�(r��d��yy|WM� ��:�h3���[��R�g�bm0�f�*Odu�	)�AE���H?;����&��~s筠C�,߲�v�焋�/�`�����&��ח����/AN���\�4�AW��<sӴƧ"y�Z��d8����ڏ=�a���5�x�h«kp�b��"�=�\��v���X�`1V7I���t^�;ݾ�Ͱa�G�Q����հ[�8�zL��L��j�
����6#>Ҡ�Z?k�S��@���2�K�R���8�:����A�p��ǈ9��"�RW�EA�ȴ��O�6��>�W� ���m]�?V�T�?vS��^I~d��l��=.�p��8�E��@#:�$I���c4Z���� �|�yhi�Ѧ����$���]w_�副�d�|K"C-��Yb������a`�Q�#]`�|�;�ǂ�?�J!`B���Z\Q�����j�IM�v�]�3(s����^vR���ȶ�P͸!Jߢ���)Z�^�� ������oU�2� h k�cM��m�ب;�ٝ�I���0�<�DY]��= �Z�#��u3p_�RT�ia?ǈ��]0vlH�N�/�F��3��=ĥ&_.s�
N����0c����Z��C��'Vx�Օ�����\S��,�*}-5�����xLjZ��p]D`�����,��Ν�Ȩ�a�_bQ������P���t�-]w"��}2��\IQL��{9�
��ط�c)��9��7B��x\�r *��֩���o�]k[���G�����C�K]e��5����($o�df��@bV���ʦJ9�y�򏣥|[�B���'e���-�:�"!�Ա^���R>p�8V׋��m��s�O�Τ�A�x,���g�]nW�H֦�6�`P�Sy��(��������e�t�7����E���fʀ�R����"y��E�*ٲ�Β ��Z@�L���T�1��gni�����EY6�W���3I��2�� b�c���8v;k,��l��%X�ow3�����:�
ٸ'�e�/��<��>2x�7\�7}����
#;�_[%��$��3��P������pws������
P�?�n�a�p���nϝ�f��\)�,(�����C2�f�(�6�Dcٴ'��������Q5չ�5N@0"��j�#��w�g����|%�ʾ���6�������g@�?iP�Ⱥ��-0�2�����eoK]��N>y9Ӊc���c����6�[������ǋ�,'������}�����
�(B-�m�D�w����I�LJ�$��Q��L`��f�f���ˮ�5����! _C���W��B���ӣ�ZfZ���$}g�~e��}�@�"�=fg��ou֛f�)y�n�X��h�#���hv�E�Cv����֎�[ECd�-�,�}¹}ǐN+��j'9�>�zZz}��1J��֘k��a�`O��3P2³,��cy��h�Q�b�K���D��;�؛/�'�o�G��yP��?�7�g��I��r�{�p�c�-���F�c>;sZg��	����y��2���R���c'�'��뿒�4!H��,Jy�Zk�J�.�]�
!ޓK��z ���}X�Y�ڪ����F��Ϙk�"��"�ZP�k��Y`�C��&�V����fhKRx�Z�5�V�̚.�;I���Q��8e@mw�ǂ��9�3��j�i���׻1Ʈ��F�z�euźV#�^�s+�]��5�l�4�r�O��U��n�!�aA�"u5� �zo��^�sVՃx�W����V,�j?���A�hj�؊7~(��я9l�x���=6wԍm��4�>/��+Wf{1qf��w��b6�m�Dp���4_�t�J]��#�p��cGM�~��ٌ�̝~Ol�}6�!��{]������Ϲ~����I6�LYϐr��b~�&'V��gס66�̜�R�޹��婰_�("A[
�)��z���VO���Б	��,�^��5�VXSz.���/�1���ȫ�XM=օ(i=��?�҂g�T٩TЉ�`K�f�W���S�����a�F�\ ���)�}#:YJ��G>&7pSw��dc�'��3��a�w#j��4� ��t�+�^Hm�a�^A�D�����I��hN	�c���x����ʜ����ؚ���g��1!��+ː3Y����Y���e��\z|�pvQ�!X��1'F=�2S�H������
��8������m����H��b�q�T�~r��b?���p��"��Z*-)�݈>��" ���D﵍��gTwS���Lb{� U��)�h�U����!a2{�9V�7H��6�dr��z�a��D�O�Chѝ�~�Ȳ�����]o}����s�,��(��y����{t�̞�UB巙�@�E��?_w��c�v�u�ա��	��K�E?7�IEaS�ң]%O�g�bCV��$�$Ӛ���lh��� C"/HP�W�35��1�������䷺��>$�c�5�q\.���gȂ�'�B�������j��_���������P��	�p�Kduo���8r,�9�e̡��7m����Y��@���F�	eL��B��p��l5���M�:fsf�q�_8��`�#��p��H"�0�r#c�GE2����I�$fx�Ϊh��K�CO�TH�kX�0e+���e��ݩ�4jR�g���˩k��ʑ���\���z�@ħOy���?y�qyV׍��Ι�fg�8�Z=d?�>$5mD�1��Ǎ���/5O�1��������ߘ�
bY4w�V������AZ �}Z��og� 
�XL��Lw;�$���2o��m�&{.�b�W�ޭxw2yA��˸��\y���!q6KVb9 �7�eh���M���� &	"P���R�DI��ӷ�%o]N"�Űe��� h@���M{��Tn����ǎ�Y������f�glI/U�Z�p��#�,�`���:&���W]]O�x��v�����zǧ����svkh�62�͒8q����~�=�V����%��V�
�hX���U���\b�t��p���X)���Wl�JB�(m��Y�d?AxI*¦%~�ԇ�K�4s�ц��ih���@D)��f�I���77�}h�YA�d�Y�Xtk���;���㋧=��ы,�GI�G����\<����7ZN�+�ܝ[��pV��+^ߪ^��t闑ظ��{4������n�ׇ�WL,�5�{�Fh�U�H���y@|����w`z�D��ˈ}����Dh��̨�D�X��}����Y��ȁ�V8п��ҲU7�+�K\����e֠_������0�)9�Xe��%��w���X��۟�-G�p|�R����m3�