��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0&Y�y�OX�GK�!���%V"7O��r<"p���6���	�e�MS��"+ qn���gØAld4�!��D��:����+G���5�S��d{�G����c��4E��/&K��ۮXXYB��ɓE�$�
Q�0Y?�@X�<g6qӘ+�K��u^��ַ�'j��1pP=�Y�{n��Aܺ#�<Q�t���#Mξ�2TR� �m���XE�w����}%̚Qo�0���2�~��c�o_wL� �x_����e�k62�v��d�����z�: 7!�g�ەiL��f��	��M�y�-Kh��1��x^�b�cVE���;W�3kw,�5�3�ۧ`2Wf��OrP���y ��d�v%��y�&�t_@�dj�6,jh6�b3	�[�_��8��&����Q.��"�%�?!Q�)5�CU�3��1t�sB�mq�4'�����~�e�'����u�kO�|UZT��(QA^�0�9ns�����K>u�]7ͯUCp���r�r*:d�B��HN�d֩Q�{T����x��W�i�=:oe��Մ"�bJ�6&E�����-{p̅�WSG�wjIV7b9�|TF�Q��%��kùR���=zwZ���у8}e0"&	%��.X�����T'���0%��b��v�*؊�=�E/����aA�<f��@w!�	L?�yج�N�C������Ғ��(��M��7)��W����Much�x����>'��P^�*�s�qxV�9m���AM\�#�?�N)w��> F�缌ǵ"Q��-TrH�oV�2�1�4A�.t˃J���4�������6�E��3��W�2��((($w�}�Nr�э�$� ߷�aB��}��Z�!�/j�v����0�V�H��7��r?o�C�����tA����t��f�ǡ[2P�4���>�7�u$��\��(a`1I$2^���l.y��ޝF���&�e�q&��G���y�����˚����L���Sj���0��v9�&,�2U����_���T�&�I)��}�,0��1($�}yMsb!*��������Q��r�$:�x�*�q�H-I���W�u�C�G�y�-GP�O����n�y4#��ݣzq@��Y2�{tt�Ml�gk��4��-�a{`]^�7�xşTjM����t�tZK!&��-��5��V�����tp����*a���5�H� %����)���GpA�8^���"���1]�)C2��/�i�7J��b��!���h�}+8(�G��}�����9!�Ⅷґ��)���e����P~f@+G�/�IW�ի�w�"t�Tc^^����p}eT�����)���Ew���{76ʂZ��w@�/.��@�ҁ���]��|�'���ɲ]Hk*��X��Rt' �]�pE_S�����f��w�&�{xڲ������>2] ��Ĩ�cg.C�(����Aj�/&�3��f�_[W3ẛ:{]�_�}Gr?c�u�p����[%1ʻP��p�7!��]��f=ec2Pq"
��Y,+�T��s1��ڼ�� ��T:}3�
���z�]u��vQ�<<��٤��`T�wSha$��r5sì	���a�QflO��*�(o[~ln� &]W���٥��-㔾$�ג���e�V�@)�N�DZk�J/#��\K:9��F� _L��1Sl�A�Һ��`�Ĝ�O�=�,qRj���BF'���n�ȸ�{��|�j�:�e�	c���\���	(=���Q���#��z���
���%�n_�;�~dӒ����E5FgW�%�cV�(i�M�Z�<��*75*!������q������Y�嫄�p�\��S!Lg��Uo ����i?<��w�HXO�~-�Z^��m��3@v���Li;���=�?E`��M	��:��ŠtD!��N���˒�P��bn��?����{��GU4�	HU�=mG�╫0xg�K��D��y)^��w������d�2�s㬠|:�[����PIV%c�ɵ��#x�����ŸE`]��2������+r�������ϡ[�zR�wq>���L���,:$&V,ӕ�H	G)����:��m��9j\&��n�ӳ	(�d�	�~omp>�5ݟtZ1>:f��.6��&5�W˴ g�˱�����L�q0��mr"����ob�p.ir�$���}9�x}� �hv���E�j��A4(�^�[s��$��%:�a;�����\J�������>�V�@xjVPg0���Pԩ�'�lZ<��'a����z)2���9>�쟕��<��x<��7o��0xw?v|�j��s�12��S�`?z����'�	]&2�����*3`y���R=�U��R�4X6������
T��fc�+�W�l��ՙ-�gIQ7��,7�_j�Ӯ�,I��2|g̋V�>�ڷjm� *�أ'���:��ȬwF�c��{@-[�s����_�H�e��T�8&je��V��Zc
V����sX�hCTt̨?�: ��S�|�"q�����9�������BfA<�8)�;Ő��d&���ƿ�V�rL��o��X�훻�ZֲJ�,vfy��)]%��ÉY��, hB"�+T����'E�/�v�yc�<�i�����H?gĄ;^��
+�B��\�gS´r}�f��:� �GX様������Tq��糑��-��F�#}X�f;C5�	�Gٿn[ �"��o ��%��� 8�/&U�2�R���Pm[d(Aډ㷛%l�h�zr)N+S�@;�4"��»��|����B�)���7b��I�ӌV[�^[rt�Y�])�!5�GX�7o�����D1�k�("C�@��)�����3j%:"Z��-��$�Ћ�Lm�vlJاR���������3~�5nhN�)��q�~�U}���f���\J4nO��j���8��4�A����s?� y1��B�0��I�]�����H�<����7���] �����r˿|�Gf|� @��Ki�ٜ\fn+F�t�)����+�3ԁb����&�6S.�,�%i�1WH�D��-|"Wf��s�K��.f��-�"Q���� @m�-k,K,�/�
_��/7��e�.�a�Z]]Rj{�AG�����+��������1` ��d����Sc /R����0����44
qb΅6�W��������g1������'/!�X~�3���Nxg��3�p]g��������ˊv�|�N���B��\ ��:�x҉@�jX��[|K�����Z���������ꛩ��vM����d��n��dJ�Qot�p�1x�s\������78�p#\��2?E�r�L�P^��X�� C�ͽ�  J�2���G���ĥ �,�,���@j��� mT��o�<@\(
�Fvk�&pO�άc8�t�*���?4zCaDF�˩}��T_�&�5�;�3�Z�|���%��U�t=��8�5뢓$m� 5�i6�v�Y�Z(gϽ0@�ɓ���CV۴h��;8�`K��{_�@{��B%M��fʍۂSJ��4�}?����p����U��ٯ�Ra�W�~/S��s*S�4�p$^���dRF��s^*�d9���Uz�^:���{���@~��ra�)º�(q���Ѷg��M�9b3�T̬���H� Sa���9�d��"�y�C���'S`$��<D�2�5����vň?E��0����D�y�4	�����Uā�^�2� ��G���7>�1�o�������x9��]̓C�9������:�����P_Ϡ�t�$C&�n�[��aPB��qL���A��iҡ���XB��Է��A�t���8
�ե�k4b�Ʒ���H�&>���.D4G"���=YA>:$Q�3�9PS�	S,��䱻o��
q����^���B��{_��~�flUYq{yT&�w�Jh�:ߣ*ڀe�_��݊�4@��zԒ��hf�3l>��5���.�������A�%��(�Q?q��D:y-����/�Zږ�U� ��9o�.p��q��Q�����D��u����"N�o�B{����%��h�љ��i�TK\嶺���$�,�8q*N���p�d� L$�0~Ƕ��sI��EU	E�'XA�Wȫ�$�����!
R2����*[z0��dG�A�ǚ�Tɿ��7�w�e�|U��X��{^O��Ǔ�!�H���6:�6<u�;�=60�V�_�fm;�E�cnಡz�3�k���v���g�n��ɩiW�o�����=�T�ۚB��{L�?�ý���F��q�d<i��s����I��"���4�P��uR��=-����z|	h,���n+��_O�~�jH_G]�c�Nr_ N����j�^��C%Ic�8�^8�U�^��!�5�uha��׬8�m������6H��M��7��ߑ��Jʎ(Y�nX��S����޽��|���&��x���TOs�6��%JB�<�2T6�������3�\�ܱ3��J'�g���?���D�Ǟ�M�ӂ �"�J�g�����%������ڊ�}����u*�GS+Ǳ�I,P��p�����c��+7�/lw\����<��={<�$��<�{'LC���@ef�Rގ��Y�EΜѽ~e�~/���	�CQ�L�y5Y��s�Y8��/�QmJh|��:I�`ZG-�3b��M�Z:\r�>	�h��ȵ}�l�� }�TQG]�T�v�c4f�o'�6�[�T���
@�#zL_[����0��=s�������������t���eX��($�1���|_����lw��0����К���]�w�F�]�lh��2��kΕ3���VD�K쳃��rj(�����k�+CdJ�.���&G��o)�}ݤ�}�-�$�̲�㉱�,W�Zjl�Zr@�Xt{V���u�?oaV��*a��8�$���{���r���A����j۠7|�?���Sˬ��s�?�~�8�u2>��aD�m�GV��Is�_����֜f�/�Hz'D�tk�bLOe@�{�S<�y?E��[���B�^��^+�ō��@����Ϋ �%��ؘNx�?��wܨ����ˑHmP4T�N���k��r�+xa��*/�m 0N�pT�k���ѳ�C�!��BF??`@BOi�<9���
ޅ�a�U]��v��+�ڶ��qN�F�)�؉�p�?Y��ؚ;��r������c ��0?^�����B'͹�L޿����רm�S���ŵ����ڦ?�Ȁ�T�W���m����-ͯ���g�\���4�2��3�P�X�_�Cش�!�n���8~~�18.���w�%� ۰c���yO#�р���G7�nY|�K�a��`�,�$�}�0��I��v�
ޓ�oT!��yS�I���Ӣ?�����9�oZ�?�2IX'a�~���)	�@����Y�5}=��Ֆ.��Wk��P�>����EMu���MT�i�������L�����%w���@K�X�ǚ���Ϝ����dX!;KBZ6��f8ؔ?Y<]�y�|7�V#ä������O/<����և-
��~9�^x���A`�;Ni���D^����T�O�.i�҂��;�c���^�P'9&�nW�SZ�/<kVk���6��}��7�v��T�J�����P>�(��z��vM ����ܳe� ��4��9�?�����'�d�^1-Ň~͘���[���H��|J$��`�ݞ�mZbTZ��5�e�ZY��x��Nd,[�Ƀ�<I5�Ũ*ކf�Ş��#����Y$�Rj��g*��#2Qא��Z��}0����ƙ�Fd�q4�����B� 
ٻ����߂YX1�M���AH5:�u `KX���gP��mq��N�V_PR�zi���;\Jf޵1�u7wD�Z�v�#̀]q^��������ڟB�w��;zt�K�l�ri����71y��C=5�1�ͼ00)���"�p*?�B��c)��>rc��W�� �}ȧ&�k��G�������������;�+]=�M��!�|
��Jc�0ϙ,��#�X��wP+ʷ���?���UK]%I����jg��E�`f3Gwf��X�����
u0B{�0�'mDP҆!B�
��5>bnT��9?��izo Xb<��.(�m�C/���{+r��|�0�2(�5����*8��8>����痑R�[���OB�|�%*V�����Rx!p��fJ�)@�^�Ӱ1ĵ^{����r��{���]J:�Y!�Q�
�(�-���Ro��p$I�oﲒ��t���1r� ���P���>���@`�?�/�]N|�z���ևQ%��a�	�TbQi7�G[����b���*{,������e��S��	Tx�G��Z:��x!��z�!-����y��bxlʢ�����}2.���@@&�'�3v�3*M۵Qr���8����)���F����h#�2�+HX��/qՠ$h	�}=M�1?U��7VM��a8=�q;Y�e�&�/<T��%�39�/�x�?Kj�A�'xL~S�A�4}$�\r��8�o1�@k�}t�[�{.�9�#��j�J?���������_��%i�_Z5%0�Y���lTGb�ƶ�����W�B�cz^+��T� A�����C�����&2�ğcm�ם����L)�D�F��Ƹ�%5��}[�'}�!��6�삊C���zA�F�9��|�'���2�i�$^�롷�S}��:DQ*#_h������8�B�֦���-D,��"l���� �Z�D�n;}��x/���rVp�l���������˅�"}Ȱ�zڳK��v���bA]�~Ӊij��[�qoȓ���B3�����@V���;�UѮ��Ȃ{%�z��K)*mj�����\إl�̜�z[����)H�����ٲ�.u�����1&�J�"�.h��D�j�4��WK�7�#�q`(���#�OU/U�c=���}�>�M�N�dagg�}���^�aF�S��)���Afh��%Ar|;�*@��j6U�k1@"/ǒ�陨-��n:YT��]Z��Ab`�W3��s L5<9�$9�_	)i�K�Ek��z��x�ӏ��dr��ǵ4&U)��B��o��Ʒ�%u�#/��n��Q�nyTa/J�-��u���$��ܤ����_���u�gnXM)�`����$HE���ٴl��#(̺;M�`�Q҆�P��4���~����٧�ω��@h$��0����MJ�aLme�/��@'����5��Z�J�����=d�X��&��C�i6s�vݨA"�a��D��	b�Pm�v�XJ�+�1W�P�鍦a�]��1��hb�\;�Cub�M`~���;0!�p3��!�:�����&�J�ۇȯ�ܾ�I����dW4m��f�H�����h��zN��\�]��"��q��X�Ő��%�6[���5��b��V��T0{�R�����z���]�j-�|����b��u���-��I��`8�5�m�r��=@&Z��9Sp��j-ezH�}��X���(�e��s��E���-\Hj	&ѡ���r��ٻf���w#�c�/�3��P,���'�]��/�Žħ>k:e�h�x����Z�M�ax�V5+��w�k��/���;7m������->11嗍QXzIr�H�}h�w�l��6�Y����8���Ӕ����P:
.j,0����J?�S4���M���i>?'�Bg�"�#΁��5�0�r�:_g�:��}|�($�p%������}���|,Yi�0��(/�.�?Ȏ��OE��\	I�$^q���Q��n�/��^Jf����Ts��aގ��6EM�W�� �+_����룍�)�9t��d4��͙�nƫ���=��*f@�BS-�����bd:?3�$�|��cۭV��N2# /(��n�^��gY3m5Y��'� RB ��<=�,i�GC)���f�����x�h����{���J���y�+߀w��η��<
x��w�iTp��D���?"r��,!�C���-m5W�L$=	��1Mc��6�,�CKɍz:y�J��7AXo6�i�/�M�jDCý����{s.I4�J}M�B����˹>�?�n��M��ZS҅�&�ӳ�KO��8��k��7<:ҥ�,kagl��I�]����Z�dUUi����*�'������W�I�91!A��=��~��,�1���?�Yc�i�dG����G��o��$?��`Hru{� P&@��G�U%�V����	k��i�ѪA�^OV���;��>vR��;��6��H�;��A�G%bK,�Ty��~%^���r�\N��+�.uoz��PN�i�[4�В=�����B�mE7r��,b��hĉV�Yl�|T�󌔝<E� �������2x�vB��Z����J��A����G�a��D�:O&����+]�����%P��gc���B<l���Q�͇!��	�(+��;�ΐ3`��Կ�]������bm��jt��T(F��w֖��kh�'챏��f��	�2�i��+��-���;�w�]?�,�v�$C�d�V�y��q �4���`&���%�'��P�ul�mW���6A��m|�4�6���!��Q``I&|��fjP��u;�p`�HA[�S��	�d����%jC�Е�7��K틈�t;~����z��9W�[�<@~����w��g��=��됽��Ct?'����vv�d�Y]�(��u �me����q�M���P->��$a���P����UB��🻧�/���&/Ǯ9+�\��W��(f˸|���
�g��Ь�0|N쏷�<��Hmv.ﱩc�nq��_m;�҂�we���fM.Ae� ?���g3ò2��c34��}�UHB�֗%_�Ʉڗ9ٮ��2_��z@b���[,]d�� ����ϭ�o���t��4� 	�	�I®�,Qwt�1�vy�`�^5�pɔ0��"Ұ ?�yv���b3��\�W{��?:|��n�@��I.��e*}�L3�ϒ6�
|U �m{��01=��N�t�Q+�ǎt���y�W�v ��4�_��H�T���㑑E��8-4�z>��"d�%gq{�xֱ�nR�T)|LX�hh�=��٬wO�_��M����,����W�]�E�.eݡ�<��N�`#谌���_#Z_�����=��G%�܂��ن^҂��-��Z�i~�w1��J����hHa��
�?�D��W/܈��A��Ook�S�t��,�n�>��# \Z���L�n<�=♒NTꈦ�`���9i�.#+T���9M�����/��_�w�/i�e��$�0�1��sA��h'�/O��^Y��~j�,��fL���]�i��WG �����Bc��T3��j"X��M�W��n<�"�qƣ��8���E�Q>^+e���`�O2��[�4��q�6rҡ�k0�����`I���])o7�p�D�!)O��k�t�Q�6e�dˀt��>Ψ
��y��Z���=���@Q��Ǻ'3敭��z����2����k�w�#h���t�;���  *��P���|��|����U�2)�4�f��@��e�a�Ų�82����t-��U"6;���A,G������$S��MC�J�d�W�0��Z�1�՜__��sj�����!�*MϞH���T΄z\l�M�K
�z�$���$L��y��sz���d�� �1I���@#ru�ͬ���D5��X���u�m���x�t���*���yz
�p��\�ӫVh챣f2shm���d�J����̑�m��\a���3W6��%�o<��o͹d�0�pin�R���"up��K��<7#����c�ʚ6SK?|�ϼ�vs�'�+;�<	�o��5ў���pҠ�P�r���	D�Y�w�� U&���%��ty��f_�o[�tw�����	�;����c1r�
���gaނ��A�><�+�Ks��;�X���+vQ���s�&u�T'_�T�р�i�|�k�P�7� �I�����b��H?6O�<]/���[�*t8��'5� ������n�o@��2��ҁ�%���E G�鳥ą"7N�R{^�L�X�U~x���Oe@Q��+�ɳ/#z�*�ӛ�*��#���O����e�\*߄6�X���ۉ˃��ں�E��r���aoF2�����Z?\)U��'7��I�3{8��	�y���� lҌ ����/$4�n(Y�0`����}���U��$b��L U�&L�yXnz�vY�P�trpǠR���F��rZiHr���5-4�e�Kݾ2�]
��C�`�x��9�د<�,g��J����V'��c����Eq�����t�f���h�Im�[f���/����#�v��r��PRg��w� ��=~{�|���&_>�⳷՚���7�t�[���a�����5��R�щHϵ�'�������w��xuo�iHy	[�*������ui#!b�t �Ĭ)l�B�Bù=j�fZ��uwQ-��_8�6�;�}��(%��=O�Z�qU�6�3��4�� �^h������;x�f�<��CcB�ѯ�Q)s����f��a�r!A�=,6�ܽw����j��ި�G����ƾ��+��"$Zȧ-��u�ßC,��b::�j�kN�F�!��\ZY�=�w�ke���A��|�?(�+�f��}����;��I	�	��v�����4ϤT��&8��\�����j,ʩ/�Pc��-(��z��k;N�\Y�nNV9�饣=ػc�S5���ʂV�ߒX� �d���('�a��H��xӌ�ؑ��@�q<�ӹ�rǖTkMe��T6ek➣�(���|s�G���A����a��ފ��y ,H���㰔�x�k'�KQ��_���t��I�< /[�Qdw�+��4�1_y̻�$V��,�YL�z�},�E�_(������i��l����b)d�Q�|�(������cS�;W6������á�y.kL�}�����.�.]�K���V�Q���v�D�y�e4w'w�\i�Ӛ�bP�@\Qe�[�WiWo{�G�j���ǽJ���pr��j�Vu�!�{�ɹv���e�����4gB؍X�bto��͠���@x��gJ2x�kK���.1Q�5���UO�ȯ�U�g$������	�VC*�IQ��{QfŎ����n�nR�5*O�(?��$��n��c�H0�r��[�&�/!�?ʴk�)����2��G�vLp�M~���
�������^U`�mb(�\UDՄ�*ܹ̭�
B��0��)�N���@�G1�M�O���n�yc<�;��ۯf��L4�~O,�˂��bB3���:�$��t*$I��
�{d�̛���7�ob�7�n>0K哊6&K�TB�kK@.�/>�����KT���𔋥^e���!���ώ����F�&�ݟ�C��2����?B�{Gp0�|�nʱ�8́��l�s֧�t���
�uB�/�R !�t�0 s��݉���`���f��O�͒4>GB~�r����3v�{��+���X?8N�!1�`o�sNB_���5�_��h�NV"E�+��M��`bN��}�`)�=�y�Q�O��`H���<s&1_Uz`E�ڦ�ſ�z�kY�?gǀf�XL�aa0���ݐ�$���XRV1�lE���Mcp RJh��Cԁ �L&�e���X���Gdh�F�{�\��fԏ y�i�ǫ3h��,�Gn��}��H%��[{��`�nE�<�����������G����=��	����"��ͽ�>WG��Qfq]���r#vg������qʸ%*m�1�%��D^{�BG� g��do�s�Ef�{Sv�*���;@L�Z���νztWw5�MF�&����#uE/�A�"�&	!L-t?���f<),^����j�5���Ć��.�.����7
��C	<6?N�>S�c���&������`7RU�
b�}t!/���l�XZ/e�����=9���W�����pƤ��{(A�~]�!B~�;�_0�U'ϰ�mux�v�G�]��7qg�uR8�-a��*�띞�L=w�qz���`ǩL��ĩ	O\4[0RY�]f������T����65��\b�tgq��{�̀U�N�阼�33mO�]�m%%M��-!W�/��{�㔵/��t�~��lրH
J�bN���\������Lĉ5�l��}��`@�fR�x@#�{W(�鵚0���n��2�3+��ܘ,T��������_M�rJ��]-�����ˮ	ÀW���<��@�L\�f�+uS��V�n�sV�DDG�nK�u.���?z,R�6��m��V�ȃ@?�p�w��I�0>*��vOziZ�z�Qe�C��i�>�8\�Yk�4nv5ڡ�dU������c��{�8k���
7�V(aM�<���s�"S�qh�\�5���i����
Sj��"�Pih�����[�Z��	/�/$bo��H겲S�%{���x�E�D�v8�G奱�]�.n�Ks}�C��Ꝯ�,�C��H���*gؑ?�+T�}zL��hlWL\&�+����.�ɚ���gH�Y��Ĩ@Qg��e0;�za���z'��BK5}�;l3�l4F����[�D�y��y>�	�A�u���"*���;1W�ٖ)-r��mesK�S���z�a��9 �����Lo�P�i����ag�f�o<�@3hюE����t��~�}F���.D_9W=-kM�>��6��ӑ�H@�B��S�Q�%c]U��������8{'���t��z�LW{���i�M�j��1*��3���o0֭1K�&p�@Cd=8���@ֵ'�{��7N���	�l(�Z׼0�i����S�o��:\�rj>��W����w�I5A�ԇútz�-�T0�ە��L���.IV�%D8��\��uOg���m��ڽ�T�w��ǲW�8J
�zc�z�W7*���uEԇ�E�Q��L������d��V�V�����m�2͎Z�+�y�ƭNY��p�;*'���Ⱥf�����Uf2!�IK�_��k�͸�x8��3FL�<w�Sk�� ��O�7>���� ���*�d��ß���uc�4J��3d�-�����,�}��~��C)M���w�o\(!8�qd���]L��a��jxhH��a%�VH�8��� �ez�@{v܄7�C������z-�X���%ք��<+���,����������i������;�_�/'��ao)���~��3���!�"��J��D^�	T�y@���f�(�ԡ{����.���u�y�IGl�kJi��r�7fG*h5��"��(֭��W�/�q��Lۀ=$�g�~��;-��3�u��r�H���vD���H'��m�S?s�B�7aS�J���\S�L$֩(�Q���m�i8)�sJ��E����o�d�1�02��T1Fp�JR63�l���S��#�bjF�D_ؠ���KO�waN^��0�| ���(�����"*� ��5�g$���."�[�K0{ZI�j5*�:�O�v����GM ���mT����=����=s�Ե9��nN������b2���:�A�Qf��}���X6�MnG0���!���a=���°Lq����͘������B��w$��e�sIs�I1ڧI�C�mE�	i룃*��F�6��d-�eG���h������ �&>��'φ��PSzFE=*͈W�c�3B��.qF�6�g�R�!Nf=�_OڹQ�_I�Tԏ��� ֔�P�Rⵛ`�3��H��rix��u5�B[��N�u����^|��I#a8�ƺ��}�)�
��+m�t$��9��7�x�>���W�t-dbR7���p{�ǊA�~/�ᣜ����ŦAJs��iJj��"��܅˻�V �A\s������d�����2�D�P����´ʆW\&y��Z(�ö9՛����B�bd����6kE}`DL��ð}	��s�z^:B����`�!s[���d�#�9Uw+�|�I�4���5d����*?X���R���c\5���=���Xe�":�
�n�'�女gN�3Ne��#�識����Ѐ�������Փr`��)�X�Jjqz4*�4���6�@f}}�W�q��'��'��qAܬ�?�&�.tB�3�lɨ�89t:�|�#�d�'���kQ|�J��|Ӵ�x�R�ׯ&Q��C���q��7�1�KZ=�T���d�r�qt$�{�-#+���yӝv�K�0J��҆BBu�.P!؛$�S��]X��c�⡓�g$r���3�8��8���M�a�d9��S_K���4��&�ڱgl�i9�� l�u�;�Z���4 F\^�]����N����_*�~w�h�%)"��w0̓q��ė5R�x�U�q��}��p��"��Ē���-�"�|Z�&a����s(k"��.��^��X)�z�X�qr���w�OV����� ����
̧����K�V���R���A��r�(�������ǘ��v���A��5�{L1��VV�,��-J�ddt|�{�ڱ���Έ�ܵʃ�L9�$�3��F\�-:��	�k"��w&��,�r�d=��p��q��~�m����U��+�L�O�ef#�hgW�������96؀���}Ϛ�9P�r[��B���%���Z���0;)'�+���ۙ�7�� ��t+��6����2�4�ȁ�]4�%�䳣�q�3�ɚ���9�;oPI��3�,��|��vʯ3q3���ƆH�4�t7 .���'��v���W�78�ƙP��[�lD��W��zU������7�@��l��=����5�a�8������6S��!�>b� T֬��s˥�@�p;~^c١�Ä�$%8g�:�n�H�̠H�kn'G�5J�A����*�u�:�=����~���b��r~�^��V?��%�����8vcQL���N�m+Z~��ͬ�O�
ʑ(`�Ͼ~]e������64"0ZsQ������z�.�~� ρj�a��E��<�0UO�߻Fk 'N2�w�"RX7xUNa�����
���j����%O�_A~$�k�����3�Ƶ�W���ڲL��'�� :�z�K^��2�t P�?��1�^9���B�Zf8��i~ʭwg�����HXkn��H|G���;�5�bU��̄o>���{����)j��oSY��(�J��x����b>�Tn̆L~C�=�>����'�Z;�����w��$	�q_��.fm��aӞ�o���a�����bi�j�yl �(*'?��)7��c���f�������7K���Wk������Ͷ p�y�]�h������KL9]ZFD�,��������S��_��Du?��F*g�o�t���nM9T/�,(.;��]�Ӣ���T���]<~����{��Buk�n���1`X�Nv��ڌ�d�M�b+,O��%qa����8������2]e3>�8�ደ\��YdS'*�ʪ���$ޱ(�Cʥ��q'�ˑ����\}\
B�Wx�#������φ+��1B`�G�)�Q�Euv�X뽿(-��2�m��(�3�i�n=�a�v�o��׌u5��|{����1r�2��
~�ʩ�FWOqD�T?ĭ'K�9D�R�8���z9�]98#n����}����q3G�� �V��W>�P���������hP�N���\�[Sp��kFx�N)u!8n�/w�93�G��˲T���)������$
�G�缑K�y^�6]��g��7�����E���<����(�~q�n*�7$|\L���[��F�|�)r��4��QӃ�T�ˉ��t7`M 8��ұ."�0m�ȯӄŒ��B����<J�K�*E��.J�u����)6�8tOt.���) Px�V7M�n����g�M��lK���fP�����BҚ\?��5��P�2�K�O$��D:�����̌T���?�l���rY�`�%\TJ��GJ�r����>�o)8#��?0<
�T*���k7���3���y��?(�p�F]+V�o�-f֪��Kf���v����\䊨��N�f�Y�+�A��,uA,yw^��+ɳ�?7�����
��ĸ���7c��޿��Ww�S�	��՜�Cչ�
�����KN�^{��6#��(��U�`�c�H�y��Il��%h�	�5�i���_�9BEm�� lS0��;�(0V���
p���'����0[9��Q�*��YG
���;Uw�.hQ�2 x�Ӹ���o`���tґbaz9/+~���2��	�����J6��&h�كH\�P�+^QT��&n�`,��q�ހpS��U�7�:�Yޓ�Q�bt�0R]�GT˖�+?���	�#fssϊ����Ń�j��M"VH��!���<���Z\&��7�_T	�3?z�8�@����Y:�u��n}__P�"�Q0[o���.�PE:�毯��D�p��x̏���b�KQƷ��s8�:�AaBi��6�+��Tc�(e��{�&�?���ނE��=d��d����J}:����{N�#��ݯ�,I�)��e/	'~� ��͚�
�Fj}��ܚx���\.��OY^X��F�/b�+GlFf��R.5'����b��-ГpF!
��ʟ� v3#�.�4�o}O�
�H�y2C��m�ČB&��"��s��8p��Ŕ�����0M<��D�� �9`��m��fX��ӡ��7��I̝�͵�#����0���I��V�ճ���<Q�V�xU��Z?���yz�_N�%�G�=HȢ�(�#r�9կi�P��?������Ņ�?��	�.p�����tǾ�L2ۢ�`���C#n�q��W?Q�2����f8�8@��HF�:����gu+��
hkhn��>�M�--B�}yE!<�K��BGv����aVQ�*x��7�i՟=���jTG�n�`t���۳"�!��EFn0�j�P�|��je���D���R�!��^3��������4�x�"S�1(�P1���;��p�s�x��D�PG��p|�9�(�d�<�Pk_��Kx1$f���g&�8f�@��]��������տ��/hcG���G���CH�j[-�N�κ�|܆PL]Gwm�}�#���`��`���2���yF����ɺF^{�tΦ"	��!̮��(� W��B&<�<)FU���>���?}f+�Ss!a4a�p�v��҈�E��/�<�����G3��.�!7��?�Ͼ*�8b�]?'�#��o�V�g�0�e�����`zI>c��m{0�@����d���ӛ�$�>,nZ��7|o$_�,�ڵ�����Tƞ7���۽Ӌ$��Ѷ,���.1w����a��i�\�'j�G��|3�ݹq�B�(�J/���j݂��i"�!�x]4[������G�Mi�1$N�f<
0J�����O>-s`��&�|X�������+g��P��n��+�]m:M�?B�Z�CJ�Al�9�y8 Q�uG��q�
��C>�k��@��/��`��abz�n�C�$�����ƈ<����$��]Vm�>�A ���'}��r1h��n�q���q,���vQ�y�;_`����Jk4)bL/��y�4}��I�J���ڙ&�wݫ\;L
!5�3����O
��D�������=^�����w��qD�F��:Fp��A`P�@�.��� I"]��Q,�g��9����������5ѓQ��Od~1Q����9�_��l��<������a~f9�H݊�I&F�,)EĨZi�d�i#T�4�k�p~8h�TT��BB���ۅO�isN�Q��K\��(E�7H<iXĥn������u� 7�bV��N��Rȕ��xx��s���=��x� G�~�8MYB󳆕����pJR	�H@����WL97hҵ���r�֏'��:��P��YE��=;.v�yA��ɜ����i��y��)"d��LE�h�4��|�ް���(����;K�o��]���Z�	ͽEJ٩f=�1_ٺW�%�%��ZM�٢�$��,7E���,t_�X�}���vT��?�tp^�X	t��e)NF� �r�������"�'WLQ=�('��7��x<=�-�§`)N�� �f�
<�7�=�C�\uBN��ޖ����ΕH( ��e�>��Lk���\�R �%���v7L���wf2��g�4O)I:y-38�"�2@H
/	�}��
Z�3�R�m���)��l��\�/��	 >/��]�L�㐠h�r��t*kD���}|K'����N�OWw�z�2!��D�+��[+�ӰihN/7��PU��w.4�/�ӳ5��l�o��R��{�-!����-�*�{D4~�� &c.�����e��!a����m�T[(m�O��sYCG�Oj�������l��"w	�����w�'��V|Y`�lJQk8cHO8�����wC�F��*f]T��A��|W"�R�'�9B�]��\�DW���Tb���0ǳ =���W����OQ�ɺ��T������m���E�)���ޭi�n�˱���iZ�;>��Nr��0H�xFA�ˤj����|p�:���uٺ�m<P�C|�=}�.+�����I��!c!"2��9gƝ:l��Rq�[��X�ݞE9P��d�e@޺j��c32!:LP�A�����K(|	��D���ʋ����>�h����چ�T c.���e+7�~
����I;#y���6`��".�e�Æ&d_"��aĳR�G��-��,�R�_�Gg��W*&��}���"6��A�ό�c։W|y<$��Ș���J�cP ''��U-ST��n<_t�'���A�lʍb�F��X-��K��d�F��sW}$���Ȭ��2I���G?H�%����ȩP�K�^t�bv��!/Q����f�NDh�d�#ش�ο��%���a�g֘V���*�t�ѳ+����Τ ��sS)L(�/�5f�dy8�eiUwR��9|����)�p�sJ.&W�G�|��/�f�(��p����q���6�\�� 1_�L-lS������ t��u��ZY�@/��)	_�3�ä��'0���ji��x��oL��C$t�1���٭��������ЪC�]���dIQ�~-�=V ÿ!�Zjlb���O��1�����#�a�l���ta$�P��žTP�Z���}%c^�x���� ��`���lmQ_�I��wR��H���si'*�.���i�~J��dX��,�I��栕��Y3�����L��Ȍ���
�;٘���
8����6�Ǳ��!U�c\(���ɞ2��`��ߣOE`�b�kK6�x��/��u�_A�����g����U�@O�xM[P\�=�Z$-�֔,��c9l~1�:ĸ
kY]6&��p*�z��)	#Am͗3&��D�'��ij��~���(L�E������F�?��vj�,BZ�������gd�~%d���n����)bAsu���&�jEd����ˉ[���l�'�~�u��fT���������Hi5W�Z��CO\X�&_0o���Y�f���1����
���Q��}]�����\{������/ئ���D��h�d����3��|A�V�f8=>{�Z�[�k�1��C�Y�SD5��/$��R� ��h?��4%$��7t|�'��@i��H�n0�@qy\h��
"�,��YAD.���!Ar��z�Qk�`ρ1Q:aV���"�Mb�G��g��DoY�Π��\��\֛���=N>}�Į����qX�����9�/�.E� ���H!�HoE7(��M_v�YX//4��N����X ����)���V�Q�2�BcL�H���Wo,;;a���bvW�J.��Tɦ��H� \��QW��>};<\�#�>��6���6t��^<�q��g!�f���ŭ���`Q�v��j� ���Y)-����[�|Ng�Gli��!|�M�)t:5vD�P8wv��_�|�"֊�`;����v>�J�6��}� :h]��}ƪ$��.��Ne�wL���Ў���C�{i�T <� Y��A뎪`���wW��&���g���5x
K�������#5X��fC��t�z�����$��r����Gh.R����W�$��x�� �y^�u��Zl�R��X��<��c���4��$����+�.�!_�!�寽ξ�VW�B �m����G��=7q���Z�P�Rœ���	�Q#��оֱ/wk��X>����jU�@#�?m��H� �aQ�&f��r4t�U@m��x�[�*a�_U캉���9�sz��ǯS�g3�۬a���f/�	�O���8�&����L�O�XI9 �"C��GÅ���	�uܰ�5����R��yK[�¶������~7;w�����_�cО��"�v����v��D`�L��e\@�p�ٻi|������Ub��rm�[Nv�R�;�*lǍ��5�cBq�����)t��]H0��dQ�GtL�����&�)���,������yz��/a}ȶ��.����c�M7����.$uo��f9�����'�%�X
�KܔRk��lDf���j��f����i�w��+Ǡ���>�յ$ӂ�&& '͋&๗+V�bA)�l��9�0�܆XT"�-��L���0��т��
h)aa�� �1���H����Kz˾��E���/��\O���fF$T�O^ܴ�:��쵳�����&h���㞨�i(�Q�F.�Ձ�9��گ#�kjӗ�`E��=M�ae��o�Co)*Wx43��ҧ��	W�V>��~�0F>fjF�'��n�A���w��~A�
�=�Ѐ����{_
�w!6VϤ�!���Fz�/!�G�f��f$��V������H�3dc�WS��[l'��0�RWSp�!�d��4�ۚ��k#^�.]�ȴPl7x�%�� ,�1Zx��Q�R��FBUU7���o��k����^ ���$����i8A���=QW٦x��[6Z�D�q����ԝ�%��TKr�pUƩ��^��������rE7��ѫ�[SO�ɦ <�!P�Ѩ,(����\��z'=Bz��G�ھ�#��N�L|��y�yh���W�'͉���**r���z�������j�	�D=s�t���G���N�]�.lw���="�Ij;O��j�ntѝx���`]���:g蓎�7TF�/$�s�x������-��v����cfo�d�5�-��0��l�ٖD,��a4� a���9��̕
]�E�Z�/ ����W3�ۢ�Z
%�]�%{��8��-���b���)�2�v�ٮx�qPF��&�$̓�U��`S<t�o�7��Fn�k�Ų�q���R�JrsɄ���P� ��G��,t�o��ߌ^7�����è�Y�r�J|~!Lo/��S�w�q�]<Ѽ�?��-�,E!��0��T�3��BN~E���ߡ��_��})tq�{��Ժ��-U[�Ɯg�ns�$K)�K<1�#�x��R͠2�)�ш�9�]w�%���B�X�E��-��h���{6u"Y"4��w��gv���O�w��6xh��xIˮ�\���@�?�D�cҠh�fx����찯X��}u0ܔ�P�������&|R�'�i��ɇ������ʡ���i�~�Q�)�Eu�G�,�	Qq��`C���A�u׾��'�}Q�h;���Y�o��Y8��B�=���_��h^��������pw�y�;qBm���{Ѻ5��I�j�,��i*$�}������T͟[!)���/t�.�L�x�F�bWa�M�bc�i���G������qA+�.$Q���U��]bT}6��M���H�Xe�ZQ�?$ﱦ ��.�r#u $�A�R5`?���p]�φ�AB��\�t��f����
����&���>5U��7}��I���ӽX`i,㼬�_�a�Gy�z�{��텐�lqm�$iy_Δ��Y�C:���M�v��
xS'�J��~`��=��w U����g�l(Tzf�A^ζ�e뎞
ڃ͋�;���r�����UZߨ4��K�Bԋ� �z���%x�b.^T�|��ԛ�=��5�dQ@�W�{��*W���dkI��o+(��*0��ga�J/$���b�2f�B>�rZ��j�QT�6o�i��m�UH��8�É�:��|�7�Q&_MW�>&Cy�(2z�"��2��z.��\����3���}������m��N�ݻ8���+�
�}�.�R�Gp�K$�ۥ�6F+o!���G�!��x����>D�+��ʀ9�Ô��G��Hz�+�s)k��	a�����F3�}KL)`�w�a��e*�SA&�����-��';/^�tS<̑��$�7վħ#Iӂg	��@�Q�A��1�O���IU����WĠP����qʈb�N#��g�\%���T�ܖc�Nxд�N����⛸Ny>�(��-�)�^+4���?B��יK�{���*��ð'�Ǆx:�q�O"����0
1Fe)�]������f3\zB"��H��Ǉ���G���8�1R�T>a�h�іl�OMLm1������ǵ�8��<���C�ͥ���X���gT��j�3>��*0D#��Y�� ��S1�1)�]"��)� ��uE�֖@Ar��T �m��.��.q���I��.����Y6RV�F���c���h�	��l�����k��Î�5N,)�Z��p����������㉼~6�ܯʁX�Wl��o��2\�%��1U�Ann�\��22�����]Z�>���񭪊A��ϣ�<~��-�_�oo���/��NL�Β������L!/�w��#)pR�mQ)����ۚY�
f0ym�~�4Ȫ�o��hs}�DR��ԧ�F��ѿ���,a��*;OlT��D���+��C��� �E��nz���� :Й�6T/�����m��˒��d�޽�`��My�m��2ǭ�1픭${Qi\�D���" ʦs��2�EU��k���K]�����o8� Q
�5j���+~E�*_�3d`�����C`U�k6)�\�Q3r@$˿��F\������D�µƣJl�	c�A�թ��gv�R�vQX?�}�����$$	z�0����4�K�푆�ݾo�C��?i��a�l�mRM���N;�9� <f��#��S�|w� �=���x�J�����"<D/�҈����a���X��i��!d)B��	(�!Sǲ^t�� cY����ȣC jB��0�_�ք�݆[8��{,��͜���}��ɨ��e��q���%���J�<>ux��.�[	�Ù�B�)rE�;^����u�������^Krŗ����2)�Do-Y����Q5@��!��P�<�g�=��x�l���F��B�)B�oz-oW��V��ݹ�����/פ*�
^2��!�c9p���M�ٝU��^U�hǵZ�OZ�����7(Y��ŜE'��_�ԨF��3�M5����Q:Jv���3h']9 �IA@ ����Ia�O ΃�,D�<�}��V���_ϫ:f���t8����,��iv3y&��~�V`n#A6����O��7��@��,5��;\���!P&)�_��HV^{z���q.y�҇mz\��7_�+���h}��_j�h��<����]��+y�X�W���F���u��q��DR��Pbb��Bf�h�b�-�s9`��GGv���Vz|`a�^/�zF;g���.a�J����Z �)'�VF�a��駴<r�Lw��b���j��ej��ʇ�$?-"���Q�����+��莀��k����TLdգ�;������v�>����V'���77b�X���c��!��r֐!n)�� �=˾q��c����ޖ��0��Zw0+&�3�Q_�;���*��L���Y` At��[V5,�6.�{�+wLs��g#y�7lZ�+d���� ��� Vu1W��K_�R�Q{ܲ���*ox��F�J�z+˾h$�;��W�1}�dy����lʐ�,/�g�h��Z�<x6�N�ǥ��+U�����m6���hp_�8Z�)��5�T�9/~oa.G����V��[��{kMϹ����s�gA׈Y�z<`ꙤU����Ay���=V��wӪ�Y3�pO`�_���K�Y�H�'e��=���y5x�l�`[`��g�i���!���z�����rG6���e�0���k}�#D����iR��c�����9�A�N�EE%9��+`��
ń����2y1�LՔ�@�.�����:�*�����l���u���udJ,�V�zsYaۈKKmW��mK��>U|
���J�W�O�E�6-xXb/�;��:o|��_w��q�H�<�b�òH��1�$�tY�^0\Ey���7$��$�A���%�9���`�TT����n��Ϥ;s��|���]G�P���{h�ʳN��R��#��! ����Y^mQ[~Z#5�!L#z� M,TRPL��=ӏ���P�/`��T�).R��מc]�E��:���'+	(q5�J�*�A��G/�����$~���'*�EQSǯ�Gq��c��б[ ��D
!��ݰ-dXQ���v�� 8!_˹M�cNn+��������V`�i��'�.f���V����|�VT
^�Ё���g���'��2r��S9{q*�)G�EG��m0@��)�u}���܊oU ��k�f޲�L�дG;�
�(���G�_9+�$g�|Zr�����V8���<σE��f 7��8b����?��1^�����Q�D�4�q�v_D1�Y1�
҂�X2g�@���J�D׳Oo�ٶ1��'J,h%�C��q3ܯUU�$y�8�q1��r����06-q�����3��,��zȂ��L�p���i���jё�%�S6M@5�Q�-��buC�A�Mpi���OFͺ�uu�jc�Vx���D��-�ӪulR�)��gk�R�3�����Ę�#�L�3���c;�i�\��C6�d¥��}F��IN���L��c�W�~y<a�,�|�{b�C2�>�7F+<jb���	�痢�	� _k�R�͘�%��m$^�����S�|V�u�wc�L�<���rg�q�RPF�H�**`��� UQ����A;j�x�q6�1��)�����r;GL~)#�*������}M�\O�X�G#i]v:���*Å���W�A�)�����`xW���E��M*h��E���#�&M��Kr������܂����d�ۭ���Od����l��-���}�پ�8�?��9Y�TP��?��&b?]e�%?���T�Yaϰ��@C�6��c>��W�&��j�r³r�f2%WU n�D�˛��^�I�c:���[�Ͽ4�
����q9 ʍ�Wu���K�}d���Û�C�{$hU(Z��@�

���Ӧ
*�cw��6���י�ko,Ir�ɱq����阀����v�_�@��},s�(���R�ںxA�2���`ӸT����ҺI��g,[?=۾D�[�	���s�E��5	�����К��k����y�r���wW�'+�uwZ;��(p(��Q�����L7�2:��9�XY]���Jd.F�����i����c��7�*8�2 �j� �Bv�f���*2o[����Ԇ��R���ҳ�����;�.å�z�ݡ3�\�!m�l-(4�ݍ�>��&1~*���	�'�9㺕6��\ʑ�.�{f�J�t������IxJC�����,�D7.�/f�fϑA_��J�n���׹��A�&v�Nz��!z�.L'�[�Ej��l�p#^ܶ�ٓ�u�� ���@1��
�Τ�a�n+M�@V�إ��&��ѡ���{�#,7xL𐰎�{��|��^���_�BI���Z����K$�&�Hx��Jo����N�L��y�����Z�(E�2�\0I4�Y��ߍ�g��;�/�jRL� ������c? ��M�l��B7�ؔ�%�����=g����)��oq�Q�l,�w�b�-�Ի���|��r�q2��37R�'����t�R�ڧ`r5O"�u׵*���e�!8�|�!*Lt׺y��B& H�A��V�PK�ZY	(�X'I0B��м��8�t$�%�'zCX�1�e�&@��-�n'���O!�r�]�j��R��>�^)[V��}��dXS�&�@�l��f�M�X�T<ǎ#�(&Y�B���{$�D\w��k���$K�t'��wZ��H�~�q2���!~;17l�vͬ�.CƁF?�j���y-"B���X��Z���~���G� -.#�Rb�q�5�g}yr�	�f��|��q�;\n�CD�rO���</Ҏ�i�ќ���x�)�I���
e7���E�hf�Y�4	�{r�ԏ�9�6�^��\���<�������h�G�;��^������n��T�v�Q>��N�q�~4M/R���du�6Z�����[x��Ϭ��B6��q8HSl��a�N��ٴ�J�:�0��S�� ��.��Pc߷����ܭ�OLq2;��P��\f���x���t�nS�g��D��������/l�+<�C�V,A
�G}��'JR<��t�M/s� ~�C1�O�C��,��~�-4�޳5fj�&���qg$����e|�H�Xbێ�Im�:;9�����'��}��zd��y%yK\S<�����e$+EML%L�@>�u�S��4/~���U�d1��X��l���v�%u7��hrK�ct�ND�;�S���.i��/D�u=����?(���M.xJS�Vq0 ��0�r���> s�8H�a�Twt	�b�^0�>N�����Æ6ʹ��+\L%?N�7�̵�#� ��=���Y��B�)�v}�����FMe�0X�S(-dXv��*V5�%4Y��zxX�0Kz�S
w�Tjd!��C;����R�R,��0���Mⴀֲ�=mk����(����*K���w�󵡇>^��ړ�m�,\D:W@��xM+��Y�+8����,����%�w���ϸcAI���@s��{%S��[nZ��F�n:�1�i���'�y�#L���ˑU`�P.��Τ\DOī�|�I�/y@����!^=�M�P}6��Y����k�{�c)Sl)�Bٳh	V4I�P�$�J�W���4�ҡ(�#ZJC��ї5O��d�.�'��pT{�Ǉr����$����@��U�<�R��k�15�d���K ���D��MI��RgT�lL��&�@+�_��?b:H�8w_�V{��{�R4�s�3?��c�ӾA���ͳ�\�P��@$xb+���Zz�{��o�O��%}`�A����AJц�����_��D>�e�Ss)Hh�K�sϾ�y�6�0�_�;��ֿ~Z\�Mtu"���Ky��}7u��$�渗�^s�[� *!�^����-��������F�D�*0��� NKL���v�ŤZ?w�~��Q�}��m쫎�y|Zq�4����t�|�7���������w`��ћn�=��;˳ ��M�g)���q��߅=�Jh(��X�dL����8"�ҽM��c?H�0���c��& �<2��
qbU�\ݎ^EI��>j&����u��@uV����E�ċ';�A|����)���|�F?<��4�𢚩�Va�p�ha��A!��1(!<vU>��d	h�Jn���,�/��ɐn'Š��y
�IBC˳�`��9���?���;#jnbYɽ�*`;[Oe�da6"դ#�Y�x�/�rd�k6(ۢNڦ�'[;�>*��-VT4P��4���K�����Bt�;��4`I��:GtKг�Yx`17\%����-e:O`1u��!�vߊx�_��!䋯�C�'⒯�T�D�9.
!
a���y�p΂B�b��Y	?K���Nl[Au�QF �g3�C��� ���t�#�zd��QQ��V_G�"=������g���=Q|χ��c�wT{Q!
ϰ
��u�]�{�>c�� ���*�Q{��A⢖�ǐ�&&v�HӸ�rFMJ�"MSh5����/���2.i��9��nO����3���
-�I���{����픺�d������#Wz��0 �E�p�HZ2%O���
H�2z\�8� �9��w�@$�4�cuD��C�)���W͋_�p��]��Z⢸��!x�<�u�9���Y[p(�w8�{���������N���B�ڑ?�S���sdnuʫ�N��s�ñ:��_�AݕH@^b_�A�=랇>��	7՚�g�k@p*o*�R&q1�j�?&�O�S<N�Aʌir���
6-�K.��)���58	�2>R~g:�8��{֢W��y�1�����ZMհ��� �T����@��OH��曑),wL@��)�0p9���5�S�f೉g�VT��lA�.x��q�N0�/����W��LA�Ҵ��5	PE��(i��-���i��Y�b���j&�aw7lSG����[̝�`&����v�'�:e��]X����΁ԡ,x^�q��-O��Y��{���סּ��]}��wg��p�K�@�脇 $��÷�uz��z�{����p*`����ƻ�+�J�' 	?٠�8������BؕER� ���M$\]v}b����A))oc��XK��!�@�e�0�ʡ�B�LEc,�������{������6by;���#���Eյ�	7xM�%A$����+:��(
(��6����#���UU�=�U�SD�Q+��q�A�G�9����]�7˸*��gA�")6�̠['��>��0@� |,>$�R4o0�� �/��G� A�R��:��U�����[�1�7��f']�)jN�D�`���x�ty�MZ
CG/�����KJ��W���*?P[i��͓&E��{�6��AG�'w�W��`N؇�3�x�g��:����%��NX��h�a��N��}�p2��P�k�i���M �C���_�0�m����Mh|a����Q��;6*����*�%�)2[+@ ~7�>g���4�;pWI�Zwās�?]Mk2�L�^}y�.�[����n��3E9�g���f_Z�?��V���?����ڗ�,�}R�pݠ�&�T�
�N��F�15ʹ���i-���]S}�g]a��єO��!2[��u����5�$�a-S)��`+��6&ܙ�O� ��z2l��Gqbg*�/[�
�s���nͽ��l���n�twFR�^_��?"1C-�<�V4�4���V��+��eat�]�19���9 :�=���>�0
���ٞ'���7�W���w�6�����m����������J,"����<������3�B�0u�M���D�2%H��|�w�w}ɡ���U=�,6���_�T�t��<��j|�?�^9��><e�=Q'���Mx*�׉4;�"�Qh�b�摚KUQ�`Zs{�&ҫ[
⻩'�|k'
��6�B�M�E�mg�����@G���of�
�k_U\� ë$��%�8u����z#e�P�Q�	�h�\�dIO���`�l���Cx�a^��m~�0$��a�?�^�ŜM�7
�,`�AL���挅�	?z
��.,�.N� ���LUv:�������u'�?�;E���#���xyb�M賽I2ՠ�H�g��V�K����Xp(�=�e��.VB�'���;	m�֍��C̓��5���'�����?��ZR%��Bͷ�`H�S�Rj���1�!N���k�}ւ�c�Z��5+'���䘿S�E���(��i���x$�2hC5����L��Bּ,����԰K�6����?V@<�BuT^3#�oW*vRB_X�B�
����-ީ
w�]��ق
b_�9�䡇�wT��|դ%�Lׄݼ�r��hX�0eq"Z�]�0 Nn��-r}�$C���;r��ŞW�ג>�q�-0�K��F �)��� �|M�F�Ҙc�<���$���r�ÒlO�b�e7x��7|;Ih��h��$(�?�Tg�h�4��z��^`J"\lC��)���4_ �����K�w�M�'��y�E��&`��e���Q��c���t�:��z�@ʊ6�'-.��BfB}��K+)6YH�#��h��g��T�YE���}�&�U�5��yZ��b���E����+�6�1��Et"�TS�B�r ��?�A����?������` (.����!Ta�:���E
]Ԣ���K0-�Gy�@c��A�<0v�2&z;WRf����O��;:���Q�W?����j��f��w��8����V� ܀A��w?��20]>>�$T�Q�5����q�G V�����i?�|+�3
\\~u�)����\lό��o�q��[�Bau;l��}��fgN���ޚo�dU~5i���!���('����k�^-�!|�BIq,�ylHt�}�����&�)�!�&'�Z��U���e'�͕$��%���Ҍ���Z Ly�`W���<Ͼ᷾�3�%�M��x��d0���~���&���4^��a����Z��30�1hy�B���'�wy���H8zz��l�U������c�_Jm��3.Y�"2]���
qw(��/���U�.H� �j�̃|cu:r}(��^�=�g���}��u�Ȕ�@4֣�+��.�V����r��Jrf&��$���������-}��kQ�(8��W��#U[�ؾ�V^��3��x�Z.v��$�pP�t�:���	#��g�}UnU%�R)hI��<�d�����T?%�$t�x��9ٷ�=����M���SA�1�JL#�y�:(�xoi�@D �6�(P�[>��$��iFI�j@L`�-����"�&L��jU��?�&�7�������aq�Ku�t�6��N����Z�)���G<�H��0FS';���!����Tt��33��H�ر�X*���7sӋD[��N�n�t-.�i<���0��2�~�mΥg(U�J����X,�<����zc��Ai΂��m�F�T �6�a���xǾ�I�si +��P�K��zr�r�.�|cH�A��:�K:�*�ŠU���p%�ܫ%B&@;H@j�b?�&�n�{,����U�Kr
���1�)%�/�qUe++�5�A��v~��R'��@Ef��B(���4ZXj[����)��Q�����u/*}�W�r5�s&|c˙w�*�p-�.�3��(^��>02�Ҵ#>9L�8*	�m�)��[N���P�����G��ɸ�h��_W9�}�	�BV���qr�q[D�������0)�w�k�q_5���]c�J�6\d�s�c�Y�����t���B����W}}
�3��h�g�5��D쌿�����럔�'L���"��	+^�����Ȱ���b�$�*�%M�2�y�51*=	fI)�����P�S��f>��<.)_8�����M�:��7˫���i" �܆T�"�؎9�ك�{BB*�N����aoSj�(��V6w�nͫɘ�GXhw�&5�В�� Ig�U^��u(80��7�)"�#���v7�����N�2�A�b~�C�rf���h�X��`��-�!��!W�D#�
��o�jh�I~���m,fLO��8eM�v/$�1tI���p=�r��I-AĚXn��*`�=$���_�D��+몡{봙Q0���s�I3�-�y�sg�fV2B�_��g����I�matU�уRz�,�����h[��i�=_7Q��oZ�ȕ37G/���5�>�a�Q�
���F�	={�"+�Ƽ&V��ڠ�3�w��U�YXvi1�h��Sފ�~�$/ޤP��d���sAv�x�������j�b�tpiM@��E��"�z&�������!9GFG��ϫ�w��@���w��s>� m�h­���SƯ�z���n'`�.�H��m��/�&z4�:
�vr�l2>E����-gx@��EP��/'�H�緯��x�O�������?#�"�}�T��HL���X�\5cX�1�me[�:��4R�����+=[W�/1=#oD��/{B� 5�ɍ2������Vs�h�3��@�o��!k�)�)��B��G��1X��FS~nt�ؐP8��pJ���\~�k�X�c{B�WD_���WJLPֹ:݇_&�k���7]��5�a���7�e����+�z�C'�>Zh+��L�.2�t�(� ���G�����5��c�a�����u�|�A�UD���K���^XU9?о��)�:�u�6�� ���x��0өX���E��)?9�5�Ƃ��A��-S~��(����E���hT�>jJ��Ԭ�7O�!yի������X�"Q�2ՠ�fPb�`�h�"n�Dy�d;��h����~�
mkJY{e���;u]2�m����KVB�}��pq����>�"Nh�r�!�?i/ �a�Y9P=���N\��J��I�]���x(��~$���cz*[�u̫� ��y�}n0�~=~=�8���e����ԛ,�4%��>���Lb?MaI���3i��S��bLG��'锈t ���Shy a$�Ɠ�J_9���0-����d����F{�K[�������+��a֓�$�|���SR|3V�K37e�L��u8w�X��(h���xcbN6`Wpl���$�-�@�v {��K���k/ZXD�.W@�Q)l�>@�0��4�4�q�!��w�3��P����-2cj�R���Ni�9B��l��sm��q(�� �8.a$B�����X6��q�'���7�x%w4�y��H� s�QF�5#g�$n��o���3���9䵙G��-�ز]�6:���m?�H�@�bR�kĥ�mSĒ��SX�AJ�"�X�l3�_L{p-�i{��NZ���=��٭�(~
B��;'}yZ�%��Р�z����H~�b	Tvy�,ی94̗3�o�b[I��E>;�\���L����e|3�K�y��K�˧��х��(��W�]#��_܈�>;%�����{^��5�+�[$����ЉB:<~.��Z�ulML�D�.߽U�^���D<�0{G�pC
��K^,7��l*ۉޗ�ĩ�����Gu}�m(�w���{x��a�fP�׌IG���V?{>cdT�V���S ��ȇk�ǲO�߇R4/�R�Y[9,�|l���	,r�1�B<L��
eդf�Q(�*��ԳJ���;t��H�';c,���	ʰr`���m��c����.�>��!��X�v�-�#`���e�x�'N�lS�ۤ�f���xH�ɾ����l��ۏ����h0%�J�M(�Tw��p ��Z��%J�&۴W����e�<���q�H���4�!si����X`3��$�s��/ڥ��,9]�T�S�ի!q ��Ӧ�+���Ne]���|~�₽͉G�����R	�l�*�[Q`g��@��C`�Ƌ6Mû��hQt�ڈ�����t"����)ѷ��W��X�Ŧ�`��桑�`s+����SY�:�Ca�	�w�Z�yr�c]�(ApױNߵy^�� ���T[@�O����B�^�Z�%_�ڻ[?:]�p���
�H�-�&N��'M��D�8I�W(�Jޥ���PUtᑁ)�]���O�����<����eY��s�@�>����J���ч�4�R��������āSW
o'�@!SD��W*���J�g��y��4]�EP�*:ȅ�>��C3��]��J�:������z����C*��n/������!�� ��H�z�z��t!�ŋ�YSսxN{T�2�/��S�G�m*�)G~����洏�4p�oe�jb�1Zyu����*[�#����t�mܽͻ� �Kk�X{JX�o%>�wOھ���DEtz0����X�I�\]_�VZ�)a�)|t^��<v�*�B���I�ע�ݫ���+v�@I�y�"���C�2�x������cxmq.��ld�CE�E��0��N���g�[�z;�s��*Z!?�sVٸi�~��)_z#Q�t̤�R�:�_���q�U�!:��z�\���|��] �h�p�����r���{�+Se߷E6z�{S4���d������$���j��/�z�2)t�>[�벌]�����"߷EM�ϖ�I�f��FC�+VJa8�W�u	�$@�E�1TQſZK]q7^�A��ޓ�V3 B����|bD۰�}ۈ֚���d����7N�e�Y97��Y��(�Y��)M�X�d��*���ޓ4SK��;W��5)
�i�t��<��4�޿8�
����cG.~�Q/#y�@zT�a���8���+(@����	x�����B�j�����EqY�7�پ0�a�,`��_�q �9�N�V>�f���B�&�+G\q��Whɰ[�P��/OE#��t�s]BWA#�qy�0"*����$����fbZ&�wa������F6�1��ih[юٚAY��7Up��nn�p?_��g`�=���O}n�X���-��ڀ�^ ���К�>R�	&����X�Od�!��9Z�����.��;��<f<�@�(#Փ��TJr�EB��U=�/���|�¹`��n�L��Ɲ��vf= Z'���"��������'X��̲�g.m�#P�&��fpPD���D�ό+�w@\���h��udA=NYr�x�%��74�(�[��49�M��_Z���F��C# R��{
�N{S'�8�Ա �%��Ƕ�ww� |�S>�h�S�R0��L�dѯ`�	�s5H|m��?c$JCՃ���GH�]B!�Kp�G+63�X`G�ͯ�6���g2Z����@Bhy�J���i�tc8l���S���[�.7�_�l��|�B�@ ��v�}FRP^�d@L�0�ɑE�@�f���:��D�.º���i]��	��w7_ւ��y�����Q�d4�I�
D��pq�o;0��գ��,z�ʌ��6�F�;�S�Z�G��Rh�Ҵ�g�_�]��S���sYP���X�g���3�!���lU�o�e.؜���tEhچg@��+���S������e�T��i�cjB�{F��^[Y*?�Ej]���rï8���g�5R�p���*�@�7�,�}��CD\j���t��j���r���u���5��(�]ߎ�lGO�l��:�J�3�hK{M���nw.�5����J���Q�����J6��9FX�I��;g2��O�l�y6K`�C����;+΍�����>db��8Z����!�G�K^\���ö�f�S��3�%��im�=D��g嶲?�i��՗A�|ŋ�竌������P�K�ˮV�Zp��͛R�e�JU�{��'�	�U���?R˟��W{_h�vU��d�(�#���5�F���KCゥHc����7��0�b��u�֙GKt���47ʶ��6%�_�e|ߊ���@���u"+kz��0<H6t�6�t��a������`�[�_���ˏ�	����Y���R������]��ݦV�Y����i��5YS�G�H�9�@"����c���Qv�m_Tb�[�ټ�����<�͝���@P�7_:o�ȿ[�\k�)([�pM[3>Z_�#!6c����݉Q�
�0�r��mHWm
;C��v��������<�;���xw�[��*т[����5H���R&'����;繸p�W����͟p�ƀ��8X�&���bu#�d��}G�lĎV( V,l|��U��&��)I��V��q䘌]i��T� ���B��R}��]��<e������Ʉ�xl��՚"�+K��=�(w�pW���%rv�T�\T,��(FK[�V�cכBa�����y�����������֫�^�\�eP3%�(�]���׷)�O�X�d�0�_7�d���Y�WO��Ĺw ��2o�������K ��;aU��41���4�
��=[(���(�_n�u-��f����>��n����ݔ!ZЈI��|{<IN�v�S����nB��6�*s�sY�AcX&�bw�
C����Mgڷ7���7&��KR4�!h�D�����E���>�aY$=�zu�QM�|�#˫�ou�� P#*7�����j�Pvڟ6���G�[�GMz$%c��)�Z�}ޜ�	k�%Ʉ��B��y_^:U���	�����ݱ�=��d��Px�<mq�"�	W���2ЎN����¾fK����٧x���鉘�ɸ�;
�M�9-�<"Mwf>��}�4΅̳w,j⾙�:���-2�Cq@@���R�f���ho<��ò���t���{<tw�_EO�0������d6��~&�3o���8Y~�<�㒕2�0�,ݘ�c�C�ZiAk���'`�ٿu�Á�l��;Lj��Z��;�C�3<�������躛F? .kă����k��>Ie��������p8�܈QB�f��F~��d��e�M����tT��;3���81�E�.j�X'3�p�
��C҉�.���_��>j��1Z��kՉ�Cf�=ЎCD�M��@���l���+�#E�l�Ά���R��삝,�y�[;;���~�\��J�W������ �r���nI�&N��,��=t�d{�y(Q����%���zӭ��Wތ!��(X
�v(����֠����א ��q?mY�i�ģ�-��Tt��]�"���r�cf��JB�9A-��H)��x�I,�AL\|ҐZ��="t ����Oɝ  ��Ѓ ��u��Kh.�c8�]Wf̣�>R'0$�1+�+�W���XiҘ���]����o�-�b�Z�A���|N��я��o#י�o��:���);����i��T���8���|�Cfу1����j����:wnciƢn��s���k�7a���R�a�X��撅�#.�M6�iP��!��L��u�X�dN�ufHT�X����D�6�V>k�`;��&�[�d��*���AM3��f�R����VD�u����C^}z������s�TI��?fS�ǀۙ~>��a�I=�9V���bP��]�u��1o��ҟ_���B�4��>�/�׵��K�-	���v����G��-�>���@R�{�HA��<���Q��V���8p���y��|��B�5�S�$��w�9G(c�+��B�� Q��M�[ȩiܠ�%���}4�LT�~��U�ݣJ.���{b��-o���S������B@�S�ط.ʡ��Ĝٔ\�.�*�Ў����KV��͛�����N}�ͣ�����6u
����Xo��,�(��}ؒv���W�_���Ե�~QL4�	�D%D�D�g2IL�Q`{/��B�p�m*��u��&La�Z d��yq�:��yjBu`��{�R̺��g>� n
ߓ�����͔�-�E����/&��s�k�E��Ρ��sr �'U�Q+toA�����^	��Axs�z}�Vf�~���_��f[5Ͳev��H����ո[I	�d�3��gћ��$Z�Q�K��--�뗑�ɖ����dB)Q���d��*���.��1ᐔ���_�>����K�)yp ��.���l��_+��g�гh���[S ��QRm�w4�ʭ�xӽ%ƽR�y�nFh�)�&��0X ���W���^qd�H0$�cTQ��;��Z��asfɼܣ���Y���2ĸ�6rK���6�W���2u��7���'�)!s�y䰆��}��у2��:|N�P�a�ˍˈ���=/S�q�F�/k��.L]�D]�V�
�g�E4�L_K�e�i�؁�{Mꢕ�ɦЄ�o�_w���'ώ��i����V���HG�x�n�:�6�> �Q��&_���Ip/���Z(�g��O�O����K��I����PQf�`��8���ka�`Ң� TA��~@5կ�D>��C4+��J��:ě*@m6����M��f���V�:t��.T؜Xe
�U4���4�T���N��?m�0,?�zۿ}�^ ))���h6�E�,�����>�^��g�C^��o���Uf�ۥ���W���l�7�Ep���~w=k��z7\O�K�ҋQ�td�� ���k:;�Ki��M~�>s���"�A�r���l,W+�ad� J	����`��Y�V�?�e�T�ͥ��#�~ݽ1��Ѐq6�	�y��\���K��W9Ǩ1����~�#�:X�������Լ��0v�R��#yÐڑ�	���˹���d��n��?h��Il���Z��ǛV?q*�4ve�ϢG��#ra-&��9�y�}8�����)Yp�Mg��>�H����{�-^VB���>��V�A�N���"*�$���ڮ�5V�du��L�P[NL� ��Mk���St��S�D~����\{�<�9�4y�8�'�B�,\O�M�G��rKS4� ?�G'�IƩ��hu�Xթ7=R��([p��6Lz_�#�ް� 5�]ZBx`��5�H�H���2"�@����&�I��y[�|�m�A1e$c�@K���͜KۇN=��{�
��?�E��6w��&c=��S�V�W�
~�l�J~���V��T��a'�Lʉ%Kʡ�}Mܚ"�Q�Z1�b�f%�mU�0���7�z[��˚`ʦ�(q�x���A�q��n<� � �Y�y�[�+q����b��P؜$��Z�2Ea'�x=���"�3و2�H:�����%LbӸ��Aa)j]����z�q�^����ג�#]�� 9�'��2O��uf�dYc?E�R�����u����7#s 
d��tG)ѓ�{��A*�if����u�����o�V���e��p]X ��O�<��3�/�N�S}޺���Z�����w˼�o��>�zV�]x���O���0WB�*���K�}jB�u4{>�wI\O�
�/4���!'��q� _��H����~ow!/�9J������1��v�\��j^a�y@4��]�0]hjN�"�p�f�XM������V��[��x7�(W�Qx[��N?>|T��b���蚚_GHp�����ݍ�` ,ζ��	z����U�@m4~J�(��d��E�[Dj��1،���J7�Z�ō[��pp�R���]dֶ3�a�����{ʓ3p�o��w���*a��'ց��r^H�>�47ʧ���d�{;Cn�D�;��� ���M�h���_�����>6f(�AM����D���Z@���b,��ҹ%�+'���9�7YRЄ�2,�h�G�S%��j�E=�P]B��G j�+i�M��^ ��}U/�8��(�yb�Sk4�� ��엜;�P,1u�}���ae"��.�u����/6?*��l���� Ѥθ�����7F�z�k��3F������#5	�V�	�J�K�x����-�wPO}C����g$�v��?�֣���қ�v(�i��s<�j��P!�M�#��X�xG|�C���VxR�Ę>��O���اKp{�[EY�Շ���ѿ��U�R��{Cĸ�LQ��i����్hR�Qa#�U*�j��k�T9�a�屄�R�Z#�qH��4����E��5_-����^�;&r�vQ}��?o_��o��m����9���v!�$�ۯ��]]��3+��j��{T�k4�L������2��ݞPyg����)P����	f��v|ҴX����3d'����F`(�Til9jy�3�_x^�5�	$��d
k6R�7�{�kOϧ
���=ɧ��D+NrH[U�	�Z=��r�P����,!����賬������G㔈��=^�R-}�cV���?��yk*�F2W�Qās[�	x��'�.�2�I�ʌU��Vʆ,6q6kk
���|"�2��{))���i=��X�x�o��P:b�:��l����$r���LeԆ)�p���0(��^x�J��W��+�]LrXk,��ڠ?��Ypa�6�S����E�$�;[�.���L]���i 1O���ǚ���T���+�%��B4��}��e�U�6����2�1��+�T`� my����}Ofa3�Q��t���Y�78�3�����l4�p+��]&�!��WY��둋���F
{8��X`F]@0��{�������S��3Ț��f�Q��i_CP'Z� \�4��h{o:��T���6��LD OJ��z] ����K����Y����UddH_�J��V2�n�c!���SWR�Y�8Z�i�u !�?�D�tD3r�OGI�Xd�=�|�h#i��J�-C�ʼM�p�)E����p�OV�a����uw��-�T/.�_�4�����y'Ll�\xkG�vC}6�P�mw/q8�My㵖m�}=z]��Y�_Rh]��^��C�==I��C�0�#Z�w���n�"%0���<q��M�«�gmw��"?}^��ۢ���Qt��D'�-�����d#���lǞ�KI�1��/{[�lr�1���W1~+c��S���ŠR�������A!]���c����n��\����c~L�3 �P<T���망��۷�Vu������U�
K+�,�VY�v�ă0�������Y��zSQ��|�ԡ^�rHJ��=�O���I��r��9=W���	��i�V�چ4ۮ��R�e��u7�A��v;�)6Ÿ��;Z������[&4τ�@8����EY�������i͓XD��6#�����>���|�U�q�NeY&dneHh�ɘv�#+{��U�=�(J& 6o�҈���ޙP&��%�|*���8JV���'@������Z�cX��-�%"^B
 �uǓ\�DlP�.��Qqj�hL��Cdg���"����`�۶�_?l��߼(�7�K�r_����No�ԏ�l�Q�~eg��}�A��;;�aa��� ��i�]��wu�!}Pt1k��v����g�g�П�,��5��41�ω�v߼��K�L@��(�e�ӓtL4�e�1ڷ�
��г,�3�>b�3��E��[�������9�=����8J:�)cf�_y�oݗΪ�0z���O��7��w��ׂ�s��u���k�`ฅb�\}�d��A]��Z���V��q�'4t��s����Ӕ����aMЮ��re�>f���'n��E��;��Kp^��M��3��G�П+�_����a�
G]��BTyl�����9�Y9�hх3�	���ξ�l�H�5�s��1�	r�3z�8ʑ���׍�����e�`����һa��1�&'�C��ӛ*�c��o�Hz���E���~���
:i��ȯ���ۚ�Y���qw�f�R��jW=U��[]�d?
�,f����yZ�$�՘��/�$���g��il��Kƥ�1��T��	\��	�u��3#�M:b�@P�4������?�l�Y�����s�}�?�dM�*��N�[kEs���hz ������w�ߗ� �]�}�0+�P�*��9Α��{��"�p��	����_��Հ��se�O/]���  �(:�ں?*zG�PR��/'\�з�#���tc��GO����wv�����۽S����|��G���H�[�Y&����[����b�pk�OJ����@jr�ȴ!��3$�b\����RR�U��]S�`���̊�$ʏc���V��>P��]˄�<� ���1lm��f����bz�/N�
R̛��&�36c4�˧��fn�VqֿY.�d�9J~'/����]��/0���.<�ҢX���Br�/���Ygǀ���A��|GAb�B�Z��:Kp���.
.w�Hu�P��)?��eW��s�c�����v��ui��
��13Pa{`�[^�!::�>�����gD���._*��E�Gc��1���.2୯�Y��
�� �,։�y�0%�1%��0H h&^�"�7�Lϲ+5�K��O;�Y������p����lk,ZQ��d�æwamm�,��RW D�h�\9hV�ߑ|o�7cۙ�3@ N���G-U�.�;�&O�,��?���]����]�e~p"@���� ;���83w�:���t+��:�,i/��cۧ<�-�N5�B��eސ���T����TGܤƮp��ʅ���RVCWLϒ܂\�hI�����W�=ǧ�%��;�byj�/�=mY���	�9�|�4'(��*�*���a���:O,���0'�f�i7�Ƚ���e(p`�p�/usbp�z)E���#T�I��"�(;��O:ڭ�vʟ�fr�g!L����;*qjL~x��?�[T��{�ܯ@$�k�Z���߆�~l�D�յϭ���y�v�k�2#��7�s��{����i����u�oss7��K(;dm��l�8��j������H�t�Ð'h�_��ۉ|�>xYT@B�6�8QE��{�����A���zN�n�r�p^�$��pzy#��A�(�l���㣭�_� ���&?�7�X���,T���J�xy=�n��V��>w�#���ً(ݢ;�/k:��k5 a�#��t��zA��C�4{s� W���U9{��������$<�>G3wCzr����szb.EHŇ�(6ޞ0�b��[cr������c�n�bi�ff8[+i �0s`�ߌI�;���l䦛��ډ|�5wy6�e����D��y�?L����B$��UA�i~��1Ao9J��cw3�v�M5Ɓ^+@��v��α�A�c� �{�s����WJ㉿�K�(�_n)G܅�MqpUI�CM�Q�RQT�R9�Ǒ͎n*��..��΅G�v�ۉ�! �(���,�KH��.3C�z:9�FQ�rRp/6. ����N�d���X���0�]��	�K�U���M�5�������6��(a��nՓ�xș��b��#��D�v��̀k�/7��6�/�i%0�jx�b�x�$t�<�G�;ZE�D[9 +_�i{���h���HL4�mB���~�+_�|�C5��=�pbvj�䟬R,R���%L�,��a��B�Y��$���-9�4�|M"B+��r	�s��������h�wPIp���L{q��P���|�J�]��D#��h�74��+�ߊ���S����.b����A����r	'�ь�=�L$�2N�2O�Q��щV�/P�N�:�J2���"Zk��!�9R�o�o8SZ��p�FE�K��^]��"p��P@�����~ S�jYA!K/�����e�-||���l�D?��a��أ��)u��#�J��m�@(t���X#�Q����, *K�LO���Um�r`��{~�$/�T便�xA]�C��	�:t���$�;"g�&�'o��A1��SJ�Bce�U���,��N;�Qb���ZŚ�[�S�vd�Q�90�
��>-����6^l�ګBc�Ķ�9�ۂ؛������j��,��A�R�rF���g<i��Xܒ�X�{��^�G@	t��&��5aOa#����yݎ�H6ƿۀ���R}�ݠТG}���N�hW������Jه���,$~��	�ܠ�@)&�4&F�)k���}��O#eT�_ L���L`��%<Ԓ� �6����;��1:��[Q1��H���rN٬.1� �e
�)x���V�u�$�	�A����ݲ�Þ�9�Y�E�FF���`�e�E�c��˪s��L(�4�/١�́/���#��f����C+��:��-r�sܵQ(����p�G&	������<�4�羚0���-S~!��N/Z��c���%�ҁ��*�S������8T��t]��؅�pߟ�O?�N=*&6�}$t���t_=Ͷ��X�A�1�!�~��t��_��=��4E���pcQJ�%�w�PEW-%����a��p\�2��^��K�<�yn�+Z�����q�GnƧ���U���%��<��04�m%R�Lǻ�W�\�`>=�o-����-�$� �'����%L�ؔ��d�1i������_�y������� ���J��!�N���������a�����A8��"�.Shڀ�?�>�ǬZuݟ����!¢���	tP�4/�3���c���LE��$�:W��̿�"Hq�#0h,]ק
y\
�/�,z]�4g�wq>Է��°\^�z���*���	�� qmo� �;;_誶�|DWQ�v��'�}L��d��Ů�.�왊S�x���������f����"�x�RM��^��PCTc�:~�ť������&�p�vL�a=$�~���k]xY���u�G����n�̩S4��~ҲK|�]�)���E���%��$K��s�7�u�;�ȿ��d�z*|5��[�Sҏ��
��<e��M�D \�P���:ha����BZ�%��Fw�Aq4�J�}3_/�覠4c���v�_ej;��c�,���t�.�GM^��$�>I�C�k�2�k\R�H��Z�����%i��|�.�47
����;O�`�u��(UF_�\=<a_!���Q��Ɵ��ˎ�٬�A��5��}r1����z>�+����Fl�����7b��a�P.��ڜސ`�Yi1�%����O"�j�F��h�<��ڂ<�~�?a�2���,*�w��&���Q�j,��m��ѩirn���3����?ތ��LR;��0�q���t���R��qm�f0ֻ����P�%t�s��.R���LL�S�x�;�-���?c��k�;#N���,mU�Jƈc��V��Q�S��Oܩ�K���2����ɖg�[Gا�&��$�OV���o���w�eE��4'&��b�)�;״gyK�/����T��W�����V��&2���:���kr��C*�J����t��{5���ڧJ{\���+�����ٳ���Mtt��8">_NF�g�ք���A<�u3��Q��d���Wn�GB��=�j������>r��n��"���>>tC�������hY��@���ےD�)l�"���C�5ﺸ�K_]��G�ݬ�:X�rؑͷF#�ԑP�?j_N?͜)�B�;94<A������9���a�%hs�R���kyުr����tPˮ��2�W���?� �j:q%��l�\�I�����C���:�K�����
�Y��(Ɖ�$�1�{SnN>�ZA#T�i��0W|��m��r��R;���)jj}����@�q��R���*B#��=t�����i�����WGMZ����P!c�K����σ�V4���P���)����O��9}58QN
�<6��0Z)G/b�I��z�LEMýW&�i�E� \#~����.a*Gj���@��DĶ36���⍳�R�[���C��~���;\�
��s:��|������B	����\4�<	���o�5�Xg�+�� M'��ʘ��@����-8F�P0=�{N.����n��KjN���L�&���M��͡�e䅝�dt푃�Ψl�=��?�?7)eĠK����hb��k)�����&-h#T	���ߠs�-Ed�!tb~��w��n�������r������ca0���#e	u�� ڸ?��p���A��7"�ݲm�R�X-���J��2	�]�Gvx�b��E�䐏>������N��fST�҆;�l]��S�v
*EOWOB���cx�g.DahuX���n�^�Gh�&��G2Z+���>�Q��#��>/��]�Rҿ����n-�r�1���c�uNy�V��S��֑|DQ�u�:�k��R�ݎ�J�9�P�)�Z��#X�8�T�!	�B��3 �.�`�+�c:ɖ�Ka�x3�IUnL�q�v{dX�N{h�W���S�gz�k�������#����=���NE�J�a!������O����B�	ؿdx(y��ȹ���F���������R,�"��mz�ܟ#K�P�_����%s�d�$⦛����r(�؁�["�o�v�k�/ ��.o�������k�6(Qwޣ������얱{J�-B�K�.(�$�X��-���\3�]kd�����m�*���l^��1��FCP��dB*��e^��pܨHݨ��.�T�}ο�Ѿ�"�Ƃt��+�ޟκ!a����5�����e��-�0�f9���z>n��7�U�2$_�\���9"*���"B�U9���IXW�V���O6�;Lϒ]��]P�RH�Af�y���QA��,��C��)��y��! ��eІf�g���U��V�RkV�/�yE�R�3~�I�O�
3�?� �� �#���&��Gn(�	�+J�,�m�G������$�uΛ�24wC������r�ԯ�c-����u�	ɞ��GnyLh	M$T܇�|�u�3�Ue��;�% ɲ�P� %	JO`�J�p�ʺs�������chw63�R��k)c�Z��/�dҰ)�Qv,��vUMn~X�5�^�/�}S�&��:�Qғ���G���]��Z���i؁{Ao�B�Z��,¨\�"4���J"���P�6� ��Y,|��L��rR5��&K;+�O����!�bj:��"�T�l.���V\��}Κ`�g�,E�ȴ�ae%�v� ���G#3u���k��5��}�CY����I�.����Oq�Xc�k|ʡ��yC�v�l��ģǥ�\Oʼo��e�#��O�x�a�>��+���/i����D��q�B�-��n/���� ��E��y��h�ʵ�{�#�܏�ʩ(!��d$�l�q���5 ��=�ս#%�5^~���C{�@������" {�II�`s�[J���v�1�u�&�[W���(2B��=��X�����qx,b�:׌����m������!xk�����RǶ��X�^�&=�F�d�C޺�R:j��H3BMS��\��a�{Z�?h[�SG�W������s(�=��L�5q�j�,� T�jZA�Ê����~�N�-�
zR�yk)�.	A�+����?��LJj�H��h�����:�n�0G	r=o&]�[9��]�p�8`^�2k���z�=����Y�zA�|��v@�� =���V<�[E׈�B�s �y���p��T@��,8�am��"{�5c��{��3���AGԆ�E�����Ds_q�
��JB�T�u�Z���(�[G�L7^�>�A�b~��01�8�܏^Z#r{����
D�߆�U �Mݐf:�^��\V},�L#����c^��c�G�rN�γ����s<:�U�:b����y��o�Ԇ,�=��d������k]qe2�"�g�U�= 1X���r'0 ~֤ƦlNyK��E�t��r|}�ʸ�խ�a �Ʈv4Wߦ�;�Z�s��y�t�CE^��W�����;Ǫ�MK��xT�R�z��ڒ�i�糀��1�
�I��^U߸��#V� �]�E����$�e|"8eSi��+T��1^�E���{/_3b�De� �р�cC�f&����gR�,_hz��m ~�6�pЩѽvC/"�/ȭ�.4�)�av�bH(�g�̵!TX[iw���+ e����֊>��L�16�;�#�V½�"O�iL�%~ۉ)*AH�x��M.&�=:��������6�%�3xS�J�h9&Mb-��U��A�W$�^<����1p?N�s����C���Q�eX
�_o�
^�Z �#�?^�/L�����sN�Y�t2=~������}Q��ƠXq���y�a]9�+A��ň��,Y�ΐٱ�5����7=,�3_��ߩ���\�bK�����٩��u�\Qi��M1�j;�Y����<���J��R5g1���js��4�g/qg+0��	� �z�M��2��˺8Y�ˡvE��,������ߺ|�X����K��ʫ�xI� 婽 e��q։U�c����~�gQ�c��%0� 	�ew3�98�X�z�PD��}M�%nj:Y�GD���/�FP�Y2��� QL>I��ye��u�����6��f��?Y6TouV��*?�C��A=|��}�������s�7����M��g������~��ܔ?��c�_Z�]��V�&\��0xߠd%��!���[&����
�d`��>�%d����c�k��>�f.��m �C��:/5�l�vd��nʨ k8�lk�k�U���h���.���Wi3�+n�w���)�Sd��T�Н��;�tH��z�"���bZ��ނuw��n���<K���Y�ͬ�[3{s��w;w6Sߚ��8�={%��S�sK��&��3�˺$_|�_h܇`b��+��ͿW9�\�2=e�o���Ú}7�$˦�T��I�6����e~��2 m7��u���V:��RY;T��*���P����4M8��e�d�-=������~)tLJ����֛�s���!�C`g�yJe��u����^�c�6ݿ�ս���u5=Y��Tk�@b&+z�����ӷ��|�%�S����s�]	��P��p�ܐGZ����M��I%����^_����ӄ~2rF%�� (�m{�iH�X=cA�z�؏�ʆ��JB�@�}���H�ӥV$����⠙���Џ���l�n�L�����#io��ft��h�5�r'�h��Oi�\��r) EXԂ����5wZ�K������sA��^>:������:~���0���6�x��"���"��>����Z���������
�a*� v�Ӳ�t�o��CP԰��qNi�y��q��N�3�\���6]"�Z���p��{6L��L���
ш������{����䬖44�Q�Z�G��Vhm��|�a���C����z��T����Vz���UX�B� !nN~.[d��^̚u�#H�I���T���It65�>�{�_?I�ƿ�Nb2S��ew�rPƑ����y���W(�0���=�}��I�B�Z��-�6 y�������^�O%trAh�N��bg�O0��>얎^�U�`��A�0�e0��!��l�J�u錮�g�84�bTu�5�f�Fd�pZ;��2i�Y�7}�=j��*��k�$�?��<�:��u�˼3��d.�F��*�����]ۀԴ���H�A��s�]�H!	�(�4z�����%�1͠�5�7ƃ���y	��O�{��oՓ��vy�w�4��Ŀc�:�A�r .����%U2:�-�GMVz��ʃ�8����YAʅ�Ԉ��+�0���@݆r�\'u���N�O'4���BFu� �� �����p�(<��n�۰�?�S��)�Ӹ'�d���@��/�ߣs�?L��	�CC4CpU�艱i�B��"���QUz5�f�m �OM���"B�aA��}� 4���3�>�F/8W��@�v#5�ӛ7��.	�D��{�-^#��V�ۙ�t^�2��S&��*�����E=��?��V�ff�~�e�]�D��D9o�'�ϪϨ�z��eUpG��f��-�h7]nQ�hl�i����:/��,��l�w����_��E���A�}_2��wm��bL A��=3�����Xˊg7��5�ed@�����U�JV��e#��ct��\��߇���������8j�x�:�MR�,���|���F��{F֋�uE�L��7=|�pq�N49��P��[XwgeFx�^="�Q֗��?�TL���%\�����������|�L]T�%��SM���nz�@�"�|F�9 }%s}�B�+�23_{i�3c�YU3�̀���Vl�:�����x�"R>s���wV��Ue�-\㾸]z�4Ǵ8��w�u�qh	57#QC�D��N,4�l\��{O��/Qrr��T:�!C�~�� ^�PR�ӌ%xTb_�b�j�Z[�qϙ5�Ņը��V��=F��[���(3�.�2�_C8F�/��F
#�8%��R�#�^F�*��n9����}+�A�pa��E�|���3�aU�D���s< �}���B��+
��,}ѧr�j]�H궱��RsR�#l�O�����n��~�5��X�e^\���_o���|�M�]>6C��z�|:I)"~�� �]��˯�?�c���MӐW�aY��lf�a@��En�}���&��3�rA d���F�Ψ�6��� lC@R�q����K�%; ��"���aK5���|�a���K";0��$j����	���㣯[;���s=6�p��j4