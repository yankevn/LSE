��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۧwѸB�;Q�)�q�ǥ̥N�y�7x�S���1+��Aҏk�A�hg�S����	�㳰SC�����Ylj�;��Ɉ/yl�Xь�}G�X؊����;�'��VG^:0�y��F�	���D�:j�k̷��u��F'U��X��ù-�h��b`f����#0.� ���]!���豉��Q�HԞ�8of�D5!m��%am����Q�ݹ�u<��l!��@}2"�_�y�k�dì�}.3�槱�t4����$ǌ�4M7���a~�k���";d,�>߿ufj%qC�͐d%�̴�R[U]�s,��_����ȱ��`:�C��4�;��ё���5�щV�/�u�uvC��f抴��u�	_�߃G 宠+r�M��plֱe�A�v���`�˥I[��d��65���;`((��4�/dC�$	*�Fa	ֲH�ƦLea���]j����Ub����(���N��� =�p�s�<ƌ�;�n����n4�S1Pڱq�j�H�6���b���ٜz�����>8(]oQ�v��ϟ����4Μ��$�̑� nK�m��ɒ������	�j!x�L�}�����SL�����ѕ��Nc��K���!�꘣�~hyr����O��'�R����d��o�:�s_�/�\����KhxX�(3��+gެ��R|�r�Ǩ��z&e��� �b���*�YM����dM�,E�P���d1�$��������Zqg=���,���[L�3�Ii�}��m�����<���VAn&,�Q���t_9ߟ&x�C)!���{bn�|�9��7�-�E�i?`��q�R"���W1;�}5���Kj�1�I5SP���I��r��"*y������Jmq	��wS��")�ro(�`�P�"��!d���MBj�wlPa�M�qE hv�H&�<�o���aK��T�_���~����S��h�X�>���.�0�����L� 5�������:��&z�RƋ�T�ʆ��bdt�s@Т�� g���� Ǵ�b%�_ۙ[b�;	iU
����vZ�4��x���e�S�}J$�C�t����<������N�-�1�|ay M�R��+�"�Q}!~�� V�gA���|�3[���?e�\c5Ƥ߱�	���
� 0��*ˇ�B�!����\� +�}Y?�8��AM���"N��{uVBc	c&���4��Pa7+W�LW�%���"p2��a[�b�{�RW��Ĝ�^�m��qD��=���;Z&\P�.�D}�%q���z�&�n���ГG,��Yؒ�;�a`�$=�sZ5��npė���A/*��଀rj}�R[
�|�R��G�y�A]�J��S�6_���N"�I�>^���҄�J�I|��8O�,Ξ�C<��j��0]�h:VB'VW�i<�X1Z�ϛc�^W͹N!�Y�Lv`Qц�cس+y">�����ܯ�*�|��I�T�ͻw_����ἶ�1.�vEt����|���k'��`���~B&e~	N1S�Z�=�lܠ`�����L���?�(�w%m�G��*�C���#`��
�`Ư*�G�VXoy��OTj�wt�LX/�q�����h拹�?�f��@Et�:��?������W\S��$l:΋��Û��A���	$�^@��CHj*��t]Qe�
3]��: H4v��84L\�O'��'�I0Q)�����LƢ�z��Sm�*V���H6aR�[i��eˑg˖gJ�_����7�|�ROFz,cC+i_5�L��{��Ė-r� ��1�q��2~Λ�l!k�s�n_m��<���G��0꓃H�f�޻���U�P�d�C�����A.�b���Ғ�F�*���6�q����^Z\�u�b��l85bz,G�yBb��dk�O��yx��P�wu�*n"�����G����� (	0g7R�~,O��������.��Ap��%�3���R��]���԰���I�ԕE�tbl4D�j(��?�#��qfuҟj�E.ʣO����������z�[֧��nh�@�36�8Ύ0`2���焬2l%n~��>J-s����\�EӮ�&v|x�n[��:�(���@C~K�$Z����"�����e�(i�Aj���,��TqG�h
n5�:�Q��`�]C�{i�;al\E�u���v�x(8	o�#�#��k���sxn���dBv�Iq�����l���{�~t���2p�?�X��IS0���E�/���hB9�o��a�m���kb����_����(�z#���v.c�<�K�3����[��)+T��������R7*�u��9�j��;��m��05����Ԭ�c<�n�v��"$��e���ʪC< ��
���Iv(�a8ĥ��.=�xZONRc?�ɉ��ʱ�<����]@v#D�
�	ߦ��nW���F�aHѥ���\���̚����ǃ��HF��C���^�2�?��s0�!���
�[n{P�T����V}�OV�Q���8"�0/�����c'�����o{���^bz˪؇̓����*��[|ZN�6��b9�� ����f~1�ent�.ʀ褛�n�fou#ѡ*m@ �%��p�-2yj���8�`J�J�����f�^|�f�d1�4W�PC���D�sXv"v�/BR��K�7�F�4{��Zsq��m)t9�eŶ�8�Q�X���H
Z���)�`I��98����?��ߤ2�E��c��TѰ����p�+��c�Z����<ph��i��$�3g���)�)���B�� �%�
T� ��9\���5<N_��ė�P�S`�,J)��h�{���]mL"���݉��J��� +�ZM�8mB�mv�8�~��&*�@#x����& �{X��@X��P�HJ�N�hA�'�E��7/�gJ$��8C�6&M:��;��/.��R����)wD�pz=�!\ƻJ��5O_��7mG`��"��	>��Z��0>�M���q����i��0�C=u��譶ZJ-0�a�0���5���8�'���זC�}�Ӕ�yM��*���Po�$�|�Vƽ� k��3@���0�an�%Y.#��%�q�a��C^Xq�f
�s�!:+e3^�iO���J���RA�Ҝ���go�1NYKsv��)�?��Jk��d�b9M��� n��d9��E=A���/��׮X���!��8�U��K��=�}��q��D����6\�k5{�DSOS�T*}��a��6�{���)y a�-�C~�F�A���ܬK��D(^0���,S��3|�V��1R>R��^7�7ؙp��5;ǝP�)������"��J�[V�ż�PY��u�
�,N��c�]	J�؎E��Z��y;6и��Hw�n�$�8�2?�b1|\��:�+AJD�e����DYd��`ڱzG_C�k��` ��6j�4���N�<v�����z�Rɝ�c2C�H-c��rk��
2�3�T�j)u>���.��\	��M���=��S�ߗc����M�<RÓ-y>�ד�\�f���u�������2Wظa�
�mN?M����Q���V��)6����Kcp~%�X�@F������ᘪ�G�^K}�n� :� �!�`$���%9-�I�5Hfq�p��r%�m_��-�e9��Ȇ�	u�D�7$�<��H���)�+.���9��U��
�FQ�������q@�wY�RжsY8.1���� ��H\�K	��M��RY[�x���
��y�6���*�F��:��#e9o�!�x�x S#Кv�@�w�寅[�0e�����u��p�I��I�N~9Vb �^�z���pd�\ΚP��s��KN5)]�t^�l�3w����[p��?#bE�@���d�v̝l:�,8Wvƽ`�S"�&i�6�ԱH�+��v�x��LA��>[�[�a���'�`_��&�=NV-�}��)x�,Ȁ=*�"���D��t�{��W���`5�h�:���Ml#t;]��X}�.����������Z��p�JّF����ɛ����������L���[��v�]�:��C��-){(N.V�s�F�����R��߲,K���&t(۬|R4��"A�;>�@~����2���D�0M�����p�:
�'��!�h�r�\�����Ig?�$]Im���d]���N�Ơoz�7��[%�3*�
y�u!�Ĳ0O�׾�/���>���^�w�i�?��E�H�V
-�B	$�뚚�K��Kp�]�OS��R*�W��'�C��������>QTeџ�6��."9r��ݝ�{� e}�(�.i�3��t\�ލ�O�O|������S����q���R�{��05��R+i0�e;���K���`g��(J�d�毷{����飒'M-�D���ƫ\�+��쾀���Й̎r�R!wa�ĻH{��aذX�O�g������ ��NR�˺ڌ)˱U<��e+�<�O�(�=���X�0���'�n�|X�Cl'4���ǹe�,������٫��X���^6Q'�Hq��oY����A8*ʤo����)&�5$P�X��$�0�� ����ui�cfe �Tc��C笟]�Z�(K,5�uw
��öҐe��e��Y�yB|Kii�Y'0���ʲ�p!����=XW����_��[8����� ��r.!�f0����(B׈~��y�`�ǰ���
��'&o��%N�[ђ���g���P4t%��t�F(��y!�L��y\`m�G��5iYҷ*����Ga�b���dni��!sY;ǁ��az+������WV��-�nx����,�]boiv>�
��aQ�n����z�V_6��RI^�`�0��*����s�n��v���� D��h?��l�b�`4��pO�_�hu��w�!+�Du����
����m�0�
i��i���e���`�����T�lqI����y��G%R'��M�5��${����-&�2�i����:��ߣ�E�@L���݆�*.�V��,��_�����3�����MD��ֵ.��l@*.���P�G%+|��:�0L_����|�h��Tj��?t��F�Ru�K�#�b��V�k��Jj��7�B��/"���U�c,�5haaTV�*�gl�I��HL>���ݘ����+	������ž���N�3��!���ߤe�Y���(g�?�����KE��	z�W�7�	~������.v�W<C��Z*�5�H%Y�B���]��pN�U���B�n_��n/�F���\lt��m�ю�a�F�2?Ob� ���|Ñ�)R0!6*Z�@�lV�ϙZ��u�s_� i�=K�`������l,����.�}���`I��́�f��<$�k�?1��	?�Ɠ��(�����y"�%��/z�F��P�)o:9�zz�^���p=*�no��K�\T�ո��6���p��@��]���S��OR��f/��K�[|���6�@8�dZ��,M��><��o�^e̽�S`�!*�RX����FP�::wbG�:	�/�N��V/�u0�'��A1�o�Y���	d��j�:,|��n5�K�ÚS`�=ћ�O@&���Z�Nd[���FM��{��G��\���w*�k�oED<��X��&��3���"O��!�1֬pAo�C���FR�p�],�N�j_�5�{�n�-y�"`���h|{�f\�p������w�ti��6��In�_��&�٭��
��EV�:����k�֕~���]���H�� ��i���J;��R3F�=9Nl�G�p���_@����A��.CU�nn~��9��3��X��'�������<c�K�bY��{�/`;�Pݞ��Wؾv��P�仩��D�"���ձ�o}�[�P��A�ܳ���4�����'z�z8ӂ}9>��a��V~���dz���g��#��� �j�K��;�M�U�w�WɱB7T�:���5���,��	���	A5V���vk��<��0�쎷x9+�|�<�x��b�|�;�h֫@�$��@�KУ�>�B�uW�aM��?�i��!�L5�Q�\��W��ZE,���eP�}k�Od�(��W�)�]�޿�iO�������7A�7B����bH0t�^�"ޣ+'�ۢ��u������w�����`T�x��	J�u�ˢ깯T/#��:��S�����Cx�q����b5+۫�Z�2��@���F��ylIuY.�"x��w��z�
3�`���`�YG�0�.J`�<�Z�[��K��q�����?YQR�)E(�F&~~}9����eGI�K�W���;�JY["�h����g4��!���ϖ�9�z�8���O��[�-C�����魤���1�5�Bhم�qp0��
X`���C��м����(���8'6ױ>M����z��k��۪�<�OP��ڶ	���$�=�oc?�9UO~�Ix=�w$r3k�j���$뭏��n����+�v�c2�oC�љ:j���;�\R����.ӓ(��I�������3�=e��f��z�(�QW�����~�"�t�IA |�|Q���������*�I�\��<�n��ˍ���(�W�#F��[��ɳf�z#w�?��N�����r��Byo�$2+?��T���6q^��g�Axla(p�Zqa��ҔM��h��1�g1�����E���w%I���I���{p"z��	�*�V�,�@���*(�k�4�Q���gM��V��5��T�W�܀����8�;Y��z��qX�Ң�%'�Kz0���+�5���m�TԔ�[�����Y&0�L��/Y v4�d��l�7l�i�J��~خ���W^�)ȃIw�7*��mU�>��(*5��(S���F�?T�L]�M�3��s�uâ~�׫���t2��ye8� 8���3�E���`w�rt,�ɶ׷s�E{Y�N�V�w�?g1��u�~�U-���SD
p-��(��UN@����;�Fgdm�Z�A�ꬅ�V�^��85��@=��+��n\}�����O���=�lH��7R����C
�ו��
LS/��3�de^�Tx~���H��@`)(�tqcا��jAN7����7�KOpS��qt��d�+��Zs�����Mj��鞓���No����CU;v.��2��h}��d;h��p�\_5	��Swge(�,d�'(ؙ��U,8q�[BE�T�pH���pmƞS���	>���6���a�;B�i�~S��I�
Hp�
��:S-V-N4�P@3(�'��Sr��@#��F��=�����nd2�<��@���7:�W�)q=WTg��Pk��P$�K>4R�6��1w]��~;�9�'�'`�����i�f)�S�j��`�њcm]�-�v�
���A'��B��NN��w��F�	�<jk����4�\�ۄ �
"��f�im��J��jO������aMF�J������C�
<�!E�-��=�m47	H.�O��v?of$�j?�f7�HI�bד�Cx�E���\X�|'uN�?n�܈`?�B�y��F�����=s`X�t�$��1�?�tu�����j�%c Ǫ^.+��V��N�Y�mKai���aÝu^��F%�!q{8�S�H�jʣ�XJ�{�?Y�5��h$��â�'Qs�ML���&
	�6 V9� �[�]�"򍸗�3urBOH�ّ]p�^	&�)��)Pc{���߈�>��ST�<L�%�w����`��L+I�aШ�%�����R7��Z��4�Zѓ�#JO7s�����)�����;V{���:mY�˓���r^�8Q㩨N멗_�tc<H6��c�p#Qz�hb�1 <-Ϛ����䧚&d��	��1�_ ���X"U���\z��'w �߻�o�����ɒ�LlM���|E�L��H�";��p�\N����k*��l�@���{�5n�I����� �ӗ��?O{�ޤz��dT�0�I�R@���+�TI�1vr�PT�X�n�ȧwn��z����a#���ՠP*?K��U�� �c�;���s�����
��Jd��Δ��kī�?�J�(.�8h���'�+�}�m� �)����v�bf�#���qlz7KN)�(��N���~��>�VEe`�;sz,��E�N��������ʌ,7,q�ȁ�Cs�-5���0� t+�T��Ww�Y�a��]+?@i|�z��yS2'�����RҖ�����a�`[�ι��[@ڛ��́Oᴕ?֏�����[B�n���/4�v��եi/��*@�� ו���}�.W1������{ګ�\|�m.ƪ���F��������)��1!��<�	��*�R�LH�u�(LS�����9��oI\= %<�9'�Jv���琟z�\��6K�w"�f<�R��K���:������\�^�N¹�dŘ�W	�	݅W���,����^�u�Ҍ ȍ�N���y��chY�=���|S Qn�%-���9갤�������(��S�4�jAt�{7a�_&L�U.����:,� <{�������6���5��1���tb~c�a�Ju�8�APZ�%#6KV�=��	�sw�����lfa���;�d�?�Й��0F�d���LeX+O�����V?�G�="U���;h�5����zn8��|�[�Ǐ��A6�R$qt��V�&��AUw�V��}�o��Q�C�>��A���˗4qj^��"q�[
�J.���R5��{�Ե��>)�2P�ԅac
<T~� �jC��U�.4F�iWwQq2V����L�`7�s8��,��:�-��ވግKc��#
%;�i�g�P��fL+C�EH	Eޭ:'<�<7�\|��N|��GN�~���VR���2��ɶ4�XxR�_Dȝkz��%��'���Q.�3�M
N�#Z(�q�S���ia��[�ߡl��$�$1��z-����;����C��/����}v��J���,��'U�a�@�����i*&��K��x�l"�b��G?��ݡ�f�J�����xN �5�t�T���>h��n�Ċ�Wm��סSsq�~� ����=�Q�]<�7���1��#��nH�/��v�j���q�h4�tH��̪9!�W<�>7%qb��O������7�y~�z�H��*�=��7�v+��6�Ƕ��0�囔� ��������Fr11ځ�~��W���m&���-Ł�Ϩ�~��A�4��P=��[_}���Yvq��ī���}���5� `�E8����~� ��2c��eغ�j����-۰�;�M�d'D�)�P�)�F��4�5�jh֑G��{E$� ��~Y�*������F��F'��"��H�|���p|J4�e[o=����	�%߽Ң����&$�'�Wl�U4	����A�%��/�M2��e��$鹅�I�;����ʷ�t4 
P����`�=4H�I��̜bW�ϲ�h�$�~՛ּq-ԈP5X��HND�l` �d��ly�"+}������
���Q	Z�/�[�^ݢ�nunP��e����v+JH묵���V�R��{�<����^kM�(mE�<��O���xN�u��Y�s�m��;$ͤ�9��ا�p���rU�����vR徴K�^�E!��
��W=� ���J����d�g�W+�L�$z&�$�^2��f�5!):�.f`���]�4�v��8���&�HS��L����ӡ�hiǙ.�7�X����EubnC��1Q����&s{[�\DQ����������G�?E����7R*"���*�:%�T��A�M�_s�ǁk�&O�&��Iu�Zw��j/bH�&<�U�"?�\ɻ�[����!��ct�U�ǜ�{�T�{�8~����׳�2?��:wT>Li0g>	H��UE)N6�<���n�*n�<[�"-���4w vC6�~�B�o��M#��
�QF_�9���3��B�}�:Y`���6����Zq��  ��,���M�e�!��i^H�}4Lq��%�+T7:� �8H�M�'�5��w�-A��vH��M�&]���sA$���i�q�#'�;�����fXjg ����(�|~���߶�ќڏ�.$D��cu ���Ң�Ml�X�O��;����b>����C�$����U{ �A;�YH�q��3����'��+���n�X�ҏh��F	�W�"��fn�o��u�f[�ļ��x��0ȻI��t��Gq9�`�2^k_N`�j1�Շ����}� sg7��yK}�e:�8*@7��@��
!&%���R��Re��f��<�O@��K�e\ӗ�Kx�7�d�� }�p�a�.��b>L�/�M��������;�v��{͎�!)Ŷ#���l��D�m�ũ0�X��Ǝ�1a�	{i�Y0�ï�Y��?�/'�"��YwX��Y��|Z(p���e�p�&�K)��[d�:�kV�˭����N)5��,D�('��y9ǔo��w ��k��e�)g^s���"�V�ݿ��;-Ǿ�QNޚ$vs��b��P5��t:�U�`���E����O�_�k��ue�f�Ƴ3r��P��g���ш�SE<H�e��F`�� �_|�F��fo1�P螿2/-<Zrp-r]����:���&V��O��<�Mq�h��~+p����!���m	��kNH���/�<o��c�ts�º��56W�a���ls�3�H�]b���5����C�Xl�����C��#�^ț�dnv!��*���1cK���\K�`ݧ`��p#�nT����7��[�-Z(pH�	�����6l�';�k\I0�Ht�r˗���d��p��+�p�m�@r(�<��U��Y�E�R�u6��O�'���N<�j�fl��0��ǒ�i��O$���O|l����%x�%��9y�u�E��X!_���R��af�2җ)���U#�(,BKLS;�u�P���(��q����ڑ��i�^������-)��F�e7]�} ˢ��~��g��P.�Q�Os��Hu�B|w��Ӥ�W��`Ű�yO������e��w���%#4㉟v8�-��V)��9,X�U��'�Q`��%�˼�.`����Dh�BJN��&N��u�Q��&L�E�\���&��n�� 
?؍s���wY�
�WaJ���(�ʹj�U2=my�X���g|�� 5$3��5��$]3��s@]}���ӿ�	 S�Q��7?b��}#��>D�U���҃fuBjă��M��
0�G'�;���zŃ���!�X��TԶ �Һ�_� QP�O,:EN���H
t�|/c)��мҥ��q�j)��޸�mѪ�P�ud%�H�hI"'bZ�i�ybq��cu���I�+L'��bcΚ1�r!�W�/d�C�s7��VN0�4I{�9r�������;?�l �xF�,>���-��<*@Hs�{��ȶuL]�GP=�q ������Ó�Ƴդ,����3�L��M2�F��,5���<_�_�@q�^��798 Z0����KN�I`#>9�=y*kȭ��E੹>s�a[���=����>�����qc��A��w ���X�Bq`Ltɝ�d��"�*�ct������:�6#'��y��Se�o<8r�̏U;�GHD|�5���M� ٱ�4�P��g��3;�IC���!�-���v=� ��ޖ���fRw��CL�� ��Y�8)V��i#�{z�ۡ�o���/|�1�S��+�ݩ�g��L��� <I
> :x��T�̃���{7��L�3Iؚ���.ma���tކ9��;^X�[T�j��d�1낖z��P�D�I�e���nZ�f���s��xK9ӤM7t�����S�Y��9�<��q�=�#�����R�
� �.D�>XQ3��rv��>�E���V��j�R�"~���R{�kK�8�O�ʇM�IM#a���ӗVJ�B��;�&@h=�k�F�U����kpY�+����W�0� кo �)ѵ�aɧE�#S�$�2Y��`jH`����S
�9�R�&ܯ���q�h��ri��9�����:�s�Stc��U��B&��r��?��.d�(E�EKc؈�����aC�F���&sX�r<E(������\g�� \�:e�_���z��u�81��8�,7L��w{�ϖXI�|����As%�B��F'�~���)ws�6�!����3ȺS�H)��n��S<�O�#V �;I�c��;�8Q�!m�ڪp�ς��(Lb����[�S�[��pD[��:Se����`-eA�.�^@����]���� �r�rU����]���CF28����O|��+:�w&3&E��
h��6S��^�˰���׶� h�`> Y��/My�?OX����o����xI�$�ͅ����G���
y@_RUh����3v��$�i�pg!��$������$�ɢ�!⦃�_=_�k�$�c��P3��tB��Us��?O�����~a�l&P�x�i��p�L�=���}$��[��ܡD��5���DJ�9;1XԏW��h=S��O�����W��2/�6�����'�"<p0� ?�����s����s?~�҂e���Gp���PB��������g:��m�z�H���[�*��CS#��(�R1?���̒�\���5�M���k=p ��`ւ���Xq�L��Q��HtfU�,BW�ɍ4j��`���(H�q����6%-p9(=ҟ��x����R5��r#����P�E<�ئpB0�1�HD���<�Fٽ��ղ��Z�Ń<@	��Lͣ�H��D��;|�ΐ]��?0K@q��?_&�g�wO��H!��T��!��/�[H�+��.E�4�e�x�$���8<7V��.ڿ��4c >Y�&)�)���UՅ̊�T�ho��7��W�	J@��X�~F����U�{Q!z�)7�ķ��L�j��V�֣k��u1H���e�Q?�,��pf��M��g�x�������a����!W�JJ��n���c1�Pu�$şCf���H_��3Sֿ�%��'vB%�74����?�`�����]�wwя��"�D���tM�ra[^�$K�9P�p3���ؐ��
�-��Ea�U|)�Nں���~�$,��<��$ėM�wpY��0��C�{Idq�Q�d���kt��	v��A�yK�'{�C�@��
��%
�8�~�����h(���[r�����ĒB�#B��e���ӻ�_վd�
��`�AN%�$/�a;t$#۽�lLw��1���٨���&��6K�gd�Yiҳr�m(9�ףn`��r����4�9����S>]�94��Aڧ�3�3���h`J�*�kRLN��^��9�F�X�-(а�8����Wo��3&�	��h��M��L���܁9(�� Wb;�+�!�B��i�L�<��m��Q圎Y4n$Y�X1�� �.m����g�\_;";=�7:JP�����B��bYJ�0՚��-�5��*����b]Q4l��8NAؓq��h	5I��f�!��\Y��]���0���;;i���繷M��d�
�avҙlY}�=o5~c�)k���}���XB��^àoLq���{�����Z�f���k!��T���a͆�;d-xL��h��v�AXo��.�*M�6�����Qp'��*�%�[P]Kn�lf��p�EH��O$��z��*>�\�pszZ`�f�x̻{z��ts�W���{����]���}�hQ��z!��q�"��)���-ޅxTk��� K��gmuq7�\����G靱U��d��R��	(}��E᮪������������C��Qv�\DF�ח�/ �����B���(>��k����f�m���XL��@CO��X%=X<�.�BAO���}���$�Z��g�J�l&�s`��H7����|��<�2"�h�յL�μ�N����30�s�2=	�+��a���x6b�JF���p���3� ��vE����ZU�k��) �mӔ)��{��9�gcܨx52fA�ٽ'��1Go�.��Uʢ�s�n� ��gf���`��n�Q�,PW����UQAS@�L�}G��0�kI��{h馕:���R9U���r̈́�V��MC��q�$�r�������;�3kI �46����F̗��P:l���3W����m��Zq(���� �d�F�� �E�	!��f�vm�_���2�x�ǅ�u����6dJw$��X�x�z����B|-Cu���o����9��"�K�rp�����W�ivSF�X��i�:.�%lY��Z�oT(CE1D�U}����\L�^��^��0���ޘW�i�Țvt�l����QUZ8`�!-0ȹfɟo�w�)1�l�H�6(c���.�p0����]`*�2CJ؃��Oo�"�;�[��n�Kf㞑���|�zAI���6�-�#�� �8�Ѭ��3�>��<$v�������$�땗W�E�|��μ��m���<m�H0��x^h#1��i�`a��c��Z3��|���U��Z��c�V��p��՚Cfݡ\,�3�a�����X������z����HR�����q�9S��g����$P��?���蠑�~tr���:jF2n��jJ�y��Ny�u ��Yx��AT��cq�Ie�fR��ݎ�~����������s^<Q�	��=t�`"C�c�#w�aM��?v�J�;��9�~Qڣ+<��^E�й���q���2�:��+��(�#�2����j`y�<S��}��m5��Y�`.
ƻ�����|B��&䵈]|��r�Z��h�A�o��v�=1�+.�2��[cuUa�����I_��(���`��-�=��}��@2�W�9)=7�[
�~3]Р���p�R}�#1�f��un��K����.�9���3R�3��˰�;3BJq�joRد�%
Ȏ )�S��pB25s�^�p;!�ՈY��pF�0�L��[�RmE��L��{ x��v9j�tdn���9�V;P�d=i�9�Zb�iX~�_#�S+?�`��

s���М6�����tj߹	�m�?Rk�tY��Ⱥ �@����+:�Y�u݅��;3wv������f� j#� �t-ÖZGN)n7�dz�Et�zrpܕ2kC�C:_J�~� �:���ˣ�(�C��#����/�*i�\Pӣ_��B�U���-���Z�4ur٥��a�)2N����۵��\�+K��I�)~#O��L+�W��Q����K�l$`�V��}����KL.��&>ql�0C�Ink78(C�L��l&CĘW8({\�8X���3z�$:�x���P�T1b=������zA*xj eoA�w`��o��Ǥ���q�r��-9c|����0г�$��~i�Ǿ�k�ԯn��:4|5;��D�gxLo�|��%��m�݄@k�Æ��/��1B ���͹�~��1b��˅�IN�پ��rtJ$5mb�������/P��pzڈ)��&��Z�f�"*v�a��*c���P�C6	�뭚Y	N^ϮH���x�7�*-��[�tܐqզї��~쩓�4}���hI4�W~��Z��``�RW���@Q귿˧_S^�Jm�>����{�ɷ�U�[��IK�����M�r��q/�BP?��Ѳ��~�~)�Fp3������y��\ˌ�v%pT��������
� �s�Mph#>Y|��E1�uY�5�R#��/	/�/�3��!᝶�10�Y2��0���k����[8v����ⲁe�f.;)kv����HV�眊<����\qEd̙�`h,Efi�rKz�y�m����V2gy���X�Ђ�y������0׿�D<�w�����rK'�kIKj���TZp�U�Ŝ���Z�+9��Eo�����+p)� oȞ8?m�­��* �j�`So<���mq���4��yib�<�c� �(�J��ב8�'4���Z���87���(��eQ'?&3���m�E���K-��M7����_~=���	D\�����2U�m=͈���e5���몯q�QԲ9ߍB�q��>����9�8�t�~�c�b�l��.�^l�N��[�s���+W_-ŵ1���Q�7��%� x�*��ٯIEUB�5(�ǁ��)z�غ�ԑ��1���Tb�7g~`ӄ��k��	���?(Q����Y��6j�^}����<1 �Y>�ߍ�hl���w?��E�0nA�%!a��~_�Ff�c���P���P�6z4�P!�	R0��H��^.EX����2\7�H�KN�������H��_T����l�o���r��ވ��_�-4��g ��J�)flG�>� 	aB��,�%:�7+Ia��.�A�Gz_H��[(z�t�ݟ� �%M��|y,��\xG���]<>p� ţ�7��B�u+1^�h��,�!Ў�B��G`0�٥��-dn{�}�j�Q�.F�ġ�5o��fKЫ���g/"�����x[q���$ı���02*���a/�)H&�nND~xR�G�Y��t�U�,�U�ղn��`�-��J�_��4�m|�8!v��%Q}+�:�&���~l	�����'��i�"��8�=�!�;�.��
n �)xy�_-Z�^Մ�4�	AN�q��2a�t�wLE޽w�����FT�m�0��v�c�-��鶃q�$R��<��mPy֮!��ͩ+�z�����ƞ�_êiOr����a�0Uϗ��ZGz�,21�ˣt횒��(<���"���Hu�F�.%�A��bQ���`��y,��Z��f"��'�Q;�!��O�����c�-%ͱS��K���@���Ņ�z�J�D�i�$ԄM�6�Ȇz��H�T,��*�(��|axC�N>�B�������T�jTR*t�rK���#�hZ����������]L��/}H,�j��kǤ�cg�p���I�WNIX�k34 �'oUyf�G?��)Q|�8xsW���g$ޜn��������s���q: �׷�}1>�q�:��2
�x"������M�\G��{�����"��]�%T-Yv�+j�]��CP�I蟹zĠ(@��N }v�Xp�_eS�Mu<K|���O˧�Iu���c+�[Z6�qr1��z`W��x�8�Kzo��!��q|���i+lhww+RA�|�m�l�~6�d0mb2��1�Բ��T�<���#��q��D�|q�n�J����*G�?5��e6�:�6h�HK\��r��_&o�d�Qj��twpJ�	z�A��x0�,���){�m'�K){����5�e$9�a����.D����	������K��0<ǋ�/Tv@;�B>����T�$a�>�N9���	o�P}�P*�*�lT�+o	Vˑ�Y�_6�|���������V��{I!����R�H������ד�!��:����훎ώ�_lM9��[�Y6���H�)���F0Ud����W����lW9El�u���+�~8T�Kq�)�7E�2�%_����~]:��AAi�4ǔ��o�������@�FId����IuG9\m�{9��mk߃7.�����Y�f5��-+�8-?�>
k���!W,���+
&&�Σ��RDz���T��m� D>��Y5����z	�r�j��x(lWm|HUi�/F�կ0��='a��S�x�Y�L�����.�J_/zl�U!�v���E�Y�U��z'��R��h6�$�^�@�t�5m�Aừ�jB$�cAA�T)��;}��/�Wr��6?��������bf9�`��m��b	��O�LQ�1"��Ȳ�K��P51.)�iP�P��^��g߷��@�_J=��>
C��4�^�Ԍ���1N鰦*��̊���o��+���xL*��mRx�L�eÉ�/5H	6��`��>���?��x�.�م�����P����:���"?�Hv��.[�P� ����Q�5r{T��|��k�H�[OL��V�����ᾓ�x�qb���Jա�$�w1��#�Ug���K1���Wg�Z�2� ���zAyU�)Q���KMʗ��ĺ�=���@by1�^. ��D�3Ң�{S��#�iʐ�茋�G��8���Ώ@��� ���T�g��@��ZF�X}w�cXw��+�S$�H0�4��PO����1�O6�n��J\�޶:�)YD܎�YnZ�"�uڃ��_�!���W��A
@#�+�,Q�`l��3 p�	a�֊�Km���4�)B�&�-���*vQ^IQ
�p3A�*�x��%�s�8�e�y�2`)���$�s���`8U�Gd���>ܪ夑4�VǌU��M(^h��a��uΰ�NW����&���{���YD���#ܒ���^��_����I+.����j����A��,yoLIK���K�U���2��mLW�������7�U����� $
%�گ�c̊�1�yg�|���>в�Q�<�>��H۴��[�A���%������W왻#\�(����}�JF����؏����fHf��Ro��[�K��kr���r�h獘�3E�Y�	)�;1�Arc��U�q�"��Лuք+;�[�;ro��n� ǡ�c<��v��_Ӗ/B�����|����.�����]��X�ߓ�a,4��C|*.���y��5֩yч��)���>��7K��W,Y+������u��2�`-����������Ӎ�mx*I�t������:�pA�Ws�=+K�Q�b�Ė��qBU����ya�� A��2|�	�#
0�-b���?��MI1�
�u/�b]�?a�u��V��jYh��5Z��+��u�����+uʫK~"��湇T��.Fq�����vZtH��z��C�?b����
�p��G`�l[��k�Q#�W'Tu6ɍB	�좓���9B�#�I9�߄�d�ב*�Sm\?�X���¸=�K�Б�u�]�Bq��J�R�t&t�&y�Y���"���;V�_��F��������dcʓY����/�/X��=�7 �U��͆<��>5G
BI��S*���J��ও֣(DK_jz�xR�}{�
{z?J��'~������F%u}��_t���d���y��A_����~�X-�c?��2��b���%[;���V1NS=fBb¤$�U�^�)3#h�F�j	���1�BR`��hbӮ:��ӟ�_�[|e��5���l�S:N�&Q�.ᔷ�$f�L�Q����d�G�9LH8=�o�� ��>��Ǚ�i��Ƞ��V��@;R����&����"����1��h�����1-_5�����2�r�#�<������/#Ϙ�zK���x�ɷB�������M�����s"��'J�P���z��m6>=�ipԜX��f���(��h)Y<x ��qZ��#�^%3���@ɀ���'�-�o]ai�<и���ǚ�y���Um�8l(����KTk�WP%c�����f���+��,N��E)4Q���v�}.;ZG�5��z��G-�\��Ӻ�fZ�c�ڶ۸Ӊ��Eb�f֊f�2-� ��d�%NC:��5iA�i�h��:r;j<R�=�Ί�M��ӑ��F@������+T$V��� ���o��Ǝő �s�(ۂF!.�������=*�"1��#}�u����9�k��w ^$b����vrN���,X6/�]��K�ү?��''�k;r�8�����˫��S,�h� ��JO���R�[fa��d@���y2��MC�OjgYl�:���S������E�\�L�0��0q`K̓�~`�y��2K!�M�cw�\��������Y#�L��`��d�:s^�w)����\��P&�mYF��S�@�rx��dQ�P��*�6ȸ��L�;�����Zľ��~���� �'��˸ì�0N6)�L�A�k��]j�u����	��hM�����#|������P N��J�լ/l�F���X�dnd�Ҧ)��@q�