��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\��1yfMA�>bpAo9�f<]B3��SN��T_�eI Ya�R���p�K1p((���*��?�������[x)�~��}�t϶��\؉�bN6%\�~�+���X�+��P�T�������
�lGi
B��}�<�(��{��B�0� ��b��{ـ&e��/�)�L����<��w�~W9����t���8-��ܵ�͑�v�^`�h�mרɤW?�R]O�8֏�$��:H]K-�T�!*bF|�޴8������舼��s����L#3�����(�^�6m�ˊ��e謺��	��C{[E!H��G�uPY�aY��$]��GA�M:|~1.�y��y$���@�������1U�d���&s�:d�|=�f�mp������� |q����Ύ�~Fe:�u\�Z2��l�iwg*�7/�n\�#�/:;�c ��Ň]P�kHϟ�DZ<�<�.�9XYb:G0�p�3��}�96�i��`O]��m���ȍ������I����JZ5B�Ȏ�	U�(m�?K����b���!9�U������)0��x���X�8�;I"���Mf�Mc%pԅ���Cx�ҥtνXq� p�'ħ��'e~ �gr�<��YU�6|�W���}�!��Dq�T�NpTR�0b�E^�|�<�<|� H�eO]"R�9�^�^0ު)��Np�=����	��dv���qO|�bhz\۴.�%G�=�TJ��d�����uQ8K/�1rQMc�AK����JU�(8Lf{P}ӻ��ʡ_J�ع�}��qU.��7��|��l��~�t����ҵ�~�_u��ѷ�@V ����o��#��������9A=�`$�ѐH�<��h"t��dH>*Mg��d�,FB�o\����Ӽ��d#�:�h+�U�=_�.0���^��}���H;���؅��Bm ������h_��3|k�E.�hʸjS56ۂ+i/��R�(�v�ς��4$4�Fn(qD��󆷲/ ϱ����©�w �IA�|�����[׫%�_(�U�%�8J���7�S;�OКAE����ɋi����Ƹ��"NX�՟���&l U�!�A��r�t�d�h�����������(�r�7�~��[� �)ڠ�:
����\�;�z�N���N�|�d\3��,���CM�e�s�7f�	F]Ӡ>m���[] �-"�f�f-�ԒQ4cԖO���,�����V����m�������s}赗v�c�Ec����y�\�5�|�P2�A>�"��=#i�ӂ��1�Z�>�	ۀ�2����_���Fm�������6���.R<+�����ՀS���I�I'��J���|�]-��di٣������]���_�ivm=y�}?�|��4�)�z�:J-NF�?��!�^9訠}����?�0�&�D��0gӋ��"*>މ�i�=jx�H��������j.��	��G"񀖸u]'�P�f
M	B��
}������Q��[�#��O� (��w�V\&�n�vA���W�����	�o�4�᯴?��O�g�²p�cD�W�f(P�h+�q�y!�9#���k���OQ]�����e}r�q�!��3����.`.�c����	 ��?0 ܾ�:3UÞ�vL�	A��/���/���q42-��I��Ľ�V�8�g�V�?����æ��Q�G��#E��$r�44�ۙ��*���/�U��@�K6��Q�{�����צ*�O�I {~*��tc����a���7`�1	��x�Ebѿ��t�DЫ�\��)3����ʊ����#��R��:ǁ�Z�R�. =l�&R��~�8��`H���0z�Ù�u����٦g)�yݣ�4��Ҽ���1�vF,�[z*_��O��,s8����!�r��-o���X8@ZT[��4�1���A�_�	�ހ�e���Gя��Ֆ��6���یkj�N�,��^8^F�� *�Z�5�!���t�Kt�i��܋e�r"���I/�"[���U����?� �0���o��IL�ڑ�G��������Qh�]W���H�pR�Uz��yY�=e�_ʹ��s�T�Q8���y��Zq���hp.��Re�� ���B��U�LR��/Ɔ�����npA��5P蓪�w�X�x�
�\y��s�c������J�Ѕ)��|Vc����k63��5����jqϱ���g�ҍ�����4o���h�
��>E��n��+�:��T�s�(W	=�hǗ��|TH�K�t6t�
|��7y�0C�0mI�+�)º	'����O�&W�!2�4 �Ӎv�8���u�����,諱fս����f}1���v��- ��\W�8ρ�p�ս���]�3Dޅu��g��t7�����+0�����xy���k���(Ŗ�Q3�,VS��jcɦ��LPU*��Q?�iĖ��J��h��EZ�)A�������q�R���"�ە�e\4T��fh��&�:R*�-yܡRj!w�%H��|,�=�hey��*(��8���`=�&(���A3���
�>jӸ�U�M�5�;<��t���Z�=�tn�.+>\f��}�I���Z�_��s+kP��Nf4�cs��rFs��n/�A�0Q� 4\����Z�KЏW���k�ld\J�O�=�����h�2�k:XO�2������h6}�G~�>�9d��aK|ʫ��Y����Kzo�YpD�^�"0y�`���C)��4٧bHQ���QF�3��E���pH&lj��e�;�F��,��޲�K�B	��=����c�r�7�tc|_���q�����F=����u��S�5���G��Ԛ�A)�4�d��� �6}��A��Ԝ���pyxd}�CM��yӘ�p��5�5�=-����r��Ã]���f��;�#�ء��"Xr���l܋���	��A�\�=�_��ۺu�$����(I@I�S�Ȇ�����|���J<�MZh1m��mOA�G��.�p��:]�8���,l��[v�,B��M.�Y����z?Z}�r�/��%��0H�'+�5�JIc�j ���f&��#��X��e�"w
��S�m�r��W!Z��>���%iF�x�N ��6�?6�B��G��q��/�B�ns����A��ͪ��z.�	�c�	�ُ2��ae��ww�4�P��TW��˖����`5�+��8�w˹��²P�� �E�z*�?�;U�\W�'ԽD�{a$
μT(�o�z�8��#���j=�0Đ�L'쫌\�1y��Ά}%B"�҈����Ib5�;�^��x�i�L���n4�_��I���_�L�`Ny��2\��BL#��]��ć'�`)f�k�e��{H��x	�p5 K�m�1(�aQ2܂V���ڸd����S���/u��@(2JY`�@�q@�n�{��
�4��~��+��I�HIw���i��ݦhi���؊�s�w֨S��R��	���0�ͷP�ľ�ݴΧ�w'��g��ퟸ�a7k����ť3�w��NaW9����z�k����vW����ND����D�ϋ#P�n^���}Rׄ����
�N�pF��@��E��{t
�D�P�1=waU��J?����-���H�����] z��>�*�:*��4�.�~�pY#�.%�Lz ���K�)P��0x���lx/lf��y!sG�DEo���<AF��ɩ.@��-�|%�t�eVƞ�%W��?��'����,?�S�)W'
��M��U��7�Ü-V�I��И= �$a�ײ7�tlĚa~b�ߠ��>P������e�ߟ���矨�c4Ŕ��t���AI��WE�4e�қ���'�3�p|�׳��@%#��s�K��|� bi�̜�(8P�0rFI鐒���&��-�7�k��"���!�<l��lB	Y��Ϣ����LaY����&f㈆�<x�l�!���`�A��! N�ڑ�K�^��^)6Ҋ,�t�k܎,N.�}ar8�M�1��ۙnd/�A8���޼�����"�H7�� ����]q�����=d+�n�܁�86���Q��Ȥ�]���iM��^��ѣ�$vSs%�>a�SMs�	��s��S�=���I�ޖys�����n��C���\�϶U7�\���!$TesO��Z����8�I~�Qi��Lӟ��i���a����O�/U���6����E�g�1i�G��^}�
C��)���^=���2N���]nؓ60\/,hǱ�o�05�X\�%����m��U�[icR0h�f��!�Z���ۙ��T���-՜<����\��s�����2�Ey���,W�Ehg	��SilÃ� �o���\�� ����c��w��]/֏o�2z����Y������'Y�V}L���Rvv��$�[�]���װ�|ӎo�䱟��a9�5hP��8�8%�^oߠ�u`L�X��df8Ru	I��r��¿��
t#g�NdyΧ
�	���f�u��Z0*�>t�����BF?����^Rt�p�����X�@�c:��,�,��4BWw>V�Iު�1wz�ֲ�|� �>w�5@+��b4�|�wf�Z��D��G�����S|�Xp�Y���
('��e>o�p���~k����ި@+eÄ�cb�s`x]H��549ނ��/C�x�O�t���[zH0T��l��}�pj�z��W��(��cWX�ۦ�Q:���ˊ�����o��b��N��ă0Mm������@E�D3��__��Z_aW%�V��h�֥ ,{|�{�U�����4v9g�+���H+���ku�Z�]��T�g4>�b�Cb�&>[ws��*��N�]u�Q����B�	慕�3r�\�Г�_��-{�<J���G˴��ˁ[7^&�
�e�:�^��h �b�5w���b�s\�:_�MUtZ�ҡj���L���e(c@5x��KB7ϊ�5I����XCa�ƚݘP���,���+Z��D;���y��k:p �v�_��,�(�D�ڑ,�0!�h��YM�L���#��!�^�f�s�����~`�('QS)ERz��~�~�$	�}ҭ=K`�م���7b���������D�d��[�	�fe~\sj{-�%�l�o^�rr��y� �|����y2T,�����8^8ڥ�Go�/�]#ZAQ��q�j?1o�»�~#0�+X�ChMڙ4F���]���]B�ߚ!�H��FYn��Ќ������WX�x��S%����R���D���T�i�9��R&8�����i<�����kN<�q�e�u�K��`j�cs��O����1��*��gf�����,�	���HyC����c +�5��e�Hl�g���(�,t�~��:0=)e��j����H~��E��N6��*u2��Ϩj���Pc;�r�1���/i;�� �?Պf���)FzPTZ�jĉzc+ ���M2q,"�PDC�CC�iV�����]IWu~�k��;ޮ2f��+��N���%c��%Nގ�MV�V���rO�Ұ��!�.���{���3u��%Jt2^���:Ȭ	|$4������~c4A(+-[0�R�O�M�i��%;O���I��Y�~gk��@�����4q��a���2
Hh���SS�<�7!�2S	Hی�y�$k���-�A:�y��sO����~�*����*V���C��8����0u�H�wWC�pd#���ր��6AjL<8/6�q"��Q���r�5S����i���g�L���~l��sR:j���(�Ee���탛U���_�S}�[����n'�g����G˘k#�?,�7_kp�b�)g�H�z�ew6������ϝV�ѽߌ-r�� &b��������#�YI��P��~9ڇs1��<Di�l*Rj�'�^��l�ზ�=�y	��A�z�[�`G���Q�s��:$A�u�n��G���`�ߘ��E8��3�Q����.�>��1}c@�����V�׭S<.c�͓�Eo��c� 4eI�
7.�0���]���-9�?+�.� ���:<���<U-�uu;m@��q�Rz��`�/�Ǹ�x�n5���?�!�!0�޿�j,[�4�c�ݯ꒳��h+Աp���a���wM���'Gs����sKK�n:E�sd���R~h2�C\����Z��������A�@+a(ؙkf�eOޟn ���{0[��pc���36 �6n�(=���>��FD��p�|�&��U���~I���j�#z�b5(i�$���Y�!��ұhK������8�ROc��n�x�k�����ucp��]vROC���^�s�O�����ốL��VsIp��[u�J�a�񩾥�����w��A'�ޚ�R��$W!jN�v�h��"��C&p� I�LQ��ؼ���}r� ����*�j'�H�A$��Ȯ�qY���Gn`L� ;���ޏ:2l��I9�=rzߕ"/K��
�)�Ǚ��bf魝�8s�E���P�n��m������(R�J��6�tT`x�\9߷�Ik>,��p���Y��	T�����Ȅ��b�5�����Z{���O��Ki�v#��-gU	|ҏb�d�3{��a��x:������)y�#����d����M�/��Iu)�_�����Oa�L��t'��_F�y��L-�����é��b%?��SI]��uIȝϴt�5� |'@�Pl>l˹& �޿��t�I�����ׅt�
��u����k����?M�O��^�i�`>W3^���,���m�<	���m E4�޿��}��q�7܍�����zX��Ԡ�i�L5�o�I�)�_���a�Om�;�D�'��xm�,�����&����+�숲�޻tb�v��GC�u��FV}1f�Gߗq�$�ZC�"j�����0
�#n9��'����/�E�zrv�K��������f��l9k�=�����E�s��*M���d�#����� 	�ژ̎dݗ�pDx<��Y�(���D~�AA[�_}�����o� .V����\�S���Q��E�¬')��'�a���dI�?��`e�>����Ɏ7��-����<ϸ]e��%��B�l�C��2�a�xUz <�l�FR���D@s��1�b6L#/�M�}�!)x/	�V�\_����Zp�-��Nj���y�w�羏����Y�����I���hJz��� q*K�R����k�۲�h�4�y'��m�e*	�:�a�_�jS�W�RO�Pe58;�0~ �E�D5S��~�v���k�������袕�����I���d�>���L��;��:�kS��Dz�>{��cV܇'Ά����R<RTq.�M�n�0�-u�x�>�MB��c وK#!Il�|�\�%�?g�B�0y�;�=�0���ۗ�����:�"�3w��Tx���+f��Q)�75,�W�b#�*FsX��O͟�e��G�`�r'1J�'Y��s�nY�n��r	�ߨ se�C1�Z�^5�Y��Nh�+�V�k�HIݑLȾ��.�L�"잒���J�L���;��SB��F�%Ǥ������/2;Ծ��|_�N.b�SW~�˶�/�
�t���V��)���Զ���d45%+�S�uT�R�X7$F2}� t���z7K���BJ��y%@���.䇍2��H��%��Z������ ��W��5�����6H�4�S�-6��z�����i|H��T�X����� �[��$��������RKX5�U��W|d\k7�H�AE����`��R�T��������KK�H>�6���g��4���E�?��W�BjF:�ӓ�d>��ӕ'C���
��� �'��ݯ��)i����,��~9��th9������-m������P�z#��l�/8�:5��� ��&Y�ψ�b�1
ʤ�DF)Q�C��k:׷��\�Y�|���~��h��ې�R~;�J��E4�(_|eY��#C�j�\_�J�d��ݱ;�̰�gˌ�w�q﮳���wD��5_�S�`���CB�}�l4K���~�]��.TI����y�罘�_9	�C��3Wi��f�m�G�#s��\�a�� ��u #xP�\Z�pq�/�#�lÌ.��[2�O�f�ڗ�r~Tw"�nwrxu������\=�9���P��9�|<j�ҟ&W訔��a���up��'w�[q
ώ�z9�rP9WA���K���(�V�Q?t�Яq}��!Oȃ�d N�J���}r�up�ר����F(f�՜k����&@���T�ڎ�b�&y�.e�gL���	�������%�KG;��@�g¬����������z�s��p�J*�y�j�-�86�;YOu��n)��$�n�F�v?_N�*B�~ARw@�wW�]�O5���Ew���p&	�
(��{�b�q��J����� ����p��?Vif ��2?W���م����SI 6`fY��F�j�k�:(�*�hy.&�4��HqFN���R&��R�Ι����T��:�~��j3�>����8/|���e�ď�Dݳ�S��<y`m�^��wL��	j�3�už>�NP�+,��`�Ж�7�����G'H�7�01�ǘ���+ϖ;x���>56Z�+<=��RT-��_5+�G�)P�L�!���!a�]��ͷ6P�J�m�� /'�ņs<4�#� ���,��M.�T��u����mVI�%�:�d�� 뭫rU����/v���n��v$hy�$b�p��:����+��wt�l���m �j5��Zu l&G�4����m%�X$�8�(6���'�J�Q�ۗ3�J��g��W�(�!��q'�fr�seNd"�'����0s�l3se�>�����!�b�o��kgw������7�Hӫ1�zGR���گ�	�1��c�a�Kk
l��8�9]���Ƹ8��)�`�v�
 ���%�m+y�%c��h�đb�M���Y���	O�n:P�p���t(��\�ݚ֗[�W|D_k�|�y��Ǫ���%�9��[&m9}p��_�,���?��@=�xD�����O!�����v�y�� hB�5�-�	�{�C���69�1]i?o-x&p�����iTѩ��c�8g�-��y�O�.�h*7YL���p����8�X �yY�Iw��]�T�[�+�\3*�o�o���q�ܹk�q7��*Y�g�9;�r��j=?�/�g����aFb��fO7
/uW��闩�I�wǆ|��o2�t� z�/oˑ��hF��1|L�~�Y���~�L��S]���'��E�Ş@� m�a����s��4Ɨp���'7�)<d?����ePPy$��>R�M1�w���'ů�r-MG�dVq0z���<G�4�������=g=	>�*��_�P��i�!F�g��#J���A��N�"M��:IV��(�ĵp�՘	1�k���lv��b�
y�a��D�"��(�-�w�'�4<G�k���=��W����H?`��h�����z���0�����jl���o\�_���	�;�߱O�:��1�ة����J�3=�y,���W
M�p��l�H�hB��I���m�]%�C���P3�r�{�s��s���b�]Wp��"/�����Al�N����ӹr���әi��&�*p�����Dm������PwQU@-G���X�����[��W$�n�'��}*�Z�jv2�d����������ս��n�
@�Y��E�h�ԇٗ2�����пK��гAu���{U�[H�W=���BV�J����CBA�F����{�r`y1�!PQ��f�$E���M��AW�]�9��<D0fFڪ����yޔ�+1T�!�)L:~gy�� �Xb�x6�|�V��7�ncΥ�쩞�w�f����s��ܷ���x:�&oi�t�X����s����&ݬ��F��7�%�=��!���A���Z�����KP�A���s3�:��q>����?pX:�����V�i
=&|��NUsS��p��qb�Y4�>�@,�uǐ� W�6�|�z��}|�<�8�<hL��z<���>������H�nU\�`ݻ%Z-F��ڒ���E�/1��`�Ħ��P���:��6�<�B�;M���G�Fɇ��"�����(YR������gVF �T1S����[�F ���^��,��H}0:��v��$i��f[a$���{��(�6��4���c�{׹�f��Y;ɣkB���#�����51� �b�JQ�Ee�'���B`Hv�I��9ѥ����fB̨�:�`	:�WU��k�)N�Y����f�y���Ck ���@�g�H��rr�졎n�}Ѱ�X&>���?���uS��4���'�S��w_��;�t��C+�F��E��Ϗ��*T��6g���>=����2�bGGx�4�z��c�,�r�0L�\>����a6�ɷb@���ZI�*��:8_gͱ[F~%z�T���� �l���S�a�635��5n�1|"J����J�S��60(�?�K��ww��Pe;��Y.��'{�a��♭��4감����1UKJ|t)�	0�R�m�b��x`o��w��������y-J�'�V589aT���+���z�������%/O&�U�"������`�s*��$�0%�/�R 2쎾�D�L��ybj|:<\�,#��P3�-�zvث&Ƈ���9O��=~�R{F�
�#x��Iv�o�� ��u�[A3.�?���K%T��-�	�̾� j�@���R���=���l�ϼ����U�pX�Κ�����(;�:���V�90��.~�c?�Z
2���m� 5���'�:�do4����hY�p�gw�� ��� 'n^"����#�e��"8?4�m��i���G�ۦ�AX�R%�?<�}<���w�J[�=�rWx�M���p5IY�+��R��΃;ҽG�Ą�V�4�$��m!l�"�ƧeRq���d*�U�m����'盳S�X�2����Ư�y��\1���G����V�]L�?ގr�Z�W8�|�Q@����\�ܡ4+h7~��'�<��L6�I�Ƨ�CP-d���[���A%�bʀ�2R
M��n�^�N��*A��|ek�h?�<�Ԝ���3/��:�nɫ��Se�PNuZ�
[��p]V���T���H��鰍��m���o`�9�~΀eBӑ���k4;��x7�(���
�	>���ɣ
t���ܭ�WN�s�y�I՟�����9k�䃇�(5����%���������rM�epXU��&��\�9�ΐY�[���������}���J���M��c����ӖU���@��zAdOxtk��n��MRo�_��Fo֑	�$+��bK��R�od���u���0��/���Ö=�"YH�e�lk�,Nfy��g������ggI��6�ұ����N���-���f�K�Lϗj����}��4!����("6c6��$=�`�b%Pl�W1�	���ڐf��s�i<`���v_!q���{���Ț6��ZZ�X�4I�cP�i�"�D��<�e���^�qهJ������m;���ׯ�>�7���9�T�RIAhL��㊃©��)	/0�	�M���y�Gg*ld�ԫB7���M'^�3D��6�OE`��l�d�K��]�#�;2�bR���S��ᗤ�\���<�89���=�:�(�5��hL�d�9���
�(�F.xk���y!Z����Ա�cC���C���\*��x��P�_`�ݯD��,BX)r�2�Js�ֹ��Iج��=��	Q悎^��V	E���4�2�BZ�j���[_'��O\F��
�l�z9<����
\�$�,�w�/K�	uP����)�&3�(e��T�$U�R�0�!!A� ل��b�/�N1.:��{F$c��l�.�3C����(5X; �mzsy�͹�ت��o���'������5	9�9��l�h�Zz�XT�����`��S3�q&�m�n�O�ơja��B�S%\>�����#��\�ᓇ����TQ�RRf�I/��"����w����u�N��S]�3 [�]�	]�/����x8W����|˺��Op����i�V����;s-��i:oJ��xT���P���O��I�L���#3P�uE�W>��5��a��]�5M��m�Z�A9I\Ege����Z5RC�U�׬%�o�h��mȊ�����4��\hl`�#*-	gJ
T�h���G~��٭��್�����|>��J!dP[w�Rl/6"���@�v8't�#Δ�]���嘚��6��.c���)`�W�=v#Y���5UJ<L7h�;�Ǥ�mL3�Q�ȃDC���!���@=nTD�Xd.��*� 9){*WS��ؚȍ0��@r0L�g�vX�)�
�a3��Z�)���0d��P�3��g;Z���}C�-S�zW�N8����iXS|�]Nq��A_�c5j��;L���*����x_R�9�2	u�K�E�4���6��(	\�����$C�j����WyXW���<ŵ�YC�S�すB�5{)�#C�hza�{�H9����E,X7��O�`�K�����βS�?<Y�m���4E�X1���	�B�ڌ�B��4�InU�޾�+9�~��h�$U�©�����xos[��������2��4����ĕ��RP�WfXx��v#L��vX����Z*S��;Y���yp��?��"�ۂ���'�y6���햟���q,�YOu��6ۊ��ⒽP�vt�2���T-bv��� ���|BUd7G/��Ϙƿ�+��;���� a2�+���ߴ���NϤ��5K��d諃N�<<�9r=�/aJ���H5�G��lcf�a)�/���Y��,&��:h*N�G�+�*����5��n��`2��.�@�@����oQ����3�&������d�̳����>	���N���6�8�z+�����{��k�+vk��d.;j�(}��'������BtƺT�8�F!#We%���鵭��S	���/tZ�B�B�Ƭ5��`P\'x���W^D�`�?����94��J�1�PGUI�<�N�����E]�trH/��]S�5K�n�1���L�r�~1D^(ď&�~���Z�L`��)N�M\���G����u��a�G��&�[��*��<�AM�����l���a�<dm�+T��:\�"Y�Q%Xiз�E���I_�7֊�v�ɍ�Ȗ����{:l�6���Ҵ���A'ߙ�4S������Wc3&e���x陦��C�燒�g�bP�E��k�6�n����7Ƅ2�s�}���3�9�@ow!,�򑯐�#nC A�g�0]t9�(iieD�xAT�)Mm�$x�`m�f�֨�������S�w���d��d��A�,�p���U�Vz�eF�f�"wii:�#�B
o���Tx�hpHn��	nSHn����T֊7����c�w��w���Fx�d�/� ��i{�CȺ",��v盨F@odV=�gZ}r�(�܄�S�T
�U��������D�1�g�Q�S��
hu���q���j����\V�����2���4_��l��c���I�y�{͊on*̦�gl���ƽʣ���� ��>���*w�����^8�'�#�e���b�UD���?�/ԏ����
oE69\�c��&lS?Ԙq`��ǡ���*=��:�+p�h)~ <��r�p����)�w�����u�j \����r�����_��	�πȇ��s�t�/i蟼*�1X�~W�u�DAc�qy�^(�޳��ٹE�R�[�(�h>�}�9h.����l�0�������c�G�}���i��q��'k
��/��
�4���g�V1��P\����χi�&�o�7gH�H� ��)�T,A�ښ��?S�Dkh�y�P�잶]��ڌ
��oK�>n�O|���6�/����Ո�Ԫ񻸓&)�:���*�����������&�X\�i�̅�m��9.s��ч�n<����<d����n..^%)4y�O�kH����A@
|WaN�*�}٘�g�BlG��n��X��T1k�t��X��~$��"�Eqe�N�8�S	
Q	�ǽCG�}��,���`�]{}�М��d<T��4ߋ���lI`����魼�h��ׄ,��G'�N��wq��9O*�����~���
�
��e�G���-��D�}0�W�(����*B��x_F�b~��B��I���x^��[����1,�X8��x?#�_쐳U_V`
���t?��r�;-&#V<5P�v�7.Y_��5(��2�f�#XN���LoH@�u��qj�J]D�x]�weF![�aD����{gN�H�
)�x�Q}��.�F=��q��
�%��h�F�w|�c��$�4���gN�#Yv�$��i\3�
roh��67Z�w�=E˷@!n����cml����[�D�S��h�����W����-EU�9p����Z@�'�r�p�$�0}JxjN�1%~��O�r�D���z�x���A:���!w1�5�lO�-�[�E+:�[l-�z��b"�x�G�oH}�N�ig�B���Xh�9��iD��&zSֱ�3>ȩKP�u�1Y��T��
[��+��칰 i	&3��6 ��ؽT]20d��6�
��E���8=$�e,���ci�^�#���6X���ʢVIy�
�7��IY�+kQ|���f�Bt�T�c���qB�4��������"X�Ҍ w�ɤP���b�5W�᭞%�iyK|���7�H�d�0�3������Z')&J����������K���R���5�A���o�HX�p���Г@�Hп"b£WP����3pZ/-�����$��Ű����0��Πg�Ѿ���)�̺36�Z�5m���A�80L-�J���{��h8ޜ�I��S���vS�R�;���9�t3<Q�7�mQ��Jn�I�"���έ@璜Sa$V�{��O�C'�aMy��iw�q,_�S�=�xW���^6�����`�Դ\�����$���,�Gr���6��k���4֢�ܐ�(X���O�(���ֺK��>\���ur�l����� i�YW�M���F��Sd���n�+�{k˽��.��r��dM�˟l�}DuiJ)�J�阴n9ǆ�d��:��sH�>)�e�$Vف��;��sد���H\��0K�I�R��{KD���C69����U��{Le��n����q�n����U)�­��cq>������-�H��p1�`�ݓ۽��1t�?.}��|H+M1��U���m%��]�T!;�x��Q��̰8u�R��`�#9�U+�!��K�M�w-�o��"N�,�K�[2�P���J��Fo"�LC��Rw�8$���;b��.�H�\d5@�J�-b���1�p�ic�m��u��쵇T5�t;�|�_��Ԍ��_�m7i��� [7֔��i��3R
��+��x�Ⱥk�n�w���`ԫB0H
�~���r��#R#�RM�w	����ͺ\<�ϣRE��#�_Z@��U������жo�6�#c?o����-��*��`�IcN%<����iTF��v��Y�!#�g �}];��}�H��1Ovc���Ԡ}�+Fy70H��G�>�(q�H���5#�C�`�0F�@��ڙC0�5;��4icUݽ�t��B4�Y)Et�B�ޚz�.f'�,wi��K~v�yѷ��b��W��\��c�6�Oը��佹L���\���
qjCA����G?��3(�nM��f��z���H����K(�0G�{@��r�+��4;@��Ls��ZQx�Ɩe��4�������U��k6�g5�t���hk������@��9��B���RI����:K�P�|l�k�A���mAn�4@�����}�sB�6�T9�Pg
�S�
dR&�b	�L�UɈ��a��Dй��Qb��8�2s��A+��TYQ�č}��xyv~R=���N���
��HY�J:ᄊ�~��yòIh9�q��-����IJ5��tֆ�:�7ZeݑC�D����Hͭ,��K�hkF4�b*A�܌�<T,#f�\���{�{����Bs�|�17zE�)Y��-Z�v��K���^֘zߙ =7���UD�������������6	���ń�y�3/�c?U~{)�Y�q�.tpA�
^�f�b���u��S[҄��'@�ƛ f�/x�ߨ�]�������/A�(��'��M���6��b�����n@�a�d!I��Y˥��"�JJhW設�Z-�iR�hE�8�}6x%��N
9�@'� ~��G�}�� �#���֏�p$�-�T�aj��"�Z�IW��-��Xɥ�Q �����'����;H�����k|���;u�	k�_���H ��pTK��q���-ڝ�v�i��*r���S�����o��G���:^�窣=j^�w���?�	4E"�!{Q[��J��~�����<���w�,H��p@�D�t^%��Z���(��G��oŌ+�Vs�x,g@^�U0�'*'�{�[�����ƒ���)	͐Wݕ���Wp�yFՓ�����-��=ݺ����2���M��U�X�rP7*�����tM)��V��?�W]�RP��z���G�C%Qb�;:��Q�F�ojw�,D� ~�B��6P���\�ΐ� T;'S����g�W5����Ё�?a|\2��F){��Y�8�GW�X5�9�M�`o��o�u#�]���������E?�}e�����+���~AȹlX��q��j�KE�1�YQ=�M
�~�:���o�?�}n�X't�tPz���?���+�u?�_�`'jjOպ��\nkD�}�3�B��<��o��.{�$Z���:�W��C/���\��~���+_�2���Q�
�D����y��F���'��5�tn�%
}��VI��5���g���b>��g݀�z���{o�-+R��̛r�kIp��|o��n�_����;�DUп����2D~��Ϋ�u�;��Q?�w�Q�]
�����BN