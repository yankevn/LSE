��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۧwѸB�;Q�)�q�ǥ̥N�y�7x�S���1+��Aҏk�A�hg�S����	�㳰SC�����Ylj�;��Ɉ/yl�Xь�}G�X؊����;�'��VG^:0�y��F�	���D�:j�k̷��u��F'U��X��ù-�h��b`f����#0.� ���]!���豉��Q�HԞ�8of�D5!m��%am����Q�ݹ�u<��l!��@}2"�_�y�k�dì�}.3�槱�t4����$ǌ�4M7���a~�k���";d,�>߿ufj%qC�͐d%�̴�R[U]�s,��_����ȱ��`:�C��4�;��ё���5�щV�/�u�uvC��f抴��u�	_�߃G 宠+r�M��plֱe�A�v���`�˥I[��d��65���;`((��4�/dC�$	*�Fa	ֲH�ƦLea���]j����Ub����(���N��� =�p�s�<ƌ�;�n����n4�S1Pڱq�j�H�6���b���ٜz�����>8(]oQ�v��ϟ����4Μ��$�̑� nK�m��ɒ������	�j!x�L�}�����SL�����ѕ��Nc��K���!�꘣�~hyr����O��'�R����d��o�:�s_�/�\����KhxX�(3��+gެ��R|�r�Ǩ��z&e��� �b���*�YM����dM�,E�P���d1�$��������Zqg=���,���[L�3�Ii�}��m�����<���VAn&,�Q���t_9ߟ&x�C)!���{bn�|�9��7�-�E�i?`��q�R"���W1;�}5���Kj�1�I5SP���I��r��"*y������Jmq	��wS��")�ro(�`�P�"��!d���MBj�wlPa�M�qE hv�H&�<�o���aK��T�_���~����S��h�X�>���.�0�����L� 5�������:��&z�RƋ�T�ʆ��bdt�s@Т�� g���� Ǵ�b%�_ۙ[b�;	iU
����vZ�4��x���e�S�}J$�C�t����<������N�-�1�|ay M�R��+�"�Q}!~�� V�gA���|�3[���?e�\c5Ƥ߱�	���
� 0��*ˇ�B�!����\� +�}Y?�8��AM���"N��{uVBc	c&���4��Pa7+W�LW�%���"p2��a[�b�{�RW��Ĝ�^�m��qD��=���;Z&\P�.�D}�%q���z�&�n���ГG,��Yؒ�;�a`�$=�sZ5��npė���A/*��଀rj}�R[
�|�R��G�y�A]�J��S�6_���N"�I�>^���҄�J�I|��8O�,Ξ�C<��j��0]�h:VB'VW�i<�X1Z�ϛc�^W͹N!�Y�Lv`Qц�cس+y">�����ܯ�*�|��I�T�ͻw_����ἶ�1.�vEt����|���k'��`���~B&e~	N1S�Z�=�lܠ`�����L���?�(�w%m�G��*�C���#`��
�`Ư*�G�VXoy��OTj�wt�LX/�q�����h拹�?�f��@Et�:��?������W\S��$l:΋��Û��A���	$�^@��CHj*��t]Qe�
3]��: H4v��84L\�O'��'�I0Q)�����LƢ�z��Sm�*V���H6aR�[i��eˑg˖gJ�_����7�|�ROFz,cC+i_5�L��{��Ė-r� ��1�q��2~Λ�l!k�s�n_m��<���G��0꓃H�f�޻���U�P�d�C�����A.�b���Ғ�F�*���6�q����^Z\�u�b��l85bz,G�yBb��dk�O��yx��P�wu�*n"�����G����� (	0g7R�~,O��������.��Ap��%�3���R��]���԰���I�ԕE�tbl4D�j(��?�#��qfuҟj�E.ʣO����������z�[֧��nh�@�36�8Ύ0`2���焬2l%n~��>J-s����\�EӮ�&v|x�n[��:�(���@C~K�$Z����"�����e�(i�Aj���,��TqG�h
n5�:�Q��`�]C�{i�;al\E�u���v�x(8	o�#�#��k���sxn���dBv�Iq�����l���{�~t���2p�?�X��IS0���E�/���hB9�o��a�m���kb����_����(�z#���v.c�<�K�3����[��)+T��������R7*�u��9�j��;��m��05����Ԭ�c<�n�v��"$��e���ʪC< ��
���Iv(�a8ĥ��.=�xZONRc?�ɉ��ʱ�<����]@v#D�
�	ߦ��nW���F�aHѥ���\���̚����ǃ��HF��C���^�2�?��s0�!���
�[n{P�T����V}�OV�Q���8"�0/�����c'�����o{���^bz˪؇̓����*��[|ZN�6��b9�� ����f~1�ent�.ʀ褛�n�fou#ѡ*m@ �%��p�-2yj���8�`J�J�����f�^|�f�d1�4W�PC���D�sXv"v�/BR��K�7�F�4{��Zsq��m)t9�eŶ�8�Q�X���H
Z���)�`I��98����?��ߤ2�E��c��TѰ����p�+��c�Z����<ph��i��$�3g���)�)���B�� �%�
T� ��9\���5<N_��ė�P�S`�,J)��h�{���]mL"���݉��J��� +�ZM�8mB�mv�8�~��&*�@#x����& �{X��@X��P�HJ�N�hA�'�E��7/�gJ$��8C�6&M:��;��/.��R����)wD�pz=�!\ƻJ��5O_��7mG`��"��	>��Z��0>�M���q����i��0�C=u��譶ZJ-0�a�0���5���8�'���זC�}�Ӕ�yM��*���Po�$�|�Vƽ� k��3@���0�an�%Y.#��%�q�a��C^Xq�f
�s�!:+e3^�iO���J���RA�Ҝ���go�1NYKsv��)�?��Jk��d�b9M��� n��d9��E=A���/��׮X���!��8�U��K��=�}��q��D����6\�k5{�DSOS�T*}��a��6�{���)y a�-�C~�F�A���ܬK��D(^0���,S��3|�V��1R>R��^7�7ؙp��5;ǝP�)������"��J�[V�ż�PY��u�
�,N��c�]	J�؎E��Z��y;6и��Hw�n�$�8�2?�b1|\��:�+AJD�e����DYd��`ڱzG_C�k��` ��6j�4���N�<v�����z�Rɝ�c2C�H-c��rk��
2�3�T�j)u>���.��\	��M���=��S�ߗc����M�<RÓ-y>�ד�\�f���u�������2Wظa�
�mN?M����Q���V��)6����Kcp~%�X�@F������ᘪ�G�^K}�n� :� �!�`$���%9-�I�5Hfq�p��r%�m_��-�e9��Ȇ�	u�D�7$�<��H���)�+.n;��Yֳ��(��)�j��ޘRU!d1,�HP:�����������~	&y 7����6� ���A��h��Zy���� PC���6m'�]��[@�Ȣ�'�ry~�N����	M���1,��=��[�6yzksI�~/�U�5A(��T��I�����*�/Zb̀S�럞߂���u�=%[NAc��ыK!�%��[	P����SBy~���>BO�hP):�H����t
T��?��&Y�
��<�W��7@�{�[�I|� �]ı�ҫ�|߯�H�����!-��\�be�poDZ��+Aj�Ż�ܬ�F�,��S	ڹ�%T���7;�bTR/����^M㰋D�}��6l�ʤ��"Y]L0�3��w�y��Л�'6!m����+56[����g]>�"i��+A�-���I��P���B�r XZk��;j����eY�
K~!�6Z��O�k��l���"��ݞ�]�HZQ� �j�=G[;�.��^��o���25���hV���vZ�H�hAl��M�J�bJ�(+\��)�ϣ8?X��p��u��=]�B��PgӘ�o���H��h�,�eتk��@��͵~dq����#�Nƽ��")I�P@�Ҭ� >F��#�@��,�l��،��&�7Ls�?�9��:��R+_�I��V�5���/�Oϫ�9&��whtKy�5 ����"}��(������������ ������;���.��jo��|��n#�K#�����r`Z����<�0�NJpt�"�H�b)y��;o�	E3fM�=x�U� 6�ݎb�nO)&<���_�tAH 1�n�%��u�=x
Cb�� �~��"���X�w+�nFBj%F�1;���^�ve��ތ�r���u�W���]��ku�J�#�Ȩ�%��� ��o�Qlh�W�?"�3�f�(y���Ϫ'e���Q��U��0��2w�Ȳe��vZC����y�d��m\G6��.<��&��Q,�i����-f�o�y�gq��LE֍rY���lz�剝�B�#ՄE�V[����K�����?ɚѹ�Tv�;߰@�k��Xf���~��F���.ޙI��RëZb�o����;5�o�z�f�o���.��}�5*��]Iy$&�2���@ �F���.E�B)=M�2��ax��YH��u�-gٰ���I��#}8K��C��X~��3�$!p�pFKss�*�gF�f�5�M+o�|�����,.f�9ֈ�3
����֍��9	v F/sR�9�J
^�پ#J��B�G7�.g�`}LX���d���78	�/�:���:Vj�n�w4�i��E)�Z���c�n��Y�"o��Gd�/�F7�y[��O	�3���a���v/�2χ��	I�ͤ����	���+�@�`i�P��<��uU�i��sȹz�&s�T���'D>�&T�DM����)fók�b"\�����oO�aR��W�����<��ԯ	�"ж��?c��J*�����Bơ�x-��ԯ9���b�k��vvP��'�՛�4������o��h~����ae�1"����p@c)�S�\kX�	��r^%M���'�`��:��ݥf'q����������������:@���D���X�	o���Ѣ��A�6�y|�0��FhQ��i�71�0�k$����3}z�Z1��C�#�Jx�Vᮣr���s������3�bmW{��5���u�Fuy1�B�����@�1	o��I��x�1L�~کq倯"�[������v*���p��,T�Zݯ��\>8��qG���|Y�Q�9�dp �a��cd��3���
<�z��P}�b�z�_N�}$�Ti�����Z������4���pM�N%D�vϸ�M�Pɀ�������2{������Y�TN��В�R8ʐi:(��]1����]���uFu�i|�����S%�@d6�f���z�<�"!Rc��]C��V�����#[�� ���H�v��@�,��n�b&&ZV8w�35�xc. Hbt����7�<C����ٞ�A��cǥm�B�	D�A��d�j�������s%�s ��oP�T�*�0��C��j���E=���|��">��A���n[�S��C
+�z�/�r����j�� �S^�K��LCQi�h<�Ll��7�i���aptk���n�Gf�VN�d�J��� ,0�s�^Ck�7�E!�$s��Q�ܷ�L���(F3s��A>�k��4�y�o;�z��$%�Z���N],dx8�,��^To"��;�q�	��U��SQa
	�O�CWj��������c��Ũ��������
(�4��D�8����,2��0([k��I�|�>5�|[z�߬�68�����t%��&Ƒg�����y�X��«�~�Q|�1����n	_��8�,��`G;�H�T��t����o�m� L;�u�xk��e����<mN�A�`��a�{�N��cO�������W�H5Si��_�ǡ7FOAط�2*�ElMKB*h���7�]f!{:�8��8�8t �c
c� �x�gGrSg�^���ΐ ���7v�		3��5M���^�%�U����eCd0�U���C�w�6P���s�M�kO*E���"d�Y��oB1p�r�0�]���YO�J�h�N�)Ē�v�HL�QG	R�L_e%�܁q� �M_*�ŝ�FP�}f���y8-3Cdpe�ZG�׽l��	�W�L�)�W;��]Zx�����-��s�qtj�1�����~b�e��6�EA��9���I[�LW�)��hZ�l����*i�q7!�z�s��er�K�#���g��'#��)�){�<L(-6t�ߤ�'�+t��A������[�����0�h>@��1+�A�j��rX�*~)�$/�`�e���F��$���݅P܆�*�?��l V�Y�	I26��+T�=mfq��Ix�M��#����N�E��Z�+	 9���M�X���d�˿L4�R=�9C����r|P��ηL��L t޳�W�H�:z��bv,�c���@_���ߥ���s���ʙ��w����`kݻW��9�Tp�1g�]�l��c�D���7ϓ�S���+[u_�(���UT�6<Vۀw��[���L��?NC*v-f������?�?L�b~��?"��H�t�{��b��"���TV�Q;:uq���\���
�AE8�T�j�ݝ��%�>Z�B�@�W�o�)$���8<�ӯ���rAP��**G\��L&�C���e{��!�J��%Ϣ����cZ�ћ;�k��o�v�AC���0���ܣ=�sYCC*z�v����f�8؍��.���:v~��]��>6i�ʞz>d�PZY�*�LrJv������ݲN�ٍ@����X�퀑�'v(.-��z'���C��&�ck�r��7���E�1���-�I=�N�\���Tc?C���r�}K+ж,p_%�Hr!�� =������~!�f{�~S���1�9�ߢ!�L��Z���2M��?e�F�3k��p(�ʴ���h��9�^�fV�-��W7�vw�+��'-&�oF�	b�����e�{fbGg5>س�t���ީ(���e�Ɏ�(O�$�ec�e�����rD:�u�ɡV�ׄ�~8���yF�6n-�y�S�P���@���j:ʘ\���9mG!]��+3AQU��l'��>7l����A?B��R֟mS��HeO^��Y�r����{���V\�ޅ$�Z��??7�fL�A��ѴP��uJT�L�w���g�Ԅ�c|RW|:�]��aq���A�N�ڗ�)tz`S78�ݯ�._���g�I-'Q^%~�����}�x@����*�����<j$ʞo�Ƃ�ص� `��ӷx�OȠ4C`���6���a@§j=A� c����V~,�^J��"0f��)l��):�&�%�c�ۅ?[*ڽ��^� A��2������Caeg��A�\��0�_�����Ĳ�M�d.T\$H�׀�mw�W{F��V�}�r�#���J���d�_���TH�%U��?&��S��n�g{�2A�V>���0feJo���c���$� h���Nl]K�3!�;��n5�͑j��vC���lح�'�{��$wџ%���=uI*_�y�e������@�I�#~X	m�J�|{ �����
�D;���;a3�T1Ҙ�6��`D��e��Q��w��O��7s�󃷫�h�k����6��w��*�G��⭦I�[U��b����`5�H��E��Ƈ�n[�w:��BZv�(���G��C�)t����m�_��͏���:DI�Z�kyC;�ԑ��
��Q����Qs�;���a[kC�'��L�� ;l_�c�H�"s{5�ZD ����
?��Cva���o��`92ߣ�`j��w*=��N����]M26a���ܛ�t�BA�l���j_V^����7ʯR��K�]�} ��%�^�
�|Gn�w�ғK���{��e�K��!�ARdf�A��t�%������<YCXa��ѕZ`��a�o_�W:I[COY�p�M�Ț�`�8�+��#��H?:��g7��($N1�^��G����NK���MQ��G�y��v#�U���H��!���e���3��*^L&��7v�#T�6/����Z>1�)�\�b+{��Y��;�1������$�u�����z�y7,��0e�+I��¹�&r)ś�ȖTYU~�1fL�מ�꨿�������E� ��}�<�ŝ��ĩgk��awS�зG���\��0�f���MaEV�ڷ?�h���\����ԖI�����T�,x4�a#�B���wgiԗFć����
%��q�<MR0�fN�]���q��r�y{Qi����Y��jă��E�ʴc�+��3�~���<�0a5��C� �M2[�����P�$c!��o�k�q�˿'���BZ��R91`�>*C:	� ֝�%�,�x�4h��5U���T~���$�G��h�N�b!0�J�N�م8�7�{�����-d\�������Ǫ]
�^�2T����[=���ko� {l�j\L9$�kj�m�����r���c�X�����_p)�.\���R��+� �[$v��*P)]�93��̧������̟N?uy�
�m�G��(-x�M1�J�0�F��F�z���~��`��\8��삊SuE��2�2
�nG*���N�[��d��d3ZCF4v�i��P� �D��0n�0g�M�"=h�
��46���2�AJ�:6/Jk�y�-z��Z���#�˂<�N�Q�/N�W�(�#"Fq�� a)S��4�����dtUx��ћ��Ȍ�hڥa
��w��^��Ƅ���W	�B��
�'����^�3���e;�N�'�d+E����|�SYL_�&���Y{�.p?i� W�5�)�5 EHc���Q��@��~�g�Џb��K�$3Z����R��5_"��}_�jW�0�փm�C����vǋ4��kx�����Wz�If�ɾ���ϭ�.[��
+V3]Z���ء&���m���=�rG���S��Y��������:����{T�/#Gs�+�����u89r��-��$�����\s��ԌLZj�=Š{�eLg�N��`��k��-.w%��e��#zO����1�r���7�AhH�wJ���T��S�Xu�ۏ4s9�K�]�}�޶O�#����������l�T�F�)�f_�_��S���4~�׹w�@�C�{������8��d�B��6X�!^��������e�oe��9��w|?�ܵ�Gl<�v5�vCE.�O|ſ�c�1@H�-Fd�euJ��\��P�FߨM����}��02�����r2hC:!6�㸡 �����c`��J�ec�b�h�%wyٵ����g�]E��}]Tu��F�LU�Ȳ���F���\;|E���
��˂T ���qE����w�k�p)��"p��	�$'��wS��}Z�E6*�-�.�;�!�D$�Sыp:U4�~2��� L���u�V�vB��M�tA@�s��n�ufjHZ]���i�l���DG�FE��M,Σ�Di�je3���>�2�Ą��Ө������||x�m^iÉN�ä��ft81��?�V0E����n+�'�T�XeX)ߠ��д՘j2�21��0��]��_�?�=��,xw��8����x�>;��Ɠg���?�B����g �b���n�yN��-=�\mc�H�6�E�=�}���r���D+� ���6tf�V����xH�#{�r=9uc�-�~n���I��x�s�ӝZU�/γ���y����/����9Z�j�6�K�,�/����������:C+W�lr���\t�P��R������	�z.+r����4	f��24W4K&l���>�k��Xl���zYw�ƓE�{3��t� ��~"��cs��~�"iy;D���Qq�����׳��:�i8i.^"��G���j��x��M��n�����g��a�v��&s���K�2��t�2���j���5�#�[�;�sye�¿�>���+��>�\�-l��|�S^J-_-�����S��#[L�d���1�����ƶ���s˯֔��A����:�̙���rS#�V;�l3��MҪ��x6���� r�a����C�����	!��A=c6�*���}B�w�sB1C���cD��P�A[��#2~��!v�V��YrN�徙�oV����5>g0�ʁ��]&-&�.��ˇ�-�p�0�TC�<��L_x��%�y���q� ץ�J�`��nK~������[��紃����!�	��u��2'Q������C_�u<�nAu%�
6���&��蘒�RJ��c+��h2F�
O9f�AA�+z��qn*#8��