��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��^A�-�;Ӡ���U@j)z���|�9;@XMM�*E�`� �k9���:�Q�OI:�0�ǰ��y�Pd�ɉLb�vg�;��t\�n"
@�//�|�r��s�������R,վ`���Ydi����J@��ـKU�FZ�w�� ��q��ک�N��N���nAE�-���EJ�f�Y����X����v�^��� Fm�.=L�������n�da\��+��K>y��h�|�m1q������2K�6�&,�y��3��i��I<�!�Ȉ�]L4}��4r�RÂ9,{�wi���bt��/�����b�g&��IT �v��XV�2Y����Ѣ���y]�_.��R��G���A��I����ԍ_�e����ۤ\y�m�&h�	���"탯�������,P�D�Z���t/�F}7qB�$C�|M����R��.3��1��~�N4'sJk�1̵����5�ⴻjS��_��3� �i6"z:�I��2"�F�4��͇�e]����K�3�TQ.;�R����/��-��r(f
�uiAJ<4e�օa�W��v����AL[�EW���>s��y�T�~;A�2�Y��=i�>Z�R�_�	Y�H�1El3��*�=<S(*0���~ך����C��=�62z�><�^�Iî,�7_Gw�7H��U� Iҏ@Fa���|s3O�;�pK��������5������VaC���Gz�GB� 8[��%l����$]��"]�1�q�����9�Vh/�I�+U��)0���r��������r�6�NhD���S��A1�S���'X�r�	e
���\�%���|+�˂��VM��TA�z"<���� W�|�_?�cg��ii��(�h�~���^G8��uy[&"'�k�����K.["��w�zI�7�e�?�(��(�,���f��,%`-v�� ���i��<��2���38hg�v*q �(Z+�)癐�W\$�b���*��PՕ��Z2]����0�H4����S����'�f@-�$��D&��"����K7fo�����u��0p���Y�檎+��j����?�p7�,_�Ѯ��~{pI���}��	��{��t����(~����x�g�o��;�>d��U�;<LGH��x���O'^x8���G�kO�~ �\R���_�B�E6U����uG* Muw]�7'��]$���Z\����$��"��'�����I!�)�@�yKK9F6UkR#FƠ��W��35��G<��� 6�W4����3J�7�'�`>e�<�*�̹�@I(y�0���@+�|���a?,j~\�IR�4���h-��>RӸ�Wi�t�N����A���Q���o�;��Nѭ��90�p��A�q�������[���t��& l�K�1��2��8U��Vd�^cǸ�#&Ǫj����F+��ؾ��\L#�+i�lU7>A9_E�O�����`��|@=�(f�7���P��Q6{p�X�R�K"$/�:�y����#��df'ڹ"���Z�����8K����Tp��׽��iͅ���f)�<F������7˵�VHr0K>?�{�0_:����@R�l�~m`�<���1��0�ϳ�e��sX�UP)A�{�����u�#���d�!�]���TW��t+���O����F �1�đ�����sYd-a�+o�@��(�*�����%14�~����2�Q��D	5akbVN~,��6�B4l�`��Sߧy��2Εf�*[�>����M�|ZJ��qS��xc\��Qq{vK�4��� ���z��%S����c���W��4	H:�>8�5WeȔIX��ae���2�N�U�,D6���~��r?ͳ\�Q�oUb3���f�Ҕ�?j�¼�yd�yEkI��_m�7�Q]f�T(��� �y��&_�@�\i@�?BkX>#!@�~q�f�pѤ#�Luw!����v�R�sz���ρ����d19�����J�e\�P��'��+��#���(G�p+��㱯N���q��"�i��r_C#l�wF��Z�|j�ם��1��X��A�����,W
�*/l҇iζ�����?�dM�^�{���Ǆ��YJ'���.!�N����@�w��Y�;(��P���L
�y�HYT�q�"Y�6��`�^j�ueM�1��ҵj�e�P�n��3���9�Fj��h�yM!���$�83n��yq�>�1e�u�p7%aY���R�(�j��j�qz�/oW5o�=����,A��jL)㕲��>��#��p�I�e�>��WUr�����"ܣJ欌J�3�������/]LIN2Z(g��B7�8j�Q��䲦��C�!��{9BH8������$η�o[�ˎK�]-"��8(�:�Xf)s������F�t�I=�b���-�d��&�yž��b�q���#d�t���'�Y�݅	��]�YK����r�T�K�ltfAR� nz����دI#+�qt�a�s�t7�]#<�
A�ô�(L)� `��L�L��i{�Tyb˦Q�ܐ�*��>����R�v�b�z������4*��؁T��!%8�g F�3?�����Oz:��ʤwR���Y-����ʦ�mk5���4u)��8�@p�|� ����)v�&DҎ���(���	`�>O��RI3� z끒A�ղ;$��|r�\Wơ��#Bq������]E�+v�⼷U�? ڄ~݅����R�h�xC�nA�{��[��O�a����1�V��8�O���W��xc�Ũ̀��2�{�uQ��u6�)톳�����HQ%-?��dv�@�O9�T.�>����dbO����������>�)�t�v��6/�%@<�S��OV;�K�,t�{r�v�6���E} .� ��%��m�{����zjH$iJyL`Q���Al�Xو���o�xY�9�@����!B������
&V�z��0���8�X@����LQ�b@�{�kQ��吣�/ļ]�¢�TH���>Si�*m~���7�a�y4"G��>;d�r���lj'm�i�hCԡ%
XD�r���j�%����t׀��
Ls��2����Y��7���jX4�)��op����p��ݔ���5銕W�'IX~��u]�8?�Ҫ,`�Z��8��l��yк㷭q������+�2�KB��9/����@ޝ�l�E�gÜQA�.�><V�)���� *���ۍoS/�2�d�T���Ko�IDF��2�_��vk;���@$�g>�HZ���+�6CJe�s�%��du�0#I�{=�ෑܠ~�D��R@T�KMm]}��F�����I�Ab��qf�hzw{��B��9�/�~=���@��-�I~��������-���Mp���'Yg8�������L�wȺ�a�!�|�}�J� <�˚BE��t5Ǖ�]x`��1�|jT��ۼV��T�l擔{-��Y��z��٠�"qk�Lm�즋 �1�(;�����&��l5���_�j���s߮X+��B8p���v�a�+� ��<�D����|p�s"8@O���6v����b+e�����;(W����{ݒ��7���A!���t~8P�����{�<[�
rɡ�Y_���t.рGS��NLKsO����oY@Op�(�������D_��~��9<wO��d�]�l��
R��s��26�v�I;���o~����W�s7ܦ��[����trQ���=в�Q����K����>ߥ�Axg��7&�6`�a�CG�6C�g��s��d��5~���T�;���n�
`z|�&���wn 3�`y��:�RP A���s?��/�T��7�hFyt����2Br�0��ÓoO��q<}wy�2��
:�S kw������-"hc#�bNJ�`�c��{��%$QqɤT
�Tݢ�Ty�T�hə���qK��Y�3U���#-Sʺ'���7� ��+iW��1`躗6,V���5/G��E�7�"����̭�ʶ"U��S�.L��2���-��,��r	������.gv���~nfjsD���8'�k�o�A+��p9^��㠄24Yٶ{)�K���Iz�!�_!^�B�.�@w^���_�0�������#�dێ�㻈&�WQA�=�6�\��޷g�JQ��r��s�T�>併_��Y�Q���Փe�	��㼃9����>
�s�k3\1��E�8��*�t/�X�!�\O�W��?����V���[.�)4T�
m�E�����dH��.5'axduJu�L����6G�& ��u����d��I����ū)͕��4�'S^�џx��	�ǹ��I��~�����f���}Nwd�?M�xP�W��ɐ�O���<�ۡ�����\8�b�xf|!)��0�,�c	Z"�$��1)�p��B��S�;G��f�\/$a�{Xf��7}����y�C\��e���f<)BR F8��}]�X��@DHbt���Y��b��K�Ax��m8D�_�\08�j����k9���G�����kE�wX����a������������1`#��J}Sl������Rɯf�G<L>�
�\R�3�,jWn���홣����oݙT�Y��ZW��cU� ��xj~�
�R��G\֒q�|�)a�0�bU�S�ǲ7�^3�s�	�-��=v��]ʞlmĦz�.�Ҏ5(�}������Y���	��ة˦�Qc��_t���R�CӅ��!8j��'Fz���SF;�����'D���l�h�ZB���I�؜ �+�9���� ̜�����P��'�0�=�Р|hC?=�|��d׊�U�r��v
�$"?I��@o���{��؜Y�Bt����q����s�R'��c
��6�g�[$���V,�Q��Q��+c�I�԰�=H���$��mN�2�-?�$�׹���G�ݢ�� � �Af�����"Np�́g�cj_�~���c:��5\�7�_ᯤ����2�s�*0H�{�D@[��e/��upF}f�� C��Ƭ�L�s�+T��{�A<jV]�F�+���9���'x��U�1�U/��.�����C�02�I�e)��%XW��!|Z������,dTX��=͠>��|#��)�$Zu�u0Gq�	�t&x],� ��:�|�\|Z�%����S�.HC�lŝ�ū�ͭ�C{�F���T����c� �,�
��j����P�IR͙�����%u�c͛Bq 首Y#�
<o�W���ZQ��� ���Ж�p���ΟS0ՀC�@�w��#���U���.G~U��N�_#��72�c>ύц�	^���^3�­*zݫ����
�+��l�/A����)�=wu1ʨ�6C��d����9�|���oc���'v��������]6����7�fPiަS�	�]��򟬭���0�0h��uG`<�ć��9]�� ��6�r�YܳA��_�ɽ�r�'�������;@1[g�³�%m	 �w9j[��',e/����ߋ*R?v;��=��E�� ��-�+�_	wUU������!��j�*�~8�[��5����Q8����$�̞q	ruZ�D3�d����\� �%�D�:[f�'n}�� )��^�h͞�z5!�d��I�[S ��<��#n6UZ�[B�/���Nu�G�����2�j���B��u㠊Y_�����ZE�t������&����K�u���m�D~����SHm�ĵ�f����|d�?{�r����2k����TM:�����Z\Aa#���X�RE��l��E��p�I�qU/-0��C�jl�%u�|>Y[?%Wo� if�>�Ͱ��+�7�����^��#���k��x�C�L�h�PLAu}���˥6�E�>��`Ae�1W�TǮ�?:�����.3q�G����|�q�+pC�兽K��bFKC���;E�ڜ�s�ԃ�J��G�� 7��B{�����m0�Z�Q�ӻ�k,��m2.%����i6��j�|�����|���
��
�W��s��*�M#kg�bK���`��.�;#Ǭ������ �;�2]����m����8_d��4��ϥ�1�	%QK=y�(�]��v�z �/�xd-���Z/�B�U:@��'GF��^���V�d��v�+�vlWH��-y&xx��ڏ�%�h���$q3���`�9�P�`R�+�5�K/�D���MQ���]|m�n����U�N���mH��uc`�}�-#}�421�gHͨt�qH����u����r�dʛ��G��ju�m�	� �
����qͪ2}��8I�Tw��Rg��F��a^��Hߟ���@^3Y�??��ئZg��֬i^�#>/��#�����Kǃ(�Q���,�훱��|�����P_��=s�|,~@�ZR!��e�\R,�S;��ѕ��F�I#q�F{�a9�p�+E	a���P^.��l9_��#E:ZI��b,\�I�#�`,�W�"g����0��͓��G"9�jXݏ�H�okť2� w~%��|p��{X�?Qc[�i�C�tE_�G� ���h���Q�?����f����{��W+Z8�40I�]
l�,�fM<���iw0X]j�����'T����m	�:�Ub�U����	eh����/b(zSs�ՠ�_Q-2q����{��{s�1^Dz Ki�u�i��6@�.5���i*��a-��	��-�O�i�4��"o���.��A|�)�����>�]S�֣�o�Lv�6,��n��2Y	����a���IZ@Ӗ�h��el�A�\�89���hl YTV��ƨ�����C��|��%v���Ӄ�`�5���R����4�_&��	�R@!q�s���Ȼ%c���T9�U�,ҀT�9� �x�M���<߶�l��>m�o(�IJ�As�D���f�up;��uT�y̚�b���y����oY$��;��g�p{��9��3C���l]"ے�*�����Ua��i�놾���ˀ9u����	3 oG��1u��bͅ'�y$�F��]|J�$E*�;��³��^k�5hy�n��cG-I!���^\zuS��W�^�w��D�BobpIG���
�J{������wԦ��&a�P��qP������A�'�`?zY�	*k���G��9�}�ڠ� ]S�C�(�/�3�(ShJ�k�Cx"3H��U|�H��2�H��l9�������0LD�J��W1�"��Ͳ�F��\6@���<���B,� �ǰC��z6`{0d�:2U�J�*�פ,r]}�}?)�q?��2���fh֖4l�${��PZ:ٷ1����+T�����^����NH,`��㰛O��q)���J鱐��&F6(���ͽO������������c������/U�F� �x��^3/)Bu5�r�wDq�)����,\�_'բ9�[h���&T(Y�A�(� re��3����Ң �C~��ZE�������Һ��(��-�_xX���o,Tb"�v�4�f�7�zϏD1�*n/�O�7�%,L��"�/��Vx����=�9E?�~1�I��ol�Q��_�)�4�Đ�j˫m�<q2N��"�
�m��&u@d�jJ����<(��W�F�������g�V��;5=>��+�8�Ǿ���۩Y� �����(�8�&u�Lԧ���ߢK���}a`�~dì����|WA�K1e���V<(�ح;�;	�ܫ��]�wvJ��^J�>to�%20�N`m%��F5U�:�?璇&l-$�&12��a����C����xd�,��A�l��O՗&Lֱ���k����蒂u�\)�@�we����EX�p]h�E���;a;�snG"�/��q�@����8N ��$��]W=Eh&G��^��.?���q2Uh������:��D�KE�jf���:~03���I,,�`����f�3w�7��K����s�;���M�$�
mڢ����Q�@\s��g��F�`I��fi��O��h�x�	ە}y<�Q��(��z��Te:��%�8��R�-5����"�ow[�E�7���4��y�����L����2��R��(�NG�O��?IB�yV�c�tm��Ɇ:#K�S����/j������wyΤkEz�%�<%7���އ�ؒ�a� ��1	��+\�3@�T_oU��#O�*t�>�wfb��y��s��� ���;٥گ�S�O��C��-ƶGB�<��/��mf�⡲���Ea�Cn��h��@:P�.5�*��8�Xڥn�!*��	���)]-��4���s����@I0�f`��[��ìS��&P�/O7�_/�m�V�!99������G�;3;0.�`�<�JF���PN3�-�0d�M�bt���l_�a������@�������ڣ�Ĵ��ܩϷN�6�y�6nc�˔`���jX{�;Em!�0j��^��z �����k>�4A�v�Q{:�癅��8���iE��f�d��luʒ0�����6J�)c�
��Ǌ$9ipTSsa:���BYц�fj��y�}�p�c���Cw�eZtr�W%x@���j�T�=%�,�)\<.�����؝�Vf��=d4<����+��O_�'}�R��y|S�R7��*�}�Ŀ�-q���'�9���SԶ�U�T���x�ĆY6�
�:�y�vH� ���k�EݵP�-��K ̽��s8��B ?��Ӳ\�m_�:�#2{��U����G�������e?u�738�#8����&_^R��|��,�u=t��SN��MPw��!��2d(p�����x���a��2�V�
���[����e`�|I'�J���o�������>66�r�T�4��U�Gdp�+�Cqw�m�#�Pp)���n�;?G�~�H��p,�Y�g͜(r� ;^�I��z�<��6����)~�,�$vI��6�2�@ �`�b@M@�?��v+,�iҁ;և��`N��aF��1A�H�Z�I��x�^�_�k�3;��2�8�AjN4�����EĤ'G����:�qS��z��v��K���s�.V�����3�����=��ߦ����{�M�Z.��)�f�S)ŐmEvu޳�O���:*��L�ҐjU$�m�����}с�0q�Y�	���[��a��'�0����h��<[�;����Ak��ͪ����pX;�5��)LCr��G��j�	�� ���)^�K� �m��������IW��!����a��.6 T&��L����C�Q�aGk�CTN r�j��jA���t������[ܹ�1����҆~t�L�K̂�����3؁��b�\�1W�bJ�2%�5�0)��]�c�^��>w��B��M�̹�4�8(�����QG�3K=��7���$�sIu�2G�8�М����j���������Kn�Z����S$O~w�-��~_o�vUA�K�s�+�$�9����N��rY/K�c5�ى�e�Ί�o�\|�e��N�C	���E��3��z��1����m��ڛ������"��ۺS2�z�)�<���-���%���oV������y�Zp�%�w ��M��%�դ8��U��WZ����Q�Ј�3T�.)�o(�OW0>P���<v���Y�D�f�����ER�;�5QdU&��M����uE7pם`��ˁ˚`�1)h���i��a�p�!a]ei$~�;�0�Y�~w�5�q0O��,7���G"Ǩ�iګ��{�����CO+�\t���B���S$dW�[����J ́PeCs W�(�I�Œ��Q���6E�;J�n�=r���0u��{>٫������}���B�[���3Cc�Ž��r��5��B�b`o+�?�ۋ<K����T�8V9T]Tz1a���0���z��X���T:�?�����nm�C���F�y��a,�.T6<�&�k�,18�L�{�]l�>>�(l�P)��?�m��j�<z��D<:������ͦGbCb��?{;�!/��e[�F����d���68d�\�D����ٮW��
�#nP��곇�PH���.~&���(����^���U��q�������Wf^�6SIaM�Jم
u����������Q���z�6-�����6K�y�rk}f=\�oyd�����8RY��W������u����>T�'ߚ�9�e9�^T�UJ��>p�9��4C�8�)��"	��U�΋�
Y=�������a0}�J~H�ja3�����Z�
h�����7�|u]�����z�i(����b�čkF��*�����k۔d���#��������s^QX�8�1莊zI��+�5��I���ѳ��q��lJ�z��ܣ���bD�@̶���Q���j�z�r�G6�T�Ձe�xE��֌.�Cj���ٔ.��[��Kg߬�'JwiS�wS��;�.l�_q��ǦuQp��B���<l��`㮰�����.=�d:�:_Y��'t�������`X`ތ��}�:",e?z���a�n��Fn�2�������-Pf`yFߒ5�ҴpA�z�e�����P�_��E���%BS���.O��Y�d�Ɨ�X�'��{��29<W߆H.�t��<x�p��0]�%eU���M�n��+b���Ȯ�5mĻ9^Mm�P}!��T�uP�4� �S�ض���S�HT���[���6n�L�F>�h�~B�{���n���	#`y��$�F�{��d�~����"k(Q�Y��?S �C���]���AW.M���䴄fԌgc���r�}��m�@�
L�<�������ݮB0����.���Qس��>E��ôO �~�*�&׳=�aob��C��>�Z�\y�=����9��ĆTSgn=�>M������Dת�xJL�T����)�.��nk?�����<���Z�-~�-f���M��d�S ���s�*�5qy^$_���&�}�H2	X�z6*��!nO��H�c������)2☐Û��)+��`:p֩y��b��^\�$:s�#L�����#u��f����c��g�.�u!�J�<��f:��b�����t���Ck~��{4��E!���X�ͨ'i�&UI�8`֪y�	`��@s�驘ށI�O���-!+��_�&z{��Nn�U= ��3R����y���6��r��.d�>�(]�t���E̛�w��ft�@���~!�~F�u�vV�2�ԙ4ي�W��nz9��eEw�ץ���ޔ�R�����^E-(Utb�8̇�qU0�o*�~�NX�Y1s������@^mqdX�W��݊����E������d���/�1��Z��_�$��vXSa �}�~C�_'��-ݥ�/�Vz�sO#������']��oB��:��3*S���{ș?��>H{.��\��q�:~ÔNr�if~�o���X� `ȖN�g-0(rk��-�Po���/�����
�ܪ�@�� ���Nؾ�g��j�y!�f%��T�j��:�����i��#T,�23�r�@�x��\_�lhdi�BY�ҧV�N9�O�ߐͺo���#|N�ϝ�=Զ�!�_�TN��W|@ՒZe��"v��jA�N�WK�M%gk�h~r�G��G.�r����,?��%����6��Pi���
��y��;����XI�/�A��]1���
�o}��y$�d-w�r`�
�,�,���u�'����%��,h]J	�N�����ƺL���]���ܼ�	u���@��o�8H���["&�R��Ф��d.�T������g݃΍�@th�R�|��f1���I��D�7f�X��X	�1���������2nV�' �^/���qS0n�K��'��ʛnhP�A�)V�����0-�\/}����2_�Qdx���ݽ�0Ƶ�>�͠\G�;���H=,+�n���2U^ئM��^�ɽW���ĠzJ�3Gr���G�1xV�f�Ԝ��ƻ6T�9IR_%�2�R����~�0z'�	����ĵ���N)�ź��:���^M�H�1B���Un�@d�m�)w���+,a�-L��i�A2��<�|:���,9���iD���a�:���"�4m͍���&#�p� o����W�����(l���X{�&��$�$B1v�n�,=� *�S4~��-]�}C�R�$���$kosG��O�*//U�>�T�h��c�q/6�K�G5.͎}Guj�O�1ǱA��A�V�si��FV�c��&��6_����jWPu,��O�>a�3A�����@���Nr ��a�:\���lx�����F�]	�2C{1d�;	EΚ(��@�w\��j�T�Pہ���Jg"�+e� q6�E �������u�u�S�e�-7ٸ��n`3���,b������r ���GX��Ad�	MdA�>}WE���%�)�o����O�j�DL�bir�{-$��d�cUxu���^���x�_h�=qVl��~t�[�bQڏ�/��	zY�+��w�'�����:F�h���sЧ�	U@�WjZ���� �ts~o�>��jH��QٺhM�U�:v�K��f<��Y<��va�C2���ć]4j˓�Φ��7��a�8QX�����������ئ���3��C�4y��;���~#U�J�g�(�.���K��.�Y��[�l#cQ��Ԥ�Sqv�y������]SCτL�F̓{�d�W6�Ҭ�n˺<
a�Ͻ������P���E�'�=l�?g٬Z����9��<~O{j�f��`�r��P�O�UA�'z#QK�P�J_�E������'�Іr���ӭ��T���H%�رu�Jp��fsk�W\�>/|pl�c�X����M�H�����T7`�>��_���4�V^�&S*o&�~6���jS�D��Xu���0��H�|9����i�C5n�@��C��o]v�TX�oҌ��S���x�[[���:�7(MC҂ì� ���H:�1�;7�
�.�!A�r�8X	�[����gMf���?z\�:Pf�9�O43
�E�Z�,ct}��5\19�$���/��'��p�+�۟XO�'�="��dfF��"I�
A��l���d��9x$���
����)�3���q�'��kʈG;���Ѫ���A��U+�U�}B�5sy��C�*�ws�
޶�K�?a��<~���$��CG�-W�l�G�k���)��jj�V�M۰�Q�<U�iB�=�#�,E��*�$�F&���u^1���& ۄO�}\(�_|	E���Q�6ϼ���E'0j����i�]ӴC���n}${��eU����o�}�<�F��������t�����y�I����8��o,%ΡT����h�˓��͠�������C�x��!��j.�j"=�����e�V��Z8U`�z��jAg��[������"Q���˗%����<R�-ʦ��2Zk���v,A*i	o���ݤO��"��O�j� ��^^`�Xt�P�%#e��>��Y�b�ԃ42�z����p��ʑ�q�o,<͐�*G	���
B�E��W>��K]7��H�y��3�0T��1��Yfh Y�+���pS��x'�V�>[�x:�F�̶@�݊ҽ��.Ν��
sV�����䰸n�ī�2]?8���=:Ͳڨ��0��iW�w�Ԡ,>l�M�O�<��أ��G���#���k@	ZR���t���Hb�Yzn��TCP5N�U�=�>H�����Rg���#K�4u�����>�}�4��V��&�)�X���	�q/u�W���_��3[!�����w8j�쎁ݸx���
�W|r�e��G>\�+y��0[K�����)�b�z��m{U��	Y�֯ء��4�p�r�U�d5��~���FɊ�ّ��J���k�b6ZN/:�GC?�]ݨ|��(�X�ZP�"}�Ō�b���@߃x��o"�8�u�дu(fjʱk����˶����
������d9i6�e�ղ%o{�~���ɳ�l�`�I#{*�������v� �!�x�T;��n�u��aԟ���JJ���]2#X���aEQ��M���j���UO���b�-��A�ψ�z,��ִh̸����XGaU�~��3Sm��.Z�!�2��=`��q�����k]>*7ھ��4�p[�dT�|.,�&V��'�Ygv�Uس��V�xrY���ӑ�ϫ�����W%�3�-+�U�w����Ԃ�[���Tr�Ý�\lC:�Zm�%O��N�!.c>���U��s������n*���Vb���)iܙ���ixo���Jp:�ey�Fad�Fp]\��K��_�ʡp�C�!�Z_g�O3�4S��!���'��v~��m�A��E�M4�g���,%�����Fd!�q���	r&=�eC!>�E�V�L��[����W��h�^�nca�����T9��UF������3�1�N�h,Y!؝����p�#s}��s��}�(�U�j�-���%R�9�.f�_|09ۊ��m'�
NH7�w�ƹ��=`̀l�Ha�[�=J�7@:�f��_��j_�v&�|(��h�(#>�V�;��� _S{��6u�~y���=:ʦ]ӥ:?�������j!z%=<_"��h��)2����g����������y([�Z����YDy�|��Qo���x�&m�)=�+ݺ���a�I���\�B+�p"(�ٍ�J���w�1�hJ���*�����աԨe��+����̄c�[8c����Q�#|���A,G���6�-]��<�@O�|Rp���q}b�ZV�[R�K�����w�v�oT FK���m���s�l<��"��x�\��P�0��ܤ�$V��U�9�dٯw���թ&D�0_��횅w}�f��?2C�ummiouI' ��'^�Co���b�$
�2�}�E����v���ؤ��z�;Z�u�P����e��n�����3�t����Y"��69T�RJy��9��(�^�wE݄���}Tj�BK[>B�־�y�v�7�LP��<T�tM�k��U�8��/$3��U�i�{�o�e�I�J�D�"'�ȅxNZ�o7r�\r�FE0�_�#Y�'���+���^\u� �ÛN�4SW{�8��z����������*��Ƌ�l������𤇢,��<�@�z]R��U�^M�c�#c�!��UAreV2�
����Н����O���+3�ә��E��Z�Kt�_3L�$�ns�G�O����`���zQ
 G�z[@H����#��I	f����;������i���q��e�.p�M���5��KD@��&Tz{�6�Ȇ[J��3r�`����}T��#K\��^w�����;*��Uw�`�R���X����|F2�u�HvMʁ��"
�q8�A��^�OG�����o�G��+xo��?�S�H�Ҧ�Y��y�=-8ʀ.���HJe�7��O��m��T۰}��� ��׋	�,���_�09ACRWV!O1���+���hԷx_? �^��BP���5	�&U�6�
N\%v6�}����cA���İ(=��4-%�I�_�~�*C��#���6�@S��3�W򴣮�?��]�S�n_׏g��UC_�xW0�Z�"����RK�zy`K !L��j�/z2��*BۍD%�C�Ol#��� A�N�T~_���	�S(�(�Oq�"�T!}_�&�N$ݽ`b��S_�]�W�p3ꐅt$�h�t�b��e�(5��LX�҉����ک3(D�M̛�U�j�1���?�b9#O�u5�]���a\��m.u �۴�.�p̼ �i313(8�z_����S�W�(���/��R���^G&^0�Ͻ(� S���hŞ&HQϱ8ΫK/�b0t�c͍�I���[T
C)7��4�Bv�Dn�=Jv���ZU"�fr@�l�����I�;	U�͟��+A��߻�s�C� ��Kz�1��8VK��$���^"l�1G
�A�ȔR���C[Ӧ�l^���1�3%���$9��J��=��P�^sfi���>����րbjV�����y
%w�
�R��!��]�&C���ۀ2 ����������zz8"t�����'by�^�<2���%�u�,�_t�]��p�+b������X=�a�7XFIZ�B��=Т�t ����iH��?s������ɼUuM#�)T��tPP*_�Y/6�Ǩ���7�K̆pn���pj�X^��"�|��(?��3R�L>`R2���>�YQ\��\3B�N�D��/���Ն��u�Y��+�Z��t���~⸁��0R	p
V�Z;�O�|r�)�$�;�	�?+�.�o�(�-�z`�斪�et�2EQ��ƆHr�Y젿�{0�A��Z!%8{����B�N�i2#��MZ�;�y��\�H�P�T+J3�/z�dg�iz��Z�c����Y�'ʙ���A��>������!,v���«�h����c�>���ҳz<�����C�/Z����N0�����+��s�b)��v��l��W��m:M�Bg`��vk�P^�����`�G ?�&j{@m�Y�ZQ>��z��V���-�6Y;I��o~۾����H��=_ԋ��~�/NҪ'|:ç9�Խ��faƜӸ�
Sө�m��ӿ��f��Q����a�Z���'�b��Rp^ �̓�$�os��X����~ Cٞ
֌�-�~�:qp�>�-D�6:���Ts��r��T�FmDeA`�53��w�Aw���WW������]�vRU�n�$�S^1��|�[ɔ莲uw"����h7�R�O�q��,��E��c��/q���h�T?ø���F�d^�3�EJr?�}�\�oM%�B]��'�M��Z��}�ޚ7���HJ"K�]HZf�LȀ��e�R��l�p��t��:l��S��5 E��e�*qV-�2�+�ڜ¡ϭSr���Q����U�i�i�T�Xo&��Cn]�iZ��{��� ^3��娾3������.�K{7���i�����Uo\-^��da���JZ�ۗz����b��Ե��"��j���\T�,U�V ()$�W#Y�z��\H��Ƣ���0�߀��R0t������Ǯ��Ie9�w6U����YX�:�|�&�ɹ1I�+J�f�|�	J�+����[�Gi�
�d?ͽ�nQ�&,�X�a�сG�q�_��x���B0~�⦉td5�G��v��!����k�6�-8����_�)'柁Aƚ�4�ˍ��w�i��L����$��]��Z�"�F��k��H�Xn!�c�w�sė�n�5��$ɉGDI��g�D��Դ�VP��
Vn�9-X����|q�'��Ɋ�b��R%kro�ba�TT��|������?�z:+�U�IrvF=�hVx�]k�:�AEO�I'䖂Aň�����dC������T�o�H*" |� ���{c�6��W]�%%�<ku�X�	�O��"�ʶ�:����"����љ��ن4s/�u��z�~�BN���t=y�a3�'�a�iÚ��ÝL��ifl���q>���X���@ν%�����~�C��3Q���<e���i��*�����8�e>���>jI
�+J�dp�`89�t{N7�Vs�)=H��ޠ��^!��q�d��Ox��?:����L�	�j�}��kti۸�w���5�,��:����̠me���h���
�@�՘o�|�n����(o�~f���y��G��]�Z��&���=�K+�4 �??�N[L��d�@r��FQ��9Ro����;�L�n���˗�>}Lx���OieΜ	[�
�1^��d9),X�+�`4�|*�E��W�Ɵe�d�3^kB�����i@c��Q��̐��o˭$/$��d{�b6h���
�x߮��Rn��1��ܓ�D�	�+B:�<E�������<�ֵGo ��Mv����v�wo��S�5��3|�y�FI�_�Fx�]O��Ԧ0𾒥��/��P�q�q'�{i�j��K���{���Sт]��
9!"|��	�	� �*',�Ag�Sy����X�����`a�eX� ��b΅~�=��%'T[C���c�xO��ͭB����i�\�v�:��vPv�1���KDF��A��n��է��Ê�9[XL�|I��!�� #�Q`C�Q9:�MF�Cک�l��������#\C�����*8�}�ˮxOI7rʇL2�y�Q`G6�Q�)�$�SU���#�rqb��+�yA�Z�k��TJ	���
^Iq��J�ϓ��V�ԺT
E�ps�%� P���ڬ`�|<��	~��4L��Ԛ��`(��'~���<Q��15��?	��N��Slո�Na���}�x���d�,. �%��q7.m�?S�]ãj*�82h(���4ʒ����p�ܧY�4���9|���<��X��N?���������A�U"�n��� 7<��N�Ě�loj�ۊ\�ڵ�b<@[v�0�E��4�S�6U�9�j"C	ؽ�v�x`�ҝl�@�3U4�[�:)U�lh��z�+\��K��~/D��v��z�����Y��
�+<��z��Z���'�j��G1ft���@Kc	���w^W�[h�]�Iͳ�lyMS]SO���4��YBȄ�=�t*���*߫���C5�Sj� ��że�:��h�k�\��^����x��~��,��BN�+���t��y~%�����.�a�П��{YR��Ę|�/P�?��=uMh�`�@��&�ReQ�xy�������ƥ���'�ͽ�����Sy`�\��̩�{�cɭ	R0% ������sر
j�#�o�S�xQ�d����^0�BT�ѝ?����WY���i�r�2T	.�w��8D)x+��a1I4[euV,.5�͕���L�/o����,�������n��$��g��vu 㬇 ���P��|���T/Y�wi��Su�\��C
m��c6J��Ơ}u*�/ppe��-�����䋨(�b�C|����dj�����2S^^R�3&;�
�'E-�ƌmq�.Z~���?�XL�@�..qOy�
MI�,�ތL$��Hd�_�:=��U��e���c
d�ԝ"�-�wM����tO=�m�ۮʣx�T]��g������L�s�{�M��9ͧ��!Ns13��6�)����JT��K\��h�h���v��w�$��ŗ�����2s��P�6$�p ��M��X�͚>�kp���k�v3Z�~�=��p��������������\�B��S�n���x��N=j[�O�cE&í���37�����$�k�y�楰��������\�"�>�ה�٦��yAa���b�D�
<�;
i
M�ig�w�MW�i�ʵժk��8FT �4�� �@/��Z{�<�Ë�=ZU�.�x�������P�]q�+�|��ž՘ʖ˨����?�1��+�?X��ah��MP�(����+�^��[߻��t�Lz$��5i[�_��-�0o���&c`���9�!(�S�y'u�l�������f�)s��
G�*N�� ����c�n��[��C&U�F�)'��F�Qcz��7U������!�7�f�?ڗ^�(�E+a#�a���pE<�#�"��X���AO����.s��.a��\M]������D&���R�9����Ȟx�$]�74���-�@����5���8[�Mo���1	$lB��p�7 �ەVss��fa��6����	�u�B��6o�fso���D�<�x����.�q�X��N2�������e�>�FM.��Wg���ʆ��$�"�*���Qᷪ��s����f�ǿ=���M�*��^�gZ@l@\����	^رW����]��u]�?�*�Ѱ��h��M��QH���<)!�!M�f���-�������&դ�(���mR��d"=&Nvc�O�u�]ɾ����`���^Dm7�ϼ���O����{�$�?@M�ag�\�W���ܱ���.�x9���&j��p��J.{���|���JЦ�PF�me����E���k���j�K��=2,�8#�h�;@쌕��7�����U�g�+e}`�n]��U���X��^��4� u�4=�PЬ�=�3h���$��AW*�]�i6��c�AU�l+����U�W9my��`�(����N2���"	�;���?�"�s[_����{�đ�uy�:w=�8�D�*������7mB_Ѯ:��&���9���G�d�Yt�zRxn&����=�Yv��Hj�͊���K�כ��'`%O���m���}���OmUFFz����1����]�DŁ�'����q��S��?�MQ�P��5�c�E�	�p&ވj�F�+���i���Bv��_���o�V����+OXɿe����Lk#�=_;3��+�?R��gO�܊�мO�Uj�	2�|���1�p$E ,<���Eg<W�+�G��9�>n� �</ qY�2�(	�Rdx1��1����]`��G����u� b2Z����,0�Cx3��~������<�+��uc�B[fZa/�IP^3RխF\K'�dQn��.�vv�K��ω��0(sdF�y�#H���M�ڍ3ZK%��	�
�+X��1�����I�Qh��U������
��w���ld �s���{��.l�.��PA\��42gl�,�9������Jc6��U��t=Ӥ��6��"G�ږ���\�~������w����:�g��ł z1��i�l��	�*������	m������O~]�\��D�f�f���i��r��'�6�6���XN��d �d�Ϗ���j4��]	�p{�5��W�T�w*���w��G{��Q�|*���s#��,:F	����x����I3�u�Y<P�I��{�KY�� -�ĝ�N�mf��/����l��Z60�U�{Ç�?���OZ���/~¶w�9X���6�~�y�v���;G_�aU5[����w\����B�������Ũ��0����eO/�������e�p�j���<�0�P0Y�	��#w\mm��b-YB����Ox�T����D]_1j�Xf�7�}�+MI�>t��ٺT�R������c����S��q+9�ӫA�| �/���A�n88nAU�S����wQ�Y������3����0�����
�gx�[B�&�
~}L��`�U2o�rZei�,���Z���G�-�ݍ��)�{ELow�u�B��8�'��a�y�7�\-��R"��Y��K�M&1�ix��S�h��\���ձ$�
�{�疪Tv��{f�%	�-�������]]�;��sk/�31<e""7_�!o'ŃT9ɶ�)0QP��$-�ZH��WGI+��-�'�u�(���~�Q���e���,��V�z�D���S*G:���S�$A�~��r�����g�m��B+Ჺ-Ƿ��O`?n,��$�(�Y���o��2�iW*�cP��E�D;&���$��UL�TK��0y���Rg����p"C߂�%�y���#������xe�|��A�d���\��)�S�i���M&�`�	�*�W�[�y�ζjZ����v�S�;���߶�`�����ӽ%o.�a�C���s��C�����SW`=��ZP#(&�i��2�;ǷDL5�
��e}I<� U	J��u)�%T�����(p�q�s��W�$�Z�.j�k_B�v"���ڰO
�x�K,�8����)�t���{`>�y��� �|gu���K൲�g-f6�㫹)b��I};¥��8�%�j�U69�v����N	�;{`pySu�����ok���P<�>ǡ���GfT��'�؊{x±Fqz~����f�}x����8���9 
-�=m���W��ꂄZCd�P�suj➝���z�R��Bq`S��B �b����%^��D����.�l�pЗg�o-K�{�!��Ҥ��.���'ɖ&��������mݐx�̀�)�;������kNrP�`1����Q�v��v�A1s��S�7��ӽYy�j��@T�2�Q1�O���x��=�JcDr��h��Uv����z4�J���SRJ?o� �$̈�u*���=gp�����E�N���3�u{�զ���~
�s�Sv@��S�̆nbQ��TV�����˿����W;� V���_�)�7��P��%��^��B�Y\ $�4�,����/�F�b� ��Z�DC(�c!�B�V$8�դ gN:N���̃��Կ ���Q��)m���ğw��_b�|O�[Qv������]�s0.t�~a��b-��S�Fu=�#U=����_�F����WT:c��U^ �<�f��P�g1�z�y$�<�=���iY�)I��ZБU�S�䥬����9�zE�&Y{먥���1���U�r������R���fEp�J�� �ps@�Қd�Y���uXS��/N���xM���Me�<%�a7F�4��nG7{�j�Kf/]�X w�0�>t^�b-߽m*��KtbWb��V͒:�L�'����MF� ���w��3��CX��Ni��,�?��SR�µA:%q�t�T�4}�<�.}ˢ�=*�%b�����f��Y���ZeR^yhR�m�'zTj�|@���^��'���t�H�]�����I�#UUM6�H�1����˖q���ܛ�uT"|`���s��M�PwQ+{�e��<�e^�r:|�&B���
��Okd3�+����Bj4N���k�)U7���]��O��"y%��%�Ue&��b�h�X�£��yS������s���ni0�J�h��E��pi�L�i��S뜻�/OY�%��1r9�}�	�]S?����$��D�zFW\��0t	(T�����>����qa5P4.D�Z���Q8�s���m?�~w�U�����T^�(�:���VP�+��������K��ܐ/�8�aaQ��l�S�2>��?r�`�!�B���i��-4.��ȑi2�ꕒ�Q��~q���r,���Β�P�Y���z��:F�ʡ�<z�����lX�۳^�����E���Gy�5	�� ��O��L|��+���-�o�A���2�[�d�j����xa�؆�f�x����o���^�W'ǉ�hnY�{�Wt���=qgS�����⿃7���j�)%i��9V*�k$�_
0_g�J���g����hЏ��2H�e��$��O��|^`����Gh���ڤ$x&���F��"C�����Tb�����ҥuפ��*)_���g<ז��N�s`Իn��
��xoq��,���<k��gq���}'�fd8!j!���qj���^S{�#ՊA�����1�w2σE�Ut�j���k��6���LЮ$���!�M��i�v�X��1	�s��2��r��^^�Z�J#q�0�r�K(eP��� ,���ȅ�N�4 ٸ�M^^�毡&0��5��U9�p����6�ĥ7�"��e�lIL�^h��b{<�*��W����C3�(��l!�Oߣ���[�є�׊gܓ�#�6�QZ�߾�ѱ�܉Id��Ր�(m��x�z�"*{���$!��;�K8�t��v����!��r�Dq��*�K�$��X��
]%Ӡ����3��S�H �oè�0+�\P_��DB���w7��%T�z^�H��7؍T"[W�3a�� I�4"��P`�=��ˍ�U�gM6U�y�ľ�����c1?k?3,�1X�lqrEZ��~8��̈́���u�K�6����/�蝄
� GG�HNp",��=���	r<���vB����.���S��{L�݁o�X��X'ft39�&+#�>&��/W���骳��h&����`�ܕ\�V��dW��E���4CX%5xDvۻc�PJ��m���}Jig>l�f�Bp�Pk3��o�pW�UOH��QA�M��}{RU��S~6�S�o���걮����x\�@�{dF4r��l�Zš`d�)j�y��7u��jL}Q�e��m��sH:�)%1 ֢�>��� �r1�J�c/��a�/��z>ߞ̹��+-;h ��*�m<���Mq�ٝ���~h3P��(�l�Q����_E�qi69�pE��(�����>Ş�d�܊��nw�[�$���退�1M�R"U~n^}R�Q��5��ne�!33]�Aߗ�p�ka�x���r�*X��SAh{\Bo���?s1s��C�k?}N��V�V���c�H/�B"��M?d\�^[��?�^���X����Xkؙ�@þ����2��:�0Y�_qfiS�">H:P�s0��-nrě37��ɜG��r�8�������oD3��\4p4
D�r���?ɼ�=���5G"(a�uw�m罹����$�y�}	nMp83���b�V��z�p���F�EwC����}*�g̸��N�qi ���;0���9ٿ'����ʍ�xN!Cׅs�.d��,��k��,���;�6�`.n�Dh����N��cH�o�T{�<uӭs1S��=Y��'�����f)7q�Du_g.2_ ��u����I�6��b���?���qZ?��Vp�Ǭ.@S�ؖ%鏫&��_\"�
Ԕ ����E�m�ը��؆���O�4�Ʊl
�W�&?RU�.�JX$���Uj{Wi�v2�z��V	���������h���?q}����a�eH�x��~v����2�����9��X�"X��g궞�)���'_,��l%M=8V_�9�	��
+%M�R>~��9�@V�%���R�ؐo���q:M�N��'�U�&�S��ឳ��Җ^lZ�[yc\f����X#Xĵ�Ȝ2��9�|7��L�R����-�Iq��YA�	AS�_N|m�a��-��L�nѧ���r?�XbQI��:V�J,gA�ގ���Yـiz)�ݩ�EX�`�`@�4B���_����W��t��"�*Qm��Խ�#����)�\�r��sr�J��J�K�$�M��E�����!LLp������fX
8��M�;]~�
�]�Y�}�]����}�r���#<vr���[�A���W�QJSzn�R{����A~������E�`��p��qeF?%���n�@�i%uÑ՞D���f�K$�Q�y��b]���O�����^����`�ya�\�x���_����_�.�t���(98��1�Æm�ԛ�)��
M)/kޝ;���ur&�$��n��<U��#::p�.@4���A����Ȣ�،��×V`^���LNe!�i'�������M�JMK�$G׏õ�P�&6n��*���mG�(��$C���t�f���]�[��Bj�1>�WX��mD�|�Òw��в��~�żib����2+��β��c(H�1A����y��[ﶵ�R&������^s]̱��0����$�*h)���1���@��&�C��s(��"o�(��Z�cY�^�NO���i�yw�$�b�'���OB��|�����!�Ms���[��Ր����4��J,�1;ǀDZ�W�yM+cN���~�H{���`����ft�?����3��P�d��^�f[��	]G�Ų_�pP����?���HS�E�O�}!^"E�O������6�IݣC׼�����v��`�K4e�6yk>!£A|�ύ���J�����L�.��-2��Zsk?$���A�4�(#�Dj�S��,V��8O�M�XJ+�w�(��j�!+�7ӫ<U1C��fR�����8�^i��?F���3��6�pFtmp ���0
ą��BENSNk7�T����|1]�ܔ�m�^m"���Qi�'VUѝ��P�he�H�P�6�,)���ץ�[~~x<�&�NڥV��D^��<��$�aM�N��&;;�Y�r@0����x7QN�}��;��K����Ŀ<^�!*3�m��O���q�@5���,(�$���pP��u(���y0>��k(B�����M��$~vX¸����t���z��J�
E8�۵uv����u�q����w7�B���2�m�FP�������D��~�,7�;���+�]�����Y��j5��CZ��˾Ƃ2Q��N��j�Xԟ��J�@�l�a�1g�'�W/`�.�_!iz�J�"Rؽ(�l�%��e/s�M�v�
�Or)�n<yB��PWҖ���m5��s�3�>C��o#.z���b��UCir|�׃N��t�{�I�ZV|H�(��N��7L|��߿9P%^U���:Q� !�A��X!|y�~I|�f%���?�+ƚP�`&7�4p
g���B��U�<�K8^0{W�'9�y|6A��!����7�ؼ�j[6���ww.k���sF-��#h�in^m���\k�����r���W]��|HY�:ۯ/J���ё8�*�p���Y���|t�:�
! u�!:Z�,ɿz,��(���r��0���:z�t �R��r\�:�X:n ��9X�-���w٤��"�Z!��@y^���3J����C<�6GQ5�=�Fj�b}斎Lɶ}ӭ�@��WS	6�݋�q��0$m���SO�JИ�5F�#"�R�"�o0!i��+C�����PQ垢�w(�Ϻ-�Jm �,6?]ӻ�T�^�ww�@�%�s(��$�Q��(�։޺90(��?� ]_��?''n����0�k�/�x-��\mI/��6�sGȄ�3{���ؖ������^�EI��fڸ���(UP��p^N�y2P�@H ;�|���yHy��� :�u��5�oq*h��]�h�û}.;���2������ٰ���?w��쬷��%G}�����dBc�|<�H���9��-�`q\=:��ͯ>Y7k���ս�DUWg���gB8�=&���;3�!�H))��\S@�TѢ�lN���Թh$;�����Q���\{��m���0X�q����P��W>��u���mri4t�@8���6����O�{8W���wp�7�;ᷟ�A�y���y�`Q��AcF�-ctD��j&���Yq�N��#���qM�����	.�N��"	ЩM�����rj��)�.@�hMf%��9%rK����*��Y�HJ���6�vOJ�ɑ���_P�5nwb�+��d�>����?!�\'�P�s�B�|>�N�I#9�V�Y�R�8 �K��դ7��I:�9������yi˗��>�6���p2��:��Q�I���� ��d%���y�+�!.Q/������P-������`�# ��)�D�{�~�aq��Y�w��x���l�h�/ƚ���_�0�/���#��	��<�>!��� OiTh��oH�z�IP��6jZQA�;'���Yv��b���9!��s���dÓ=��J�vTtfZ���Ö�p�$v���D���#���t��@,��_�ڵ�.1{��A�+_=�-��滛U���{�p��9Hpv��Q�nD�L�$���9Q���Jg�L�-�[Z�꠽ً��otYd� �y����,[���mH�6ap�XH��v|>�;�'��b��FØ��؉����7�j��~��1p���0�A�uH�^b�ܤr�:2���H��|΅�y<�5�\��4����&ӼVp�&y'=wƚ����N���^ ��1k.�pG_�f('�*�L}*�$��7�����Q��K�߽���5荁}3���Z�ۖ�����qF+���;,�a�5�����;���g�`~�XzGc<���.Y�^֙
�$V�_' ���&��H�?��m���^�%��i�+:X oN-
mX�d�/�I�oi��@��]J�;ҾQ�@����Z�	,��1�g�2n˾���
Z��1B�q S��6��b~���0å�Hf ��/���۬Q�z�)%�',.-x^���-����h�w�5L�~�у��S��JQv�k}"T�i���T+��^��zQ�ԡEO^�����tp��j���k�cHI���Y���� {�v�OG�,��i��<*=�Z�'�έz��?�}�o��&*�{��D�'�㊃5��D�}��G"
��)�$Ez�<q���)�p�6��	_^�S���ǭ��<n^��B�}�:�@u
�X��$���S6���,ƨݢ��w{�ղǶ�	��cΜ^t}�.g���� r��y5���C��H\3���z1U5�u�K������=�`jg���C�����Q�,�	(ʸ)�#@��S�Jl?���3l� =\��Y�c��9�0����]ń��.��#f�z�gagޕ% ��u�:��;�r���,�1�w᭧"&︂�B�m�fSep5��T�{�Iu6�Q=���_NG��wxE!��� ��4�;U̡�.�Z�zr�*����6ꋧ4E�<j�.ʔ�Q�S��
*1"k�Uf��>=��y5�_zLgg/+;k9.��w�x��OH}��c�����T��F�[}Z�y�h�L{,�Aw�)n4@!�"�o�t�)�E(��'/��sB\����^J���+*�)��4�K�^���{2םb��N��	�^"��J�8�9ބ�ks���?��D`�1��7�V斷*���̥N���4�G������S}��ĳb�k\�j����7��P�Y�	��(/�ɥ� �7m&��	��Xb-6 i2���]!wc�6�0<]�$�ľ�{�ūs��]�O�L�W:�ߨ�g:DZr��}�βT<�r�O�:|��N?��یA�'d�#N���O6�Sew���X	>tx1=9j�j:�u����y-ӏ� ��n^������V�0<�!��	k)3 ��i�+E��S�0��	���H`cjf�e���afN:�1�����B�>8	�u��>�w�9����\u��O�	qPoK,��F��oV9���_���o�D�E\5������g3z�>ݲF-�s�=�8�j|��{�ӛ�DiWA��b�+N�5l\�b��_i��p��^�mbCr�IUֈpKC7Ny�k��r�Ԁ��j��s���g��(_��0�t�� M�00ݩ��fH�/�&Er~!'�����u���WH����n�dAy0�?��N�Cx%/��Z�a��jТ�6ŉT�Υ�b�時� \?�pԀGv�ѿS�X�U�yp�����y��	�\P���|�_�jK�K6��]�[��=��n J�ݒOa���&[��y��sW?��y垓XC�Q�l�YD0�bwb�I������LE�F�n�!�w����>�#;��S���`���(�v&�Dc�\��`n�xi�aĠ�k�/��=r�S�|��u3��P�)��Z�}���)�,�y��b�x���Ϫ�ۼ-�rZU�k\�f_�M�6���qq�f)�Xep���Fsg�1֦k������lF�?�8p���@�'��t4������1l�P�7N�t���tB�	���	���#87���:o�;�1jk�\inIȟ	�)ܶ�Pp��ᚪ�&8�Y�۾�p�f��M�y�OB�r����aY�K��9)(	F�cb��9v7�(�0%ԖN
�{�����==#�n��`���_'�� `�HL�$�!C�~�FM۫9�[�ɶ�T�0TN�G�TM�JzX�r�1���L����.�lϯ9X�:2����H�B׭	@�?�r��BЗ.�6;� }'���{``]V8�'�J�"�;	U\T��D�fMhJ��$�T� I�B��I�����6pd���Rz9�ߵq���u��]Ƒ2]�S��s:��͋x+�J�{�o�%��EL�/ �-����+�mD��jBɵL��cD�|����m�yێ�/G"&Lb��^^��no*(Yu��U�Bl-�����/g��Z �M���Z����eX?�_~;n�I���P�H��1�n�O��X��9.vgq� �����,�����M���޳x}�Pm��2��Y�z�op�-y�+�`���ŉρ������\ˍ.�^�d�7�ڲ�2Ά�f��J�h���q�b�;6���[��o����+H��b�m��Q��	��?B[/�E�n�>[��p�K�������(���]�]-_e�����v+.����8����%v(��TȔ}��}*_��qb(0.�us�I������`���h���|v^|(X;,<4�&tS���~��C�!����e�hd-���a;������HJ#%���6�a�K�K4ͳBe��r��-ns��WB��l���6�+��p�K>��0���t0��0֌m5��ԙ,C���$j<�gi�2t��=ax����E�OvpD�5Rcd4wv� ���&�iF"��Ƨ��I�f	�� �J/
(,N���H�KP��¦�5Xa�PH��*�fp˷}��.��I��E/)��w䵇��ٍ�Z^Ʉ�C��^¦��Ɯ�B+n�W����Ɠu��Kv]�I�?�J9'"="�X���ĸxB�K&���w�)YC�X�%�sI�q�����$@otk�
"g3�w)fq��Nr����ȔX4:�a!��wY���>�>�k��Qd�s�@;E�P�7�B<pr`���6�r
�3��cq*�O���u1*Fa�2�x�(���II[��ڦ����:��z�E�z\b����Z��(�=Su �����G���`��?�3�<# c���uŠ0qXO����w�R�M�9�>��E��+����F8Z!��L�] ��p��4v��>��KI��8��I�]�,
ݱ�)]�w]����H�#慽`�wٹ����j�b��4g:��c�K��t,��Ei�yy�!^q��Z�ٗ�Ѥsx��%��z=�h�@��h�f���1/J=����0�Н�%��Ļ^-ӹt$��,~��̲��Ѧ \�b|G��̼Y+S@�/��}���:�㤋����M\�0Q��l�Hw�T�SMCh�4�q�M��dFX�|?��c����M���J�p�� 5����ew�|�&��8��@��UJ�~�:��
�]�T�#i��L���> 	q+�����Ғʁ;=~�c��a-eR}�[bV������xNʉgt�hi^�ձC�#S�&2�)�;��K<nD��D��et%�|�T��7I!r~���ؿ*�Q	Z����V�ί��p�m�<�Y���@�$c˻��ȱ�<M�� ��>$w������d�0�\\���Ф�	��^��ѕ村[C�&W��b�9,���m'g��ǫx��.O�*F����@������I�?�bI���̟Z@_A����\����LC���g|[���;�`�t���׋�
�r�T�k{�Cr��J�!_[#���Ѻ��@�Λj������˟�����!U�������4�/�dG��p%r���>)4��v���'���1Rh̠�*��W�EU�#�V�� 9(����Y��ͥ�9,�c��2�sA����%�/��,��=�,��n�3�?L�_İ��W�&G̊��z�9־uW&��@M1��������m��5s��蓂_�$GɣP���<p �E�3�Ag�_�]�[|]ر��iL^����m��8��I^�D�zX����+�[F�uE·a^"	�`��ِ�jSV����� �� %s�ZCY�Z��46U���w1�0���'�Ԭ��ic�nd��s��7��m�[g9"6��.���2�Q�p�}';�-�Yzk+X{��i8���g����kV��[FXP~h�'��js��s�>����K�#�"`/h�5�8g;Ĕ��R����K�-��8�,ٕ����:_K�v6��I�(�
b�wMޮR~�6�@��a��~-2C��|�M��-��Y|��	�<j�0����#u#��	Ga�Ꮳ��*Bo<5H���AHl]�S��9~���k�����s���8mϾ����(,տj!΀c&�zd�zɺ�٦���s>ìO��8'�.�s~�K,��,� ��TEԁ�@ ���tSI1C�K�Y��8� (n�i�j$Z&��B+� P��NŦ[����-o��4��+��z쀧\})?�ݬ�^��i�
y[ޜ^v���Q��}Q�@fh�"��T˳M��n�b�X�3�lS�`x��7�pf7�)Vb��a����F?qm��։��)bѾ��eb,���������e$��b��t����
�,������?38r�6y��Ƶ'�F����2vk���f���s�����XɻUXs2�C}�n9R�+4�0�Ly��T���ܽ4�y��<&�4!Kؗf�	f<X� �iȹN��h��I�S���2`\2S;~/|��iw}���UMX+r��B#����R(&z6r1O�#ܹp\�F��aP�2/��(+on
�L9:�tDbnF{�勤��_�8cYW� ���Z��i��Ѩ��{�
�)f^��ޅ��2�yJ5hz�3|��n$��M趧ql&�Y�
�{�ĝ
$�1nԫV�H�&m�4���k�b���83���]�Z�f�g������8p����-��F��G�<Z�i����;�!pS���j�ٵQ��¤�\	�� �5�ZҰ��Wh��m��V�u�.,���J?��t�JRj�9�AY���a�in���)���`�!�.���G�j��w�@�*�DI�L�S���^2�1ɑ!]H��7ƙpX>���+�L��E���:��S�Q1��V:������%pT��CUcB���s*�y��ʘ�AߗH�y/�� ~�kz7[�������e�:��C�
3���Lѡ�w�@�v4[��7���޾�U?\�x�xwޞ�/�.��,?sǧb.<����=�MX����&�J�[��i��F��bk����:ǿ^��
OU�ۻ�U���Ε�}���h�X�	�����'5���ř#��c=f�z�| �!d����)Kie�3�F�P�|#�tVb����y ����^6)-��Ne���j���d�y�]fkQչ��aj����z�a��X�wvoڧ3��ntz���p�x�Gk@"OQ����s���-R��z�覭��� 	U@{�bJI��	A)͵AL�G��>��R'���<0��2v=w��K�P:Ш4�
Ǒ�k[��E%N�B!�ag��T�n\P�ݟ�F��c�W�)͈*��Q�%�hř] � �w|�æH�m��5c�\�N�"�4pD�_G����H_	������u�2��/&�Qp�C�1�u�g[+�@2������p�.�����T):&�"!*@Q�����Q7t�Ė7�{�1�d�x%4�a��We�w ,��96�c�~�9llFQ�'� 6~߹���czL�Gw�>ۉ�\�5�.R>X{ù$c�QX���'��
N�#|G��pZ�7�f�%�O�?��9�^	W�-k5�:��z���q�	�ͥ�Jy�2�B葳�*���k� �oU���a��p�as�K+`T�� ��ge�k�bh�)�% �Z�����F͡w����7x�mm���2��򯌦����
��޿m��)��2������N�d�N1��@�9J�z�S�$D7Jh\r�D.�8��J.����vv��:妕p����g`W��~cL��H��dq��-�b|�ܪ�^r
�&�?����:��v~�e�,w�j���-8�B0�kd�K����d�����&j��`��%:�7@�a��`�%����	��C%9�ȈȗI�3T����\D�͒��������NT�x�n_M�Oh{� ���9���
�eɋ]�:"��!��c֓�ǉ�r�N����gp���Ij�ȘT�՝@#|�t������'X �|�;�HE+�y�@���\�o�٢"�<D��W��������WDk�j���~��(�;>�Ef+����a��&�k�ٳ4����7.͕�<K���V�W�2�P�1�����|�9�Z*4f���e�>:L�f���8Ġ��?�&��OQ=<wd�k�Y*.	�kƃ,"��������`)̎w����X��|7��΋����2����+=='�_#�)Ф���l�& c�fU&(�,�A�~R�?���i�ް;�����?a���h�(���钼=O�c+�`�#�|��+���#�����b��O�#�]�0V�ԝs���ʫ������%4Z��e���8g��w��bÍ�M�i�9y��R�5�xt:��p�����d)}�au�}7s������ia*k��9<'���H�~u�=�y�!/<�
�ؖ����T��Ĩ9��\�e�p�'I�t�ݷQ������;%U��8J8���M�������W^Y�g¸/OZsB|=(�w��x��_��{u+f�n�'��%����例(��~��ǵ=�!�⮉�8+W�?��'����C�,�n�ԡ1Ӗ�� :\|�I��gY��a�A�AT�C�+��z�T�ɛ�����4�򶃬q����)j3t�˦�0��O���vϩ�ڪ}���s)*t��O����oVH���P��ޙI�h!x�l��� (��fT���14xEc'��������gn��>�����M���_u#��,&1 ��'�����6ݮvB6?!����~ڦ�
���m$��a��D�ax8�cPk��i���ߕU�ꎪ����Z��{D0�g����� %��d�I�Oz��X���{����8���G��@�+Ӿ�yC���b伭+F�\f;�ȴ��<P�E�)��ַ���C�?��ZWm�W�Ui�ߝ�����T}��rܚL�=���m��� �ƃm1M��$�z/\��ڿp8���j�5JY(%Z�A�M���/87�,x���O���K����*[K�G�Ct`��[���2����;$����D3�R���|(�;)D��'�u5��if~�C�@L�D�Qn�ʅ�B�|OC����6f<oc���Fx:H{����|�s��c ��f�C�S��.R)��~QnO]��&���]/�v��72qG����j �v;�P�Є�
�|C��sf�Hg�%�u��E��
�,���^����1��@��Ѣ�`
ze�����:Ұ�^xu�K��f�*�vɼ"�h�F���f�R��4�>���^�}�絍/85u�WI��
>lthϬ�%��kW��*���x�#�#%`����i�7G�0���ݑ|�������yQ}$���Q�R�5�@����d.�,$��d���
4�UM�:P��\��7g��6uxu����|��Ʃ\��y,����?m�zqLW�k{d�:��h�#�u�
�A
TʓGu��4��8�z�/w5#S��H# R뉪�(9Ub���u��|��?�K-��1���Y�z���VN\Y�No�$�4��n%RG�{��}��������L@Ny�N�Y�GW����P�Z�`����C�*^	f��e��.I'�_OAzƜ�Q�VIp"���;�K:���X �����"�\�\n5״j�5 �"	]��Il�!�\�u%���ê��䃇qc��g��B�����C�"��ƍ�'�����%�����_8�+��A��3����{�;	��"��gd��_���<��֧��>��]t\�j�q�I:W����͏4 x��10Q������p�aV�-�(;��z��m�ئ(�
�L)�ц_:�Z��^9ǉ�8�z��8�V��4]Y���}ubPp�/��4e哹(3���%d��nQ��= &�7��=�S�����'����E)s /_��W�u��]�AQZ�7�h�buX��}y�K��k�w2iMV��״5����Ƒ��G���B�<��Xm�)��%k*v&��-�Oo�e�Xv��e��;M�|(�+�8#{�ɴ�jr�[��UE��(�����%0�G&V���{D$��[����j�j���`zG	�:>���l`*���.�k�@l�[.�={���Jx1�wL�K��$vm�V�� �Ǉ�6��q�}o&n�mc�Q�X��Ԣǂ;������Es��l�t�0�q����y6�M��e��tfd�����}c
���G~�T��nX�aS�X�Q>4�	u⦸��q/���ݸ4�ߌ��:���f7�T%J�k�B
|ͅ���J�Y9�^#��r�$��O��yn�KA�>!A҈AvQ�b>ί��q�bYoKx��^��o�����N0B?�6�A�	��G�d�A!�-�#��ew�O[{��W�^:A��ɯ��8�^�(oqTk��;��U7YMG�wQ+"yq�=_ (2��$ۚ���ؐ���G�����G�A�� �����4Sȸ��|Y�n>ֹ۱��9�;���ol��*�HjP�>�t �������}d��?�/pC���z��Q�<��gLu��Ur~�"{8���"��g��4�!�V�{F~D���L�yz$�-�k~�T�����!���"���TE"$��JF7���C�L��A�
* ��w��@�ǵ�_|�䃨v$�np�n���jcXϷ�Vσ��˥!P���c�q:^c$��cP�'�'slYؠ��!�f~��K^B�,��a��N�঩��i�?�Ԁ~a�
W�����EdF{�LQ��B�O��*��`� "�3F!
+4�/��(˂Mk��@
=x�Ѻ����VˑO��N�M��J�N�qo&�a�SB�6�`�7(s�-s
G.�e�Y	}�1*a2�'�{�H|�Ϫ&����R[�XLG��i���w��z�X%���n�!F��7�l�x6�R�ؚ�5�ɍV�R��Z�`�]-�ǖ�?5;'"�x�R:��m��xk�&����Ö��Z�a�O� V� ���1�bSav����3�Q!�D��I�o�Sb��bJ#B�Fh����Ϙ5���8H����#�
�%ak'�bɰ|@]F1�����6>�5���t{�8`l13��K�����N�u��:=���Ok]B6�R%��7�ű�A^��	|������H��+љ���4`_�o���R-�V@�#�=�hXC-���:&Q�Vu��.s{a�fm�mX�����������f����؜_��"�����Y��w��X����Q�GU�ܹ�)���;�M�Ѓ*��>�z|i����U	�v��2!�٣z��^#.G"����jѝ�e��@��Ve's�l��x<�1�Jfx�j��ʳ+)0��@�֮(��x���F�>C� \W��܉i��p�(IV���)k!�=f$a��Ӂ��;,lM��O +�	�APCx���lJX�4۾G�82�K��wL3��X��e �3q�8�(33�Դ��&)���dG5w���x�m���z���螜�*��/��;��rl��U�_�I�K������`��VԳTvN8�=�������2�:�KR�=�es�S���i:RY�-�,$O/<�b
�w7mҎ��R����^v�
x~�d�yM��-��a�Lf=��d����K-8p��NL�ܰ�Q�`ؕ���i��I��F�ң�&ޟב��7�:�ƒ,җ�����m� �cb�A��l,♙S�g)0p[s��B_���P��L�%ɕ,�7���Fd�xr�X����91|�Ⱦ)�=�T�
%�ш
�]"\�AHZ�yi��gt�$ya�5���D���yM�t7Mg���6D�&��x|�c�c����^b�	Ka٬%�����S���l%�M�F�����	X���E��K���$�k~�о������k�X?Z�v��w�>�90�c:Y�{���Y'����s�:F]^;҆M�[ �*sR����������V"`O� i�:�x���V9�|X��u��e�@n�W�!��r,3M ��v���WFX�*cp1
݌����Ȏ�Fi*f)�́c�s�f�����R��.3t��8��]F!����:
C'+�t���*�~a��(�V�c��k���`��q�k7�ć{K���S�?��6O�=44țL���8JL8}�����z6�a�l��Ԫw�^-�U���l��%z�	��4ۗˈ�y�O �9V�O&�A��׽7��%`26��ӹ�*���ܮ2n�&.��2d�<Z�!J��`d�ӏȥ�_�~��5l~=yO$��b
ƞھ�CF�~�@li2�Хi������SVVL>�za@G���,\ Ps
����S��5סN��U��\�E�v #�\/�py,Q��
�G���;�������������5��2F�B�BR|�l�}�M����'�I���B��} �*J��m�D��	�h��"]0����Z���gngx�u^�R�e��©�:b�z_y����ܬ�zy�F=wf�5ot.�4�9�ɍ4��.�}, �dz�������pQVs"�jxz4_BPK��R8��#�V�5p9�y��1�捍t�,���6O�-�g�5,V,@��-p�<|��y�Z�j_|�O��Щ\�Z����Bf� >�����_.�W��P*S ���D<vIɝ�cvT�×�� ��?4-�H:�%DU���DP�]#vhChr|�'>������R>"R�`���qߊ��vSʿI�-�d��̏��NGW����=
���R�V���0����&Ѩ@���ro?�%�w�8�V���HS��������v��n��Q�]�Z2�?P��T�H��ܟ�|�����Nw��r'�s5���Gm՛���,Q�A¿��+��ʖ����C��n9�=U�-����3���?�-��i�Kc��DL��	�l�qB�y�#��+H �T�O�������.��͐��#�e��P��v��:��9��� z.^�l)��d~�: �&����[l� 8���7Q�1I�g:ԁ���eSC^�^�������z�QWu��Iʊ�an�����WeWI=��U2Al�k�Z5�ݍE��y����?[5�E����\H�-��<�[��ӐtI\�T�qW��p�n,������W	����L����~�4H�:Px�$bxF��jg��	X�����_�k�W��/݉��9��\&{E�����8�>l֨~l� �D�g��'�&O۷Y��:���"�ˮ���#�H��׀D�t �6��~\|� ǥ�G#r�ۖ�.n|�R�>Ɩ�Ǵ��v���F�^m��1���v]8�#�%�Iv4X#��g&7�J{0D0ȴ���q[��Ӽ��_o$����%��M�g���bh�vT�	D�'�^��T�s���@<��?�V1��M���x	�4p�}�SQ������r���4�\�TM�Y[_��$�⒔���|��)%4Ş1�Բ���i��v>H��H�Ûjw1�s�虽�$n��⯫@�&�j�Y*|�IՎ��0�T�^�"�5-~[usa�94E<P�kV4ƪ�Fn�����`�L3�c���l�F�-h!)U�l�o��#�'���1�>���l�����Ս�,�--�NZ��T洯�9_ ��S�4�X݊�Qk`�$]�,��Kmd|�`�&4����q؃�4l���\��
��Z�U7��LV�7Z�(ϟP�$\xZ�k�5o؊���<���z����[_���:Tg�g:6�c��Ţ�Mf#`�GVy�R "��AM�Μgv��ݸ�
أv��������y @�g`�lI��� �G�G�F�����T�����A�����������a����V�!��ɺj�$:�	@�$O�� ��0K}��)�*@�����C�ʸf��b�&w����:�qe�n��|
858�c�E���Ҭ����Hi�@���y���74[�n7�Yy3;��y����A�)f�?-b멠f�q��9T6_F�D��B"]|}?W'��D�6���׌����\?�+�I|Kf�����_�R�TƧpo_�����c����ŧGmCʀ_���e�(�)'d��?y̱��i���6��,�E
�Uu����/����F���¬�Y��'D1(�OoW�D��s��Ԧ�tr5�لr"6��@�w\�>�n����O�W�@h�?<r�&����>�\��K����8�\?e�	���%8��V\h�q���6Vg�o�� �1$рrR��$�!{�7�A!���kX��!�^K1��0�r����$0�����x�2.b����'Nɹۥ���a��*dq�����w}�&l��n�%��r�O����IP �݉����#���ЎXֆ����g+�LG�ۿ;\�X�W��'���<a����J-Ez��5�,'q9!+�[�9�L ]���#�S��E��E\�^�擀cJ��?��_��Z�	׬�*�h��]G" �pM	�*�`�9.,�\'��ACj@B]�q8�3^���T��>�+
b�G����7���G��jp��s�Yޔ��H b������L9����	]:zn�\܉�Wu��]*a������[��%Vd"0o��PV���mA��ؕ�-6��S?G5�;Kub�[ms�'�,}TSC�4�,�r�%�MZ�M+����гw��f~���(N�����$��hP�&d9�7�?�����4�����8����'懸k�27B�%��Y�c�s�Txσ��F��k���F���/�4