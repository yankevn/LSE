��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ�Bq���F����9��	X�\|(�-��:j��ۏ�,���$��,�Y
��c��9r�?�1���\G��L�T���|Q�CN�0���cJ�H.��3`�H�:sz�+�+�:	r9r+AY�[����9'�|�]�wy�WX6>���S��:O�0��fӭ��ҍ֞���gUbo�����`"�jyᛁ����Qy�J�k� a�q^���;��u|���܃Dq�� t��֨P�����<w?%X��̮T�\��i�n#�3̓g�`DcP��J�*M�*R̺	�+',C#�ڎ�>Pm����gE�Zқ84ud��Z��LmQ_+�f��sW��|�7��rX�\J�'q���v)-�0�t��Z|~3����~$���}����,�\IW'����X`��#�l�bJ�h�U�MͽӟVӎ6�Jg\��y���3��`t5w��?.�����~�Q�D�Oϭ�x�fZ;{��ǔ�J�	���;e�e����e���X���m�p�H�<�-�OBo)�<�P�X�m��ט��}�ƃ�V� ���k{������:΍�Ɗv`_�pQ���?K�z9�\��N�����p�_R��F��X�>DZ���B�{�7<ȁ�F��L�=��QI����e/mf�sW؊�H�s����4�#7��}V�w���,�x�#�ꅤ7�����0�7k+�~�O�8�Ry̶�C���M��kd��E��1�'�E/K|Μ�Ty������U�$�߉��LO#U�y�s�qdg�r�Ȫj�q|F2O��y�3kHo$\QЋe�t�D�F���%��.��>x;�$����dd��<xRϣE�`�	ж"P{|�E|J���/�:����uV���헮��g		�4��s���M�fnlN�U3 ���Gw�Ԉ����<�5�.�k�e62��"V˦+�)�yS#4����4��q�X��Q���Ȭs��48��/5�ͬ�*&Io�r�J+������h�K�3�d��>��U�[�ܒ����ܬ-�2�	�o&~��p�M�)R!�=��۸�w�\	#�V��V~C[�j�ˤ6'q�K]O�%��*hNL��8頏��YQ�;Hw���~
O�\Љ\gK=�f�z��XeZ̤r]f���.M�U%zGߔ�[+�u����`����T�5�]Z�D�X{���
3� |l��Y�x X��ZT��ul�?���Kh��
��_naĞ����l..=G�;�7�)9v��t��7ڲ�2��n�#�_�1���`)+��sD�����G>������L\��ϐ�-�h;�]�����J��H�lsT �Im��`l�����Zx]!ʪ��B��e�$F�7��WeI��PQb�g���btA�2t\-�*��e�>��Y��Ǔī���Oׂ���	���+�^���"P�j �J����L8^��c5�ǹ���S/5w@-!�Џ0�ۄ:x�/,f��>�|�.d��F���k�Q+e����b�{��Q����x���z"�L���@�G�e�:Wu׃l�׭H����&�sQ]n�Z.un�e���q ZA�C'a�}/׵�RH�������	�H�r�˾��}��&�W���":�lu<�E_i�:�۲V�͍$��*�¹�����Y�KAܩ� �*�E���� }��P�,~�7"��D��O}֒���b��
� 	�0���G�i�i�S[QRMPnn6�����|V\����5W�?����='�ϋa����j��BϲM�����Ewv�5�,��
�CAH�����1V?�&Z]꓋,����B�S�k��F��]��WV�O��!Ed{ʔ]_O�i�	y��7�3Z�	w~�����B��YT��X^�Ô���Px��}e�����A�k��IoȀV�-sg��R*Le��(~��SC
�8����B{|��P�k k�h���}p%��ڡ�u��4xw?�~+��	�6��� �[=;�N{�`�ίFj&��"���|�~�9N�_�m�A��{{�<pM����o̧3
Zh)_�!�Ů�JZd�8���7��8��R��|~�����_/o
b�/�P�����9,�Zw&��ԇ��H>��t��{�$r���C���v]yJ�g1I�\s��h[���2�G$Bk8��'�CF(����������QBy��15�Y�{E�lﵙ;/>�/�B
�*egOzfc�B�!u4��i���ְ��Y�Ƨ��#<�R�1Iy8�vTM��CW�JqͿ�L۲��P�7V�M��S�>,��Xr�4� j0!�Y�%��Q3��$�'-��\�DƔ��w���W��
�~��]�'^���f+@�[��U�%�U�$��{t�F�8��f���z��OI�
W��$Q�h1���xu>�2;���k�ԋ_����A��?b;� %��<M�fB�?���ݞp@���OC�r��(>��
���U8
-�n�"��ə��/�Z��H���ɒ�]ʁgE���\An�x
�E����������VQ}G�p-���_���6��X1�]�~oύJ�T��PRS���(����?K���G*dZr�>�?��.(Է��W��#(���A-S\A�pO��-�A�����3DE��"A?w�V���0]/�Q�"�s�r���}�#	�,'?;�����՗`���� �B��;i�r��i�U>HE �߆8����{�}�m��_eK��O�W��؆��S�b��m����ꚴJ��m����^��~��㋯�Z72�Ea��J�gt��H�)��R'U<�T~I�[W�-.X�z�w^O#f3��\/ʲ]�ų5��.g٨�0���lQ�C[荬��-����4�c+����7��(f��bdU��nS1�w���M]�pA���2����O6�t0�?��DȽfʲ�E_��;��q�U��|O���w�W�ЙR3�k0q(cO�6�cq�X�	�qV��?|D�E���ƅz�&j�����.��Z��JZ��5��~�PYc�m�=�!��� �Ӏu�$d�߇R0�3�XRn-���ޣ��a�zav����;9t��y��?:�T�}}���㝬�;�z?�%ΊY���RD�?���C�B�,�+@�c#����P뛀���&W��\��M����Ѡu�%�z���d2��k��0.�e�7�t�2���j�r��wQ�� O�����s#؎g �尶��f!V��S�B��x�s��C�;[�<����n#��yn"$���Μ�h@�����5����I�6z�
ϳ��ߑP>�|"m������[yi#���
":"�R���}��&�e>�D[<�ð�<��#�IͲKp�c��I�M&�JN,���g��h���,.FqV.�"ɍ�?�
2rv�FH�h��KmoMg΁b�wV���|���l�K2#��q<r��������NS���^خ�������P��?]��\i����r�X��5���s�o@^&�4Ç�,���)�;؆��f��b:�e
d��`�Z����	�U�A�3��ͳ$&qO<�T�'��γ
����X����H�(�Oľ�5���:.�G:�{���K�"'s#�E��;���7v��6��fٙ+��-4�w�J+��
f��/ F��I�j^��1X�V�n��J�b}ߔ��Si\\|�!�Z�q�7T���`�%�7�@<Zf}>�.&._�������<�P��ks��`6�"8pŗ�EhS�9齕h;M���5�/��V�C�~�:�\J2\�<�H�C[�K���;�)Χ�=NS�ytsնAj���R{����zHv��!i��Q�:�A@�l�IA����Y5_K�O��$X$D#�|�1A@�>��hc�9ܨÊ��f�,'/|V��4UN�!]�hy~�F|�A�V��#B�hp��M2����C�7_ɕ���U������GI:����2>O��N
.��ί$��O����3�g�	��e$�IN�w�nC��ʧV&Tb�
�h�廒v�<��Q�.�l���Ih�٧V��Х�$�0-W-;5��Ij�R��� ��U?�r:��^�������j~/�۔�=��Dn�����j9W����k�e �gNڛr�e��w� q� �@���{�t;�2A�64���*�?>�^�jt���H���3gF���Μ^��\Y����Ҍ��r�?Bڕ<c����[5� m8�|i}(�י�cv��a�&�n�;L���#=M�
d�*o�Z�/���O}A���O�q�kɏp�+�i�۲��N�����M�-�F6t�R*�,�'�/Ɠ�`��B^rQ=yO�\����*��^n�$�&�cc�S��P�Jϣ��c��X� �a�ݳd��o趨�E�S�83��p��v�BK �>�K�d��{����Dמ��L!J�Q��c���W��U���ז��0`	�Xu�*�KǇ��;���T��O�Q�B�F��aѸ|5Zp������ہ�K��D��tZ�&�Y4�=���l���Lt�#�"�=��^%��*'��{Ȉ���|�$���PO���j]N /&T�]���.m�RT$)r@��Id�<��t��x�����c�ֳOp������dU��W��}t�G���V��.5�54&m>�F�� X��A���WH�� �G|��(N@��̻9�X���oN�αL�I둒��. �K�,%<u�٨Ũ����&4f�V	Mz��!�۬tm`�x^��D(S@�O��=>;SHQ��I&/�F�H!�|����3�����H�l'N<�l��$G+B��HR�`5�6�Sz�ϵ��*.���|'�\�N�M�!d"&�jj�6��h߃h6%z�Y6 M|.>i���Z�E�m�eǙ~E6������E4�C� Q�T�~�3���� ����O���y2�ȏiV��{�� Vg�M՞�����h]�Dl[$6e�)�����u�ID&��p��bl9��I�7}]�V�� ;�(u�E��k����X�S�C?��h	"_ϕ�M~|��M\����x\s}����
�����LB\���4���uJ/O�d��p�_��O�|��Z��\���h ����x�������3=�\_��t��[��C�\��V)��7�{?�>����P8��=�qǜL2�&����Y�Ŧ!!�����E�2C��?n �j��刪G'�|C�@G�t:��1�e
:�Go�w@��p �W3���h/x�{�3\�̽�"m��d�	#�R��~���Ԙ�%�_���{����<؄��5ăTs8�'i�1+*G+���2F�|�� p�0�MY��ӏJ����O���,PY6�Ǭ���B�WF���0{B$�ofUff���MԃY�5�꫓iK<��3.z��\l��{f-Sԝ��D�n�w�ԛK��9�����N�v����!"�58JGj澭�Z�{�瀎M\���d������ɔ�����y�$�!(����<P�d�>.с��_|?{oE5I�BP퇭��o/��G)�a -�/�/5,�O�gr�����u���UL�h��D�8��E�)�Ķǘ�]I:���_!Ś�◮���W����� �����s�	�ك!4Y��#�� �}��&w��W�i�#�i�`���� �N�$e����]�s2�\j����J=�G1��f�1��*�R�˱9/�K�@ߨh����\ȔA���{���Ա�N1v�۔Ѓ3z�kAHϲ2�K)�Q|�|	$��=OcT��b��Y�P��%�.�dCJ�������I��%�]���0�Ȧex��0 �'r�����!�U8f�k2S����h�c�m'�:��Ug�D4��{�j�!��8{R���=r��5�D:X��~1~��HVÅ�r!.�~n�������[=�M�>��Yy_	���m�C���ydf�&U�HǕ�wR�Qa#9EH�Y⦍��t��L���6]YB�`o:ڀ3����I��}ҍOߧ K�:s#�������1��ez�\	*�fz�ϭ��!	���Bx���[CW�r��s'�ג,��hnr.��I ����O����CќpJpI�5���w��Ə8��w���+��N��+I!�bw4�7��P"7$F���N��Kp3�(�:5����p̝�����2.D/6�ܩk["r��h������C�;x�n^�y���ձ��8�>�L��]>�MQ���Q7C���� ����PF!!]V���i �/�v�3,��町���ĺ������*"#gfj�H�G�--�3«{��eȳ��߁�Y`�0����٢�-�'/B͋���ʍZ�:T�ˁ��j8�T��
O�yٴ`Ĵ=H�EHM�����)����9I�cz��w2Z�T�>� .aַO(�x�d�_�ک�*��H��.e��z��P��KV�� ��l�M������O,�r9K��%pe����|���/&{D�	ڠx��ǐ��zh����>k 9c����δ8f����2�xl����[) >5��+aF4p ���;��,ߜ�S����~ZxR��xq
p���S���\�^��f������ɨ�������B����4��������W�eN��' wd���Z3��4�Q��18'l��lSm���d/����u��k���B��p��7a*�f�7+��	d"3�2�2�4��(�{���^����K��� �;�G	�OM�Y�Uԉ��mz3���w�I}����/O�/�K�l�+%Tt��r�@�>E�v;��0��m[]�|��M#�=0Pº��Yk���.�~���=�������г�f*��y��؏�����u��~r�h�J��K�-��M&ĉ�;��������T3f�,�=�f�T���IS�̡@0�,6"�ݥ�����
=��Tf=Zz�©Q�+��k����<�:���p��.���$/	F��m�>mx���=k�5Jڗ��Vz��m��nb�P���"�˂��z|���{Q����]dr\$���ݽ44~� ����u��Ɓ�w����KŐ�J�<�EIB�NU[�}J���]~�ym4v;德nc̝�'�:��m�z��aT��S��!������u � �.8�|Q��y�م-���~Fz}k��G+���E������^�"��k����ʐ�Xt8^J!���\��>l��Z�r��U��s��&kcOϭI
(�w<��C$/t|S|w��0G+D��Tp-`������O�=W��u�r��q�M�X�ȗ�~����2/ �(E�Ki	�m~j�e����]��+��������o�k[��DX�~��x=3sdͭo�5�o�B`���җ�
��j�ԝ}U�c��^��o,�w�v��XF�r�x�ۙ�84�G��Oi�L�M�Y�^D�P[3ŐG°Ǡ/ۉ�M�8�
xV+���^���h�
��B��>DX#�'��r����;��I�K��(r(�糎�ɴ��T�=��o�t7�l����!u�������f�q�j4�rb��K6�L��s��Av_�$d8:�S;�4��ÛM�E>�������HR�жS_n�0�5��E6�E,|�h]�rI���t�=���ɇ��[˭�<�1b�D���	ݛ��=�����t��P)d�!e_��8����l�/�E/��u������	̵4�c
�;;!��"N��H�m���j�=y�OgC��Z�. �h�y�ր^;��V�O� �b��-1f�rϻ/ˇ������䍿�0I�l���v2��Q��_=g��Q1�X��|,�bI��Ԭ�<���O����0���fe,���G���9���J�w=;�`���kĳ�&mfuG�uz'�.�B�i=x!�2�=%,6�=z�B�����a��g���D3L�p�$W��ؕ����v�� ֊�tŰ�{ю[lJ�'j��^Ƹq|���W���z�"���>�����j�_�7�걚I4+�u�=�ah-k�������M����Ǯיx�sFVV
����*en��yQJ�q�-��O;���x�D�אŇ�ڽ�ԅ!�:�&��3�B5�J�w�"FzW�K�0�M��T��G
,�V�Le�{��h��)�B�xv���D:�7{�3,Q<�����'�V4�eR�+��[�'3�c:��h��e�G��(ǛK ���=$��5��Q+)8���t���s��?�c��H���}�I�:i�  ��v�*bIP��zS0����q^���=�_��+y�� �̸�<�aJ�w��LL