��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�U�|�=����u��G&����B���>�e
7*>�cKZx<�lYy̑�����T��)�$OvPP����Mh�@���9=�TM�?�kq�(�F�d��|~�D��AeÖ�BQ���7��E�M��E���2쇧�A-<����T�jo-�H*����1M����cm�<\�^+��4#��<6�i'��.s�^�����P/�"�D���PSM���b`��m���-�e�}�0UW	a��$�rV����	�q~��-&��Y�ȅ��u%U6�]�c<���qC�bWm�����s:��ԭԫP�1{FQ��q�!��#`�Y��z5, a2'��9�Yd�vC��)X���?��L{Fd��kQ,YT᰼&��Ne_�ݓb�rURi�Z��׶�߹��L;.Zg�X�>	�P&�H��"���j:��F,��U�|{���7QE��ȴ��s}㵔��;k��h�d��J��DS��	�O�$�������<���!��oF�t-�\"GF3&��'���f*��/��^��d����Q�{*+^�1�u�����$v��1Ƭ]��}'�L��H[�vx�2(N���<=o�(��� ���a���)���k �Y�M���� �>�Zl��;,',�'b��Q0w�,��
{UABOO?h΢_LזS�����a�O[� eO���?)	�9}�'=�o�8֌}@2��w���l;pG�͛��C�`3�W����4�6�Oم.]�?{�N����;��lx:7l�_�����y ~5�PE4s����p��l�/� _�\��}��Wu �6�a�tG��0�e�G�V��
'K��'�\���ψk]��U�q��b�������#�,�}H'Y�q�kÊ���$n���4]4s�T�>�\�Ad[��S/
w<�g�����b���/�8d
��Q0�-0p��YV^�g'��^�F�A]9��H���,}{B� nͿ��!�x3$�n�4�����4�o��D�M!� T �1_���0��I��o��Ti�)���O����p&��¼��fH�AxEX]5 �?k:B6&yG�v����7�S�%_��f���b���P��L���8�U����I����MIE��R0�d�W����
�A(f����HK�j��y�d���TAhz{�i	|Id��,�v��V'�G��ADCpjW6�Ӱ�vJ��x!� n0^G����Z��O�v�#m���6�5���vu�cc��t�'�`�~>��=�o;y�=)��m���W������q�nV[�G�f0V�LJ��C��%��[z���V���m*�8Uy����-�3f5c�C��4K%���u����JJ�V^�y5Z@Ї��%v����Z�a�O�O�H�v���_�-(	tD��@�t<�L��~��2�L��N�L�v��b!�e�M@7��W�^�o�c���mD����]N��u>�03��S�b�}��P���/�/����y�<U��bfRztY�|Y�[@u��%u�)�`e�k��IW�o*ZZЅ�F}m��LW�����pP�m8�~��U��m�ڰ��}��}��zS��ng�<2����F:8�:?
��p��f��jIRy�׏5��<����mwuB8�R��!6�t%g�oFD��m�	�X��N��u��k&�r������?6�m�h?��/т���k�҅N�:]��ĵ������TV�_y�&/���K;��D�ۈ�rtg��f�_����`4����ѧ8��*B���FDt+F��u�6�:�9��D�oK
i�.$�c��5��m�O��m�P��mDi��?S�J,Ҋc.[fr�>Ђ���O��Y�i)K�3�n?��H.��'��dy�}v�
����	�J�aW��L�X�7�`�%y���@ޅ��uf������N��A�܅c!w��M)�1Y���jg���u6��z6�+"#F�ϓ� P9)u ��ˢ:��0)Ƴ �G��7믨��o�A�'�I^M�{�����uT�8JP�ZQF��p�X�G?)Bz�u�A��Y��UgL2�Ft��^pn�uj�(AL:hw]�8�D>K�X����P`�����c�k��h8��q���������]4m��?C��Q�qXFJնۧ ��hK��o����z��n� 4�	�u�/��X���~4��A-�"���y����J�B�B��6c��F���4_Ž����?�G�e��Ma2��q�n����#��{��B�{�0���a�k+� �B�
nP�bS ?�h=���ٟ9�L,��1�px���`)�bh�g�x��2�Ā���\8����SkE���|t���ՇiGy(������=�H(	�8i��ݜ?���ڇ���ͧ�&d�����2�6�K�j)<4~^��S�@M��e�q�{�
�n
��jAl-&v&	<��a0�>���8��˰��!`Gę�{��U򿫽�8��u�P{�����-@��:��uJM��ǤT)��S�[:��j���֠���D�a�D:o_'kbȜ5��0S��@3xWp��j��'��\Ҿl���@2��`D4p�/��W�uzY ���^@�lS8��M4��dU��ll����1��9�̎�q�=���+�O��˵Ly��Ş��z �\�8ߒ��?-ߓ��N����0#<	����[_�5Q��(C����J�R����=8zj.�w�]�\F���~�DO�]���])3\rW>I2CC���=����g�CG>*���'��
	r��<�B)� R
j�7����85�E�Ɋ/��u��p
�_�:�3�K�K@�Ӣ*\����c�y�~t ��j�/ K?�EXc���4�
�4�l�zB]@r��Ǌϸ�D�\F�L�<BX���(#R@���/�P�4_	F]�0� U� 	�*(�U�I=y����H�`Z�'Ga$�#M b�;��6��I�I��'�xw8��R���%�x���l�l�t���*_Ҟڐ�Pc%ȷ�Pl�<n�7y���_��`�p}�)���фp҅弧uj�����X�R��YN��n�����ߦ��X�T��it��M|��¯3Һ_@�͗�D�Ҵxz��Ң/a�)��T�Pm���CQ�������`8}�f�N�/����M��7T�f�2#cd3�;��2���_�1ޟ6�	-�u�7�m�f��[�0��MnG��?��X�{�]��Տ���V��������-u�[�&�}���:��}j8�9�3�z����l^�
�_.�n�P�>R�Hr�ќ�j�I6ɥo;&��湻�x��c�]W�u��/��+/�4Y�K�JH:����at��x�M`��qV�;y��r�Ú�s5��K��iPq%I*a�'ye1�6�dK�(���U�Ozhj���.R�]�@�[>v�q�R���}=�
9`RUO��Ak}8zgT�ح�C��!V�zjƠ��c��]G��g��)�v�����Q5jw�?����z��w�c������ź���Fu�-�>"��~	� � ��*��j���@���!Z����HW�0k�A�h��Vl��z>͘����a�V7QD͒�G��W�X����h��0n���BV��S��e�i�X:>t��`m��=$"���|�	�Q�Y�Ny�?__�?�<�9��rë����,���x+�!�Τ:p��E����3V���:?gi�������� Yo���u�1�ٛuG����WTrL�VR{-�}/���n�����ܛ�i�WhK�y��mA��g��[1����BzJ�E�2JǴ)m� ?e�,ɲ�
60�ň%�/ �^yX޼�:�ٴ�����F6�p����S������&.���ɉ9���°g}�I�9�(�&�¿	���gGUt����z����q����t���b�F��A��7��2�k�x��9~�X�I� "U�L���%7�����	��h�7`_V��!����7
���B��4X
�������y�����i�}E?1�5d��`��⥙�\����R�w��5҈w��ae��1��L=�s�O���U�A�A*��^�f)	{�,���0l*�Y���B��<T�`��J��3H�M~�.}F��yO���W�-��j�����G9�� �A ��e"5���� ��\崲4߁К@�|U�����R�T##^+-.�V�Ӧ���U��
��ڿH7�a櫝}U�
6 �kF�a�+!4�S5o_V�⩐���M�2�d�>�]�����8�A8^;ha ��;��	���1�%��ĔFA���䕶`�?f��m?`�珦0b�����h휅��}�&�*ZoH���!}幄xV���>����&�����%�Cӧ�._ZIS�?����	׃�$3G���&��~�?2��t�}\kL]ZY=�_�����4�L��2AD���������z1�p�!��xLĻK���ZU�Uw�-ݖ����"�^']�q�~o/54H~�[���͎	��,QQ���g�C�Ǎ�j���(-F��c}��=4g6�Ip{�@���L�?M�N��K�|:��Y��Ԭ�C"u7d Ϣ��BQԐ��X�W��M7�̜�
���1��\_%�÷�����za�L�6�_���+�
��UU|g�� 5���>�M#=|��̍������`.,��h�#o}V�Ub�8q%�t��םޅ4r{�4#��<G� �-Ɨ���{~��J铫�u��]$�'�>�����8zp��Ʃ.�~�84qŐ�Wd��+k���bkgT���
 �T����fc�	��fLm�����s�I����L�T�ŸG�h��gv�\��W	���h�ҧ�y�� ��6���G���L�P���}L��@>���,�Ro{�����{��4��^�N]��cp�sP0��.�w"^hV@>a��
mKoSؤ2>�Sˋ:�(�F+<���.^��v��!Z���:��EF6E_ha�D��x�I��rY����ɲ��E�� �]��7WP�e�k�7w��#��>��]��{�<���Y���[�����f'�k�7:z���0�wbY��{����h>�_�{��R���c��3��O�)|m��k��P�z�~�Z33�ïݎ�`�|����X�>��e.B�@�T�J?.-�(�^`�嫶�^]��#q.�dr*D.�n'�Uʜ�2����+'�,k�q�����w��ׇԄ}o�:	y��1��x$y�#�q�r�ڞ����('�-����Cf=�q$5eD!���Q�au̟e�7�sd�ĺ�)�>s0��525�/������iĵ��VWO|��΋b0�EH��7hh6�f�EN+�x姕8": |�sĭ����p
H$�_3
��G�G�($��-�vC;�����Q����??������+xߛ	��B�o�fD�@�F�HC-AK]llVr���躑��?�ޱҺ�{o0V��
d4����:ڠ���m)�Z7�� �1'l�i��՛�Yu�L�	�L=�QS�3�O���	(�V�z9�˵�Lb�8V][�3���%�f9�^7��O�-�a�_�E�IP�6]�>͗<�8i%����[M�Gŋ�����kK����L��f6"����Rz���rG���U�>�����53[�����A�R���[I	��⍿E3O.dïH4# ��q� p�V�h����OTD���H�-����WN�F0��*�ד���Ϲ��U��;�9}�e�V��w�O�U��q���k���ݳ�w��BJ#������?����mh�y�?�&,	�ai��Kb����7V��G�Fz0+��k$�)&���� \O��e�F���f銽Ј�tW�`*E��I�x�L��{�Ǵz�����ޒ�̌��fL?m��BM�i�<��W��v%D?8�{�|��'�����ˎ	�/���Z{k���ӥM��U=��+h��v\B��8�=��P�W>x�j��}�[	��<	�מt�\�?��1e}=�r�_����������z���Z�	�L��V	�q�G&��<�&[��\`<Ecwhڋz����:˕57q���,�l.w,$L�6#G'
"��T���5��������xoɐ�z�(��.�R��.��4/�^�чע�GK��r����Ȑ��yݮ�Ж��{�C��ӥf��I�pb]�$�z��:�湯��CC0�xs߱�����D�!y|�Y��l�~���f /~r�Xj�̤���gD�%� �ߓ��Qd�c��*P�{3�D
�5�^{�n��E��@�tt�hhS)��� Ǒ��颿�5~-�xr����ls&�L6�]��Q+ط���%�I��
���l���	a��bDNS��v�g��Ri\x`���j�޻̰�ʒ&qͦ-͐�ӖD}�R6��mE>�R�Ʋ�-���|߻T��)��aI���'ȝ�bPk:yJ�zy��m�:^4��	�����gJqiI��r?�j����|�I8dς�X��MzQ��0�� ��EGp\z��6J�t��jE��E( �6�S{�dز�Km�X��&�7G�)��m*��m����t4L2�h�A^�#�O��~~jh=	AsW.�����e'ٜ����F���m�]���j����V�䉒��\�������
��c�L��	���yP�=ͺ���i�§�ᣍ`=�rGT���5��pɉj<�l})���a�������܋ÿ
�Prbi���� y��B�����dcD(����I\�J�<��x@$��/��WY�����Ε�<Vs%�N�R��
��h�Z�l���t%<X�cE�ji�yGሎ$ǳO��R�}�Tt{�6�"p���kV�U�I�4>X����/p�~)jN��ݞ����<Q�!�WD����3,��Ȓ�祩���SNv���D0�6�i��S���y�)'��"'e�\���4Y�I�8A������}��=��}{CsL.�vr���l�G��t���A4��QE_�w�x�?:���^ 'o)r�/XqS���P�R8���4����Y�P"]ɞ4)�-�t2�⥻���L��a޴4S���_GVr{��`� Z�*󍉝n[ۜ�\�κ���E�dG�6*2c��jx�Έ���Z�6��ƛ�tHuJ@b�m�?�Kl�k����(���d������2�4A������6�#Rg�v#ʋ��U+9���
�g��|������A����v�����K���Iݸ)1�d�a���)�����yؤ�������h}�0��Kԫ����~*�'U�ƧX���Ym���\iP!q��k}��{�+-aB�3m}�;�����$S�l8hI�J`�E�sY��]X%��B�-�2E�v�;`.�S�HH�� ������Ln���f5��2�w�7�͖� iEo2f|�W�����C <� �n��ݑ�V(a����l��<$�VL��t<��P��;�[��y���*���oz���Ź�R������LjC���L����w|�C`j���]���k�0i2�-�2��zĸ�Z��C���R����A�[~E���?uM��⁐|<��}!
g���5J�����S,%H��_rXt��:�U������ܐ˭��HDO���T�'���?f���~O3�o�%���Sb�%���:캘�TV��w�����*~ �]Q�A�n���������c����4��9�yu�bN
��~ux�SS�6��O�*����Eb�P�|��WE<Li�C��L�
�$7m> =�Ƚn��F�T �J	���M�+�E��~ ]��J��b�,���m��r�9$mx�^���z0���u�.��c �����S@<��K|#��/	1�PQ%�ʭ\+�����ecQ:�&�(��
�b:sG2%1�J8_�"�I�ن�����E�
ͺ���A���D;�q��w<��;�y���43�U#r���%�5����B.���&~퀰�c�ھw�BX7�v����Yo���It�G2�?o��5H�yw�|�h!�&>U]lU�Y�8�9Bh��-���H>���W��I�.����(�/���GMR�]�0�a�������/�*��LnO��:�Y6�Q���ݨ��S	Rd�[�����;oM���*�5��]țcB�����x����l!a��T�}��1Dr�jc�!;�����]=���V��-�g��J�O�F��3x�1_Ou藰E�Ok�|z�@�f�3zR��Vr�KvNˋ�]�iUC��U_�MC)cgjr£&3S�B�p�(9���a�zԉE�doV)f%�(!/��	s`�t�y!v��J՟���5����"��:��
B|g�僶��=�@eW>�ށ�5%[.�6�a�a� ���n$_U(<e$#�kt���N
����։�wY5�E@� ���s���%���)~��ſ�E��p�K�MŁ�V{��a(
$/������}P578���J�Z%��&��ҳ��:D�%�[\.u ��}$H���Ի��g_���X�W�P��O��O���,���_�/�����8�E]��ƪ�]B����hN�I<|��h\���K,%��#���t�j�G�̏��*�Lk�Q��w�r9W���`@�_T��Wg���*���p�f�0�5y��DK��#�4	�.���s9�zp��,p%�}�PY����)i|�(���V����y�j��'��i���WxL�aO��,PYH�p�^!�t�\'�����e=�M�1�^��4�Z�"�v}0n�2�5�O����w���G�`�����<�ȀYj�M�ff�+����VA3i&-,hƥ5�c�e�Qg��Nx�M��