��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~�>:N��c<����x �o$��}	k���2t`&����ӼK��C�"m:�T99��N�,h8Z�j� 4�B�BZ�9�|"݆�3�,e�c�T��c� $Al8�0��� ��6`��@��C�~���!��To6�f��ct��{a�5Qt:�R��Ѣ�X����"l�)��`�����H)���\�$Pf����URڅȚ��Ch8�̠�<q��>w\�;���9�P�EyteT���@U�Ze�s�UI���[uk$0��)Dt�r����)�Kt��ځB7�V[�)5z�%P���ŧ)B����fDw6�Tq�1з��"�^�-�K�K�<ye�a���?��^���Z���[�	ػ�CO]q�}!���8��Y0T�����1�[��%ؔ��,����B�P�AH����jB$8�xnW:�=�-42�)̠"�A	��2�&n�K������F,�Z�� �X�H��`q��"�pE�1����:���b��IWk�d�Cօ�]c�oE��Jot'塗�^��EV�� �d�]Ҫ��pV��aN�yz�|Qѡ�.�{���<�7Q�]5���~�a��(v�{<����g���'o>�v����X����0Z��f%��Xi��R4���]��px�Օl��򞋌�ŅF�3HH���|������,�>v�
�8֞��ke�ک1�t�O��QE�V�Տ��Ta'Q��4ֶ+���{"�5��rI|R�]u�G~\�-� X{?��~`�D?�/�t�Y-)H+�2J��3V<0�B�����r":2ij�g[%㛃$������)���H&_֒�<+J�9H�w���JښE"��>�9�ҵJƪ�c+u������Z��� ������G��J�������Xø���iZ�0�Y��z���0��Y7��5L�ҽ�^`b���mJy�]b�Q����s�L�Za@\��(ń+=�SYI2��X��An �0�b��ý	(S�}VO�.v��f��e�.34:NQ�3�Ddm��6P�y�=��E�&���@�0g Y·�=���q��q/�8Q�	[�O��uf�'1R�v��[��etH�ǑJͪ ��Rc�[ImV0�]�)�͎��3j
������W�^	��!-�_�]�Q������D�7|a���]}��}��>��-��r���������6��JP�>��n|���淩�����r�lI��';�2=YL�{��ۗ�ah�@����L�0�{��@���5~r���D�<�hG�O���5쭧�4=�Nk_S-�W2��C
����m�QA
�.XG�����l(�;��;���F^ڕ����R^ڞ�v�"N)��/@R���5�����V,mV6���1��_n�R;�X}�B��ߤ(�КJ�ۍ�X>r����3���rr,�%Ç���L���#��:��D���/MKpqR(e�,���镫��FOMI���'�������'K��QC�1�ЍCw�8�c�,���S�5�B>AQ���l���uH���%t8t���(����C���CM��^�~qD�;|�viĔМW��8&|��֠_��̓�#.�,�DU!!��B�[n%xֿ]S�}C��!���7�^G����z^}.�9����L{�Sqv��*��0�D@C�7-K�>��m~	C@K�Gۓ��f~�Bpo�	(�9�L�ͰF�ޮGD�B0R�K		�@��p��2;��;س��^$@m�#�����1W����=1K��n�l�̮�xl���n�6���P����%��70��ib�E��.R;r6gپ;\ƴ�v ��It�jۋピq�@���uU+0$�r�x�������;dl`u�샫���w���T���њ�����`]�)B@4>�sb��ڛ�1������z��i�)!y0��6��F��f����aI�d��i�77ᚬ�7�Z&tA��b�NNK�d��,m�f��:��[���O�@��(r�>'���Z��ȮM���.��-��Z5��ޗ��o-�1�?��Q5�@}���!uB���/z#�[_B�7�	u�
.\h�`���@7a�_��a\אJsϚ&*-0�#u)f���,��{vˇ䲡?P���g�QʟVE5��=��o�1賑����|���&-:Gz:���-wQ�/V�_� h)k���� U#`$���*۪E���)�������䑽�٩��K<�I++�K,CJ�����AC���u� �آA�GT��!o�uO�s<���f�胄�k�X���S�,��Q�v�d%P��dWY��@�,�yQ�ϚNK��.�1�~�Y�$�9RÌ��Q�3s�ˀ��jl��{%�l�}��� ���ř���K�z�$���f�'6���E}��V^t���L!f>�� ����+,\n��@^�9��cEn�~��'�!U8)`��	������T��>IT�/
�� C*�P*2V˞:Vp�TT�u^3���?1��~��2I�yFWǹ�y�H�t����@�v �QC��=�W���<�� �2�Ф�L�c�Z�}k��e�h�k�/��܁�D������践_�>D�_I� >*��L�~���d�|}�x30����bV0���n�6���eܔ��)����������}0��cЍ�j��Ucǹp8��^l~�߈0�7 F�1��94�i�1tZ�H�H\J��4��:�Q��̑M!�	��ƳMV�=)�5l�����ϲ��l=��x��B�jT����q���)��"�F@�ܜ�ݫ��Q�
�� ��,Y

�ǲS�&���7����Kܨ.c��9��DZa�����Ï��5Ӻ�y� ����!�$�Q����������5�T�T���d��^rZ�`U�u:9�R�9�qHϜm���*���ʏ�r�;a�˞��q�
�Z����Ӯ0]��Y1���5^�+ېcװ���h0��2PP��yΡˈ���Z�Ta�, !���p�俙� 
2���$�⥝��m���r��iّ�?�U�ݼeyG8)������EE�ݖ�_>�G�B%u��%�|���uR��ꛩG�_�x�f>b-��� � Y١�l�F���n�����A���宅7>������Z�"��2YL�搉!Gë�M�� w���\+�D�/����F�'���W�����HM�a������l�%*OP�P�(��q4�)���*3��Z/�K�4��NuQ�9.�eB��8���I�(�V�r��`C����֊a;�u��u�ky�ֲ�_b����b����묝��_L5������E�����-k�H=W�|��B|7�Z��F�lg	�ʜ�,�w�.��3��b3����U4���MC�hްÂ_���-���cy���@�`��j�<NUe��9�	cu=�r�-Aݧ "�
�/B*?��X1�ܫ��ˇQ�]O~;5��g*&Ë-�1������N��Z�\C;&�>�-i��R��t�a�|�~$��mZ�#��oZ���f�HѼP��a�+⠲u���~���~�QIpH���2`������м���ܕ4�G���{ci�|��ب�H�J��_�4޽8B�=;�}����:�����`��o���g?ɘ+��W��I!��ܿ�ݗ&�����HīTuՑ9�O��p�c��i)G����7�ps������?CTC<gC���m���Af��Y8U��e0�>�R�[�E�D�`��`�c�D��԰`��FN4,���_��C	=C_A�P\(�?�zI��$'p�<9~�˫y�5��N����Ek[�~rË�dm<:�ء~���}���5 �O�c+�%��
H�2Lx'�P�{8������ϭ=���P�Usia�����O{FPg\�]"(�z�E��j$77"��� ��b���Ӱ"��!_�e��m�f����*tU�Cݏ�+G���3��Rn1� t�'ѵь"_��^l�P96y��vN�y��N̓I����C� �*�दi�T�����m}{"���ȖRAa׾�+X1�K9M�ҕ�<'�P-�(v+7Pl3��� ��M��e�?ܜ����p����mTv�0��yu��,����Ȝ�P��>E��}�R��_ԻO�Lr�$Y�V���q���W���L�XZ��#K���֬�ǘ�����8���g*p���bQKS9iq�֦%���ʌ�b,��y���A���m
�݂��U���[Sn�n7�^�h �u�z�̑��s�Gw�Hk��x=�bA���v?nJ^ݴD3!Mk5�o��鈖�=>�����'g��<o�Y�1��ju��>Y^R�hi-��aK�=b��jN;�ZX|
v꼰���$��� ����L"���Op�<Ϋec,�$k��;�兔�c7˙$'�¹��
�;��V|\գukFn�A<Y;�X�t��6�l�vB�3u��-�~T%Ӹ��5�hS�� 0��1��)d3�WZ[��~c;FV+��z��e��¥�S2Y��C ���\7�`�)cnb���lDή��p��L*Asr�lݘ˔�ɣ�5�~B����%�#Kk���G�`0!�,�_�Wl�V{ש���љ�������e�Q��!�\g�BS%�^�OZ��bp1͂��!�L��	x� ��y�l�|�sJS�4�׭�g��=�Eh���i
��5�4�h�9J���b[eGJ�`RHv�[.�Gs�J��UY�k�WrGL��W�xX�@��WZ� ��`pɐzoY�@9�9��مAKh�E�����N�׾#ҬXa����c{��P�7,���:ҿ��8�ڊ->�PMYiJ��Jˑwz������`�z�۸�[��n���u��R���av�,�v�����@$K;�Ǉ�7��w"s�zS���ǴƘ�4��3�IvJ8s�&h�W��N�-�SԞm6�ޯ(��}��;���AG�I�ɮ���Aؗ�1$�O����nv�<9�� �9ꎖ�0y���7�����#BٖO
�M��>�Y�$��\��-���23h��0q�S��L94fB�u��J�uŧ�N��OS��rM����&��}GK�w����j�>�r`����%�,g��A��u@�!x-�b�$��T�kR����8C!T�?w��ֈ��.JO�F/����N�Zl%7�%������mx7����'Ja2')��*~#��\��LzI�����h@��#��37�A��H�[U��u���%pǺ���c�
�x0B�f4�~1��R𵆷@��p����l���*C��}��ޚ�rG1������2m�=jX�Nm_���_��jg'팕�����p��f��߿@H�o� Z�3�k.vAe���dǣ̶c	7��1-ADx���3�(��a+�T`& ��HB��ơ8˥Od��:m=�1�X��l��`�n�p����?�;/����X��'��5�S�1ޜ�cDU��)�p.AI���94�����嬴��:q���o���.
W<�z�^��cӲ�?ȵ�L�W�@^�R==�A��r��A�3`�Ƚ�	)w�>���Z���#����R�k��K��F�W��i_���ݍ>h�L	ᗎ7
6J�a����r�w�L�l�YGY=Є��jh��*��X�O.�(��ɗ�uۖ�8����X;����C�I�i�%6�6�a��^�k2��'3��|��P	�3�^�-��m�o*���<-qv��}�0�t������O����;��v�Ԅed����Ŗ�Ζ}�0���ò�q�A��6eXn�h�ssOAQ�o`{);w�"Wl�ʆ�-/ �3�����Vm�C���X��x�L��ᝃv)���$��±�Yuh,�%%�}P��z�W�|��[~s�^�\�L:ȧ�>RW<�`\�(��r�8��t93[uj����Q���?*g�ak�����:���dKcE���lK�j0m�Q~��4�u�2p�#��!��s9YC����R�r80us/dor�3�rV=�A�[�R1�Z=7���&�!��4	$��<]��J����,��|���Ωr�jY1J߈@ J���3�RW�)K���pr��iA��Ѐ�#����b�|e�$4�pΟ<X��h����3K�8M�h��$��:e-�N76?9�If}y�LA�.��;QIl8��B��� u*���܎y2䰞�F�F D) z���%��G�^m�pz�y(�W���w�x���q~�N�� �/Ӡ�Tl�p,��ĺ�Y;��]
����������|�]S���Ƶ;G7�I5���������f��q��;�uV�cJ���L�fBB�u#��F�b��`^�CS[��9�p�wW�$vE�	9��/�;�q�Ͼ�Ua�u�*Q_CΑ�:�!��Es��6�'����^�/��+�̺b�����4ȏ�[�M�۔� �?.Suq�6w���ic��'Kͥ!����x�))�S`M��Io=�ޒp�iK;z�c�!z--LŹc�ue+Ψ~�!�[�՗BwV����;�Z�i/+e�/:�eg�Cˆ���t��l��8 �&���t�?��K���2��vBC	�H�;��9b��� '�Vf�p���P�rd̥ph� �H�w��We@��%�C�M��R�*�8+�}��40ړ2��N��!]���ʂ��A� Fd�:
�6�9e��`�t<���ԭ�\Q�+�?$��Խ_k��蕩�^�;�(E`��m�a+�p ��|���-FGD�O�ձ�9�<T�b���K��/��Y�ڳ�t�~�������m��}(��1tv� �d��%�҇��Ұe�cL�;(~Z0��ܺ��]�VGڄO;.����(�`��M����M�h�'�Uˁ����j��a���fE�&<���,^�'t��b�sF�>�����v&Z'����gg>���]l��C߸H��ͱE�|��0��|��;���b��
ƛ�9����{��6j�%���m;J�5�5N�y���R����8��K(�$1�a�Pg?�d�q���N�_�"�H�M�O��X�cA�����dQ�s�͠�ŭc�G�@]����q�lA�f-���r�~g����)V mʄn��3ڪo���Z�(�����*����Ey'���+�-��Ww�����9�aX����A�UM�fY�D� W�j���I��U\i����V�~�{���jA�H�������8��Oi�g��x�z��C��
X��8�s�� _�p,���b�I�1�Ԗ)�t�U ��Ju�7%���MD�z=Ḩ�U�t	ifO�W`Q�WȺ���V"?�ݫ?��C�p��M-f6�^C�d,8�L�s�>ъ�>�ԅ���Tc3��R��"����l�����_�E:����[�B ]l���}T��f�r�4��{$Bd**'��S�x�s[�i�`�@�<(5��#m��B��z�xU��<N0��r�K��n2�;X�)���2������G4� �G~[�]���oE�Lk�4R���kM�I+�a1����i��N��ٰ�źއ�䖿�g�aE�T.�"��J/$N�X��l���.�ߐ�2E�"���):9���F��дq�,"���D:����������I61d�id��gj�E��e���JԲ�����N�ڲ.����L�q¨�r�=�����K�Gc}�Ǥ���ǵ������H�3�	7��k|�{��� �'ƅAz$�~X��HM���M-G���y�F�� �z�3h�1��b��m���֠_t��L�4�{�;���%"A�Ăm0�4�x����	���t�+ĵ!W�%c m���F�!����^���'(.-�ݸ;f�/���
5!C�'.�(rҴ	
%�����L#,z��xî�;i���G*�)�-ɏ��D���I�0/�`�uz��]��;��=[h������[Y�|��e0G��q�����"�׎�وbz�g�p଀�"�Q��c��
������ؿ����ŵs��Q!)��J��O�lIg\��OgvLBԒ��8�VT�6��b��:GY[u��N�MI��;ѡXD��:�J�l��{��Ge�9���O�Г��Z'2±�d�N���0��p���=�T��ҥ��oWb
��Xqٷw�T��P�����1*�T��"2���f7�l�g;��y�����[��*�ҹ��"����F[-�L����oڨ���Ĭ@���#��Pdq,�f��u^O�Wa��y�@�ɱ�B�u´����_V���~�[¿و��dZ#��6��)�q��-`N��c���c�6�`|�V�&�<Ǥ��1:�<?�J5���s��9cx�u�'�5T�� �Q��k� �~���c4L��I;�dٟy�4*p��_�4������$P����LXw��"�������H��c�J �A�|x�.N>�Ͱ�M����b����>C#1>3K�Դ�o������P\�)�Ԟ�_�>&|�v�w�U��|8��:��p@���?U	��Kf�R��R�t �37�\+���f\_"���h?TP��1q,�P+�����.�( K#&�h9���n�	��uF ��\(�w