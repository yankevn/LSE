��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��?�I�J��x�H���3�2n��jmݣ*���%��#����r��a`Y��X�9O��Lii�A��P���l�M'݋�܌�
��*�����)nš�`#�90��a�z�Qy����FZ�fE����C3��#�Qw*~�JxA��uY�S��w�O�v��A��a�U�q��5m-�WZ|�4@-e���˛|/\5�@�
_ڄ�����*�a{O�V�ɮ��Iw֤lE��sξ�^C�"hJܨ�ɾ��8�FUy�!�ZCê�4�����ʦ1�f�RU���Hn ���ǇD�L~6�5�4.�G��>�-\L�ľ\ܾn�$��i�C� o(��s�UJ���SG��vڸ�m$L�f�,`�t'��?��Ka�V�aM��S!��3��`��M�&��8z%o�۠$��6xh�YUM�D��a̅,=�����v�	[N�	>;&��<�6O35�I��A�pg��aPR��'�����&����$����h���Z�<�!�^��ͩ�X��C��(�:ѩ��}��?�]���S�dp/����t?̜�����~@���"��|�e�Q�aܳ��Ȓ]S͋oZz��x׭��F#J?�����0�΋"�)$В���s��MJ:X��PA����'��)�-�s�<ߣ���Yw�@�����M�6�Т�2dM5�Ks��'����\������g��d��Y�6]�ӆ.��?��iD�
�|݁���x�3���Ff�=^M���m�<h�u�xkMY���%8Nb�<!V�*���o��M��Mݓ�L0�- c��)��q���/���ld�	]z�o���-N��YG�c�PHW��69�f���m3����E��C������PR䫑C�E��UP1ړV�W�����TĿZ����y�v[�x��)����2Af~��E�b�	�2'k=��bD���Z����OT�jM��;zh�Kc�b�=^׷��v�(>tN��5sV{u�W�)Xa�m�h�On�{��e�r3�9E�捳c��D~6��U����̣I�@�+
R�s�?IF�l|Fx�6)z0���9j?�";C����*�E\��`$t�]@��KL#������f.��%�cFjO�x�S�7E	p�Y \�ȱ����/~�)�<�Д�L� N+.�8q✾�5$���=Ƨy|e����"hX6%��jG��^q�m��Lq祖R��g�T*ͦ�����8L��\⦢�F��9�T�Lû6m5���<֫�X<�&0�_˰����0*dj�{����5�BhRS��7ہ���3�/42�F,��`,ǖ/�ۘA^��?H��NL� ��+�u��8�6�b��z�di���R�s/w�-�����J�k�o�®��c�s�6O���w"������R5��>�R7Lt@(]�덝���������G�+�W���M����^u�?/��da��.�w�M~�T�IL5�Ҋ��'~�/*��)�ೖk��zY�\#P��۵�E��G�9�T-��{ZF�Z�}w�](5)������"�m��$2��*�\[�lX��������#�<���.�|c����8�&��ˢ�]n�<��xx��������?tg�#t� ���{c`�rp��K�_%_x,W�nɲ��1K�(��]A83'��?"��&�S!��QU,g�4
뺆�UL�#��,���yT�5�FI����i&,N�l_>�x�p���i��1iW���|�/�'O'������.e#����j}�x]2��d8����(1��="�C�#��٥6�*k�jg�r����V��&ҌE}]��W�j2�b��q,�a�k��~��mx덤y!-����9��5�79,�A0��7��b.L��b�[�)V�e������d����Am���l|jaM��8Տz��᯵&`�ǎ���x߅)��R���Eha�Ppm0��T�N��/D��{���o1O1�'Qh��4*�=d9Zݨ����ţz鐥N�K����r�)�2�4��z�B��K��n��\�!@�'_&~t[�|K����TN�LH�[瓿�S�C����W��݉3�$�*��/}���Qǒ�L#FG�w�����oѥ��n�)��V��zQqa���0���cb@`vg�Q̗J�^=�u��)e�v�g�H�W<��
@�p���O���@r���0T	>t��L��U��_�׮�v�;4Aq��?�R�3�F�L�y�ۄ�H���u���g�X�*��h��cA�G�/�#J\�M^.��i�+�_]��y|�ua����?��T�~� ����=����d�I.�j�M=で)ԪҘ��B=�IF!��v�e�j���F���)Mr��vW��'}��9��{ܡ��bX��ί���T]F���)B�'1�]7_MZ���T ��Y��ױ%�d
�s��g_"�5T^"��;�x�5,}��d�h����>��5��"B�m m/6ש6���e�����0��KM��{��r7蟷V-6�7�ߵ�qN#�EV��u.�ç������@��x�1��8���w�f�w%:�>ĕ;p�긷�V�B%U�yZ7Oxoe8���)]-��:�hV�p��NB/�'��LE*��y��eݯd?�]Ւ��`�PIU�9Yߤ}�����J^��0�Pe�jk��Uy�������+�
j�Kz�K͟�~�"�[S��>d�U�g�1�+�2����%�:�*ySk��?�]��j���$H4�/ "o!,9�n(K�� ��
��մ��ˢӊ�F`c���f��a#��������<W��H����V��O"�p�����=��`���(ZM.�9�ar��n.�-��|t���҇Op���l#���h����o�rc�����,�%��oO� ���� I2�r�^�T��Wћ�����̐�[/�f4�&��  ^��Ʀ	��Z�0]�L�@t檝���!\
(}�;�j�ͅ��5+���b��A�JO>E�@���.O�B%������Aqq������@`ؿ#~�m+�ݭ���`����]kO۪�N�uZN?�Fl:�+z@�y���	Q�C���}4:c�����ௌ�{F�t�3�8���2s�x��?b	�?���dv�j�]?��x�"�_�#�hπd,��`6G��6��0�]NYu��� 9+_/��B@3�٫���o7��e��׵d�N]�as��/
$�[I��d'�3Ċ�#���0̒��}�1��T�)w�)��鸪_'T��q��Ϸ�H�����ܽQ��f��.R{0���(�L!��<���j04�pz3��)̭\E�LȘ��-H��Cg��*j�k������{���_MG�D%� m���S����1����c����$7�p�+�A�U��^]^�� ��Rs?���Ʋ�ڲ?ccP'fJZB��.�d��8}ij�q o���ȃ~|˺Dk�|����!u�3��6�	-�ECVbK�#��FX���D�� MV��Y��Tj���ˬ��eGT����;�L��1`�-�M\dk��A�A������X2/���N�dY�?9�)���鄮S U�����8�Luh҄�l"!�R�z_;#HԒ�Kn!Q%�-�����V#���v��2�@ePu[_��nF0��ͥ�Mu��W	p�YA����f8�/Y���lF����5�zp~�v�C!�P���O�.q�?.�����R��<tz�`��Z�@�ZCK���If�u�DX����v,�j�(�qZfVa(��V�VyQ�Ǹd{Ժ~Czٽ�cl�+�mm�qf���[.�WSj��D5*�'��|��4]�+l�D�����#�ǘ�����-r�<�-��Oa��D�^������u����
�~�ݏ�/��	�QV"��ؤ� ����JD:J�El��	����g�A�Oj��w߻���cxJ���+�t��z��+˃�����@��cn,eB����P��y�sSkr�����h�O�'j$1�� \Ԫ�L�h]�q"$�i��ov�Hh���y��m0>��G�>F����'�	Z��F��8jl�Rz3����U�ct���4g��Դ�uq�jyJ����.�����-�"Q�,��\_f+��0�4;�6�n���c!s�1�g��J�ZA���(*[�櫀����/�4��=1;*�0%-����H �ĕ)�J���hoS��j�p�۫U	�ӳ�?=|8_�zL\�RTa��-(��SV��X��r�1<��\n&AI#���)Z`z��k�6߳@�~��\�A���ö�W��w jM�@i���g�c�NM�d��	��xd)750���P.qB�?�QF���N==0�+Ӡ��F���_���� �^}T���.��U��)1$�\xZN���r���ʆ���o��ܟ�|wS)�L�t�&�ه�U��?��4�40XG�r�R�c�yU_H�SU�ܳݫX������V��^b�'�=' ��W�N�
�k:�Jy���/��IQSoZ��`撡]'�u��tW�\����m��
���ي`��9��5m9��YkYנF��9��_��|���o�R��)M�ui9�H�Be8��e�Ɠ�+4T���^
w����y��0k~��V/_�c��)�����b7�lx�B�_��-V��kփ�w>{�C"9��Uy"^>���A���#�e�����p��w�����X@Td�ú>萴��Ъ��o5��+3��-D���H;�H=�3>�ؕY�l��G�--~+@�w���â�U�eS��8��f�LN��^2H�֦^ �Q��4��mL(i�R���!Ro ��9�bF���/�^��u[��O������	������R"L0`��AY��J$�G�-�d��E��u"�E:���V(�F��-0�܆)V����h�^5W*}%�ݚa��<s'\�x�k�Shviy�li��5�@��J�@ƥ�Y��I"Ι"�^x^;v���"�Hź<"��L��1�y�E�ǵ�}����3���c'���h��J��G��	�&�i�&�MQRg35�|������`�@�!�K������$���1e�o�ɭ,W�]	�����d�v��"��
ڽ6{�,��<�a��lN���8�>"7�h�f�ޗe��Tl /��^��R[0� J�^���b��e��:.r��Z�]�^���x*AsU>�O��'mDF��	����$b<A����n�wm�u=�{V
�=P�D�9��	�$�3ku�%�J�Q�^ȴ�晴��S����q��J��]�����o�0/ƓiR�z,^�\�!1ZK��W�Bb`g����4�$>!Տi�k�J��$�9��VlP��dc��ߡӛ��2�H���5�R�B��]��M�r�0�}�/���;���v�IaT��S�,�rMd/�e�8��+�H�a�@Iǔ�8�֒�<v$��j��t3�|�8�C�2(����U�:r8��-=�tI�U;*/j>\y�-�=���i&_����Ծ�
���ޱ�}�� t�E(�H�E-�&ͻ)���a����X ��D×eζ��/���n���=�����HK��-�!g�bN�׭ù�����e�ב;�y��/�'��=�� ��!#�ϋt�-�,�X�D�ެż�D���#?$!6-��3*9:J���s��^u�U��u�j��.R!.rx`py��7��<�Folb� Y�B�ƍ)Ch�Ѽ�-j�y��S!�<���T䑎�s��oiw�AD��,G�4�_	L��KVv	Q�#��Rȫ2�4Vux��^�Z��њ ?5;#0~������ �"K���%�}[��,Jp_K92�~H2�p���W����mk=wq�;�X��dҘR1���Y'��7f� �r�>�q�1��鷠��s?�ƧWyT�➣�`��8Z�s�����dD�k� �)�����&�x���dl[T�տ��l�#+���L�U��_��^g����|v�R��lW�*�iY���L~*��[�[��6��5��o��-����^ux���1bR��G�$HԼ=3 q\� ���w\a6+E��x����\�f�k:Qx^D?kޏ��B�M��_����7y1L��j8��	$����M���.�4Z4e/9>gOA�Ҋ��Ob�<`L�M�B`9�Y�A`�Q��q�h��leB���O �ˬ(fR
�x���>��o��	��8�r��Kg�+��!��Q�(�E���z������1��?�+��H^@�l�����r��Dh��q|8��l�H�W�V�%x��ͽ�����;A���Ĩ� K�#�$Ė?�ӓW��1�य़�l8o�}���\�n�X�r�P��j+����`Ȃ	��|�ݼ�J�x�i��t5jS�	��L�]`�:|߻���K�I�1��#��r�uӛ��Γ�
{�q�D���� ����lg8�4�cȬ4��=z�џ���!T�|�BV���Z�>[7{�[[��l-�k�"��ۥ���O�A�|����a���(G<K�<QB�8TkK29�i��婖b)��ե���|0_��<.�PKh\�+�+��-}P������?� �r�3��I~��K�9/����?
�y������}}�U�Mѱ��3�O��	p�_w�ic젔���=�:UscG�^~2DU�t;�Ϫ!=GӹK.H/���j-�?P��>9�=�m��K��@k��?n�ē]��v�i����� JdOv4i�>o���HOC���M�IY���c>[ii5jk<a���u��;5�t�J���M�pҞ?�Z�~}��q	�Hą�FGSc�5C�� �Rۃo�b�=���������)E ?L�.�3�/�����T����B-&B<��m�Y����>�h`!�~�����R�f��@�="�7a��,�u��
�I�Hf�K p4��(.)��'��*w��� -i�9�L>`�L�+B4f���קP��d�9��j��9�F�xz���d}�f�E�)���U���9:�;67�m�"���9�(�LV�[)��.�I�W�ʠ*�1 �6h2�u�-C���=�d���,@r�by�]��b��Ns�AG*�*�:�PX��j�~����C��c�Am0������n�,�)'��Ff[���G/����ˉ��pH��Jl�K�����������_��A��uΦ�|��`[˩�-���
ø����,j�K�
���:����m���{!��5.��eѺ��2�BQ��\����w�Ųxsゔ��u�y�@`���L��,��y�j����֑��@��Js�Y�#�d�aE`�K��%�8)��|hd��7��ի�^�3(#!��=�T��3̶$��G��_ћ�A��!٬\�F�@tV�]��,]5�������$1��Q����_��-��vV��v�lAd��� h����Ң�������l��'?Q K����R�~?ŭ�t � �d�W>_�ɋ(��ۉ��X������l�����;Ra�ƃ
;_��	�e��u��q��_kW�8��5]��W��!7��B��J�Md����/�k�Y����	�rˋ6�l���5�$3�v)����Z�mA���܃F�����Ӹi���k^��-_�Ź��̈́!e�VS�������r�lx�O�N�l�!y���V�e��⢋;~Ɩ��-\tf,��;8�_���M����h(�͈�/���r`��G��{%��T"vS�~�:�%#C�o�
����|bһ���	��9k�_ g���1.~چwч��I�`�; �}��4˖�\�O��Ұ�o���xM=���M�� 
\d֠9 K飍��e�zR�|�u����,� ��t6����甜SVM$��+�i� �`�4�.�����E`�o�
T���jB޴B0W�'؈�F]Y�B��&���Z���%��jzW��lt�1�x}�lA�=%� 4�"��Q�6D08�e�����$]mҏPƄ��ӭt
�I�C��r�,e�-�P5��Do�����%~n��k�ƹ����=��>��w�M~=j0��bX�"�gOT�l���) �z� sU�5� PY�E�wxF>"�ړ�(ޅV���$ф���8�l�ķ^��Vn����� &`=7��P˗0y���0.���{R��	�i���'��,rn�I�^A]]����e0���nmI�S5�#Q�-2(��[j�;�F���X኉�LQ�p����u��h�d7	XfY�Z鰮��%b�t�j�>2v�"��U-?1d	uo4�1]�o�跫�[,;���SU��6$KPӞ�Z}����[��A�"b��"0��"�<��7�k��P��ζ���s��'�����z{�T�Á�'�L����mQS���܈���:��69��d%��>�jX�Z��^+4����"��;@r~��pym���6͹���2�%��WrO<�=�1���t��$���L�����(�4���+R�?ru/�{ƦI����=�p�~/�vJa��|���uI7E�R/�
9�����K4+��,z���̟�׌��۝ �~�&._��d�E�1�G�w�D[����`nN������ƈ�SR����b�F.X�|�I\�uX�l֙u/2�!OyO���`|鈒|�a�9�r>y'����D��{�"�V�jU���x��c�+Qqh�E&��,s�+��vS�^� ��iz�]}5�\ei�B&��P�ٓ�̅s�m&0�6n�{{�k?N��ߥq-��Z5YW����� �m}�Ƴ{��{��ȓ�ϰw*yG"@�)
�.E��>�ܖ�2E5\��#Ǳ��w�# O�kK�S{�����Uy��l��߅ՐM��J��0�%!��n��2 1�vy��h��h�;�.�c��:��R�� -V��� �*hXp7?dJ��w5�D7YAs���`���.��0�">*��"?��d�_��H�q��C,����P��8{��mL�K*���-�T�4����uJ��_!�\�gr���!џ��V+��b���kc����6�N��k0v�G��N�`RZ	W.t��|��HX�m{�f�* �A5�^oi�@q�=��[������"#�(�Nq��v�E&f�W���M�^��#ڂ�o"��Њ��U�蝲J��?T-l(����}E��V(�P|�g�_dզo�=�O�j���_�+nq��i(h��'�@օ���Q`^��q���iӱ65B�@v����)�/�i�
|�Vu�&rڣc�%!(�҅��5�ܷT?��P1�w=����Dm��Xn'��&���B#Rn��y;����͕�3+	�����]��2C�C�"�QfKo��&��.7V��L���!m^�G�3��+@��,�%<� ?��gD���������{-��U �#e�/����;B?Z�&Vke�"E��.F��5�f��U�)]�CR�w�)���F��4 �Ց�-!�'-y&g�'�Wi)�2�&J��5T<�O�K������)�&z�����Zw����4�� ��~CI7hA�_C$3u�Nȡ��yZ!�~y�n����b��7om�=Gߕ���������M-( ���x��A%��N���ls� �MaH�:����U�J��o?ڕc,�o���"->��|���Cn�RC�$7.s�Ը?�U`�}�vѳŘʻ�#����[��8l�h�Mzro��k���H�E���K���k�^< �����bv��.�b�N	�����M��!��ٴ⟆�n����^M9�%j��)6����)VZ4��8�%Or���0�8����^�̯�DIE�-�L��L|B>~SЯi�d���ysȯ�}faU���>�[��#H���8�}*��7[�*L�pBkeS$/�St�:��� �:�Fè���jUe������~��n��j�GV$��E���ae��*4��~�W���a
4V����>�#B�kdCс�
�\�oq�-��)ы����"�f�K%���i������κ��V(sJ�2��U����{���RL��%�дgFD-I���h�9hp4�UAP"M��-usϯ&��`n�x>�ʎ^�D\)A��O<O��Z�i1^ov�)�8�f_b�������GC_]�^+8���A_|t��c�i�%CZ���6Nx���
g���ș`e����f�T!- �D]6���&2�B�3�������)��'3Lg��Yʠ)�,��
�e�
�Yb5���q�=�'a�?{m��?�o���)+O�c����X�:ߺ�.��i䯥�36�"�E>%��T���;:>�P��%1�)�E�_�w/}a��8e6_S�8̭я*I]H�L�/��W����V��"S�t�|�����3��h��y9�Hfm/����t$v�T-�Cީ>q��֜�����;�W'zr`����$b� N�qdJ���[��H�X��
�꺣Z��O6]�(i8j@@�/0��*}����������7��v���'r�������5!�&�s��hך&ܴ��m_3Aq�՚+���/�<un���ߣ��@��[�S^�gz:��-����N~#�ݬ�cnP͠�]?�����NƘ%w��e���n�|���^�׵)w�72�x49�a�8j���SƆ�2l1/%/�����p�8G�L��[qCՐ�f����1�`ֽ{��3�ć�դ��d�������%
@�wg�L'pf"`�m�H��x��=c^�\�*����(V���e���!�stI0(��n�z��2rp�h��l�
Ot�-��{�=���n؟�W�Ê/��� ����kݸ�;/���Fk�P�"�@����"�1�$�lp����鸞�/X_���B�ש9��W߶J�i3�qH�e���Tn�Ռ�a%uҴ3�2��0�c�q����t��|�?y�.
��kDtt<Yۖ4���āV�!�TgGN����ؚ1�STe��I�	~E�����`� �@}Ijߚ!�BxC�LL�1��SV�0�g����b�8a��][o;PX��-fz+��Q��Q����d�,�%��L���q�f�	''{��M3�T�,��sئ��伹%%�/]�D+�[u�q�aot#)�_�t�׳'n����&���,q:��>4�6tT��T�PC�H�6U�}�׃;��b��3Ͱ]A�&��c��xH�f�ȚTV��L���ڒ�Rچ�U��U�9i@k밍�T<1��@�]��ʼ<Z'�å�D�W�Fر���Kӗ[.�C�i���[�2���^�5���$�|Z�Q׺(�qY����}
T�����#@?��-V@f� ��}�/7rCu_ɪ wLn��w(H�?4�T�}8���88N�٫����E�`c�d�b�T����2�D^w�R�:_m^%'��h����Zo}��CZ4�����Sgp��D�f����]z;��Bth����({���.E
�0?УipB6���&�Z�偄1�����:Abǂ�U��W�K�cG�g�2'��=7��������ʽ?���%*/�O�=�~`������d���7J Y�y�!�= /��:��M<E��Lp���n"+�\�n9LQU6:���j2�d�t�z� �a?�{�$�V��W�EWJd�~M��8:��ǎ#H6/h~/B��L�}}��	Z�]���E]&�W��w��/ �n٢i=D��>�,��l���:�H��0R�w�����}�2�T~��_J� BR��E_�ɥ�4A,u�]���LL�̃;ՙ����l����U�Nq1:��Or'* ����Ԩ#�[3Q��������h�R_!�,-`ylS�`ÚUI��ɦ�F����G��f^|��5>0F��1P�r����\��_�\��s�Ab��J�Eroa��9�$k�W���U�X�r�7ͼV����5��Ǿ����R��;����|/�D�`
$�$+x�jH����Ċ>tW;�qƜ)��]���w�t�4�&���i�J�pI�1��~&x�j�ɶzI���V��sB��͎W]���L�p�LK���#F��Lq7������kn]�>�e;�d~�ٍK���,���05�QQ���x��kR�d���r���Gۇ������c7Y঎���k�|��%����e�Ə��V�h�b::�W�u�؆�Z'�FB�?�����E&���ޖI�����i�CS'�������D�j���\�t���Z'�����k9>��#�4z�,�E\9ͣ�Sa!*6m�vc��H:W���[S���?���|o�ن�m{*�N+J�O��jZ^�,öPY�KWAE�q"�oҎ�B�@7Q�PcmI	��9��S�(�������@w5$Υzv���I����:S	��O�clFݮT?��3�o�m��_��Z���]�߷)���F��)R���k�a W��dy$@0;�����(�����;oA�#ӓ��/G�Ժ{���L�6ARt�m�]�¾'�Q��������'wl�������q���k��s��wߏ�y:@vN�Sg/�e~��pt���s�E�S�s�/ u7����'�1�����is�1ç����
GX����N�� p�M%}�T�PS����j�ی���ωZ�u���dC��n�w�|�d�N��ƹ6JR22�q� ��{h1|��l�c�b5j��?�b���3�p,���J�h���$��>�`��+N}ND��S�А),��!���$���|[z7���Ks bxנ�1;��8e�|����-.��d�Py\�7�JS���ҜL�eG���S�K��tSk4R LI�|R�I1e�n�d�b��o�R�(;�I����2~/0�G](H�^��*Q9^c��W;B9᩾/6X�h�݊cQ���*	X��	g���o���� ���U�V||������я���M)7D �z������j׊��0���}���Ҝּ#���ġ��̤<|5����:��u0��L�g=�ԣ�EƷ�������='���;ge�� ��L���N�K���&X�4a(D~�B����ty��W�ǿ��ǒ$�f�T���"�ΞP���t��z�#���f)B���B�#��Xx�bw�$��yJ���1��m�@��)�,z��P��{򖅉��*nk�v�^��r"�
+�S���kX,��7�:`t���Qr`�>����nBүK�إ���
��Ͷ�fc��i��{aC�.��o��@���8�;�3�{��I�r���dc/rZd�'i�
����@��K��F�t�a:�z���sB�N��`+%��5R��T_�A1�������1=�+G��g�����l��m'a�pb
����L�FD�vós�e�Ɍ���<�U.��Cs�2��z��d�	kzb�32ޮ�2��BB��#�x�&ƶ�x�O����0���r�;��{%�y������/�y&��jh�х�*���wb���P�q5P]bH��,s��J�.�/�����G�EE��A�K�E&o$�eT �4!����܈����P��V�4_F���i�R����~����	V.^���Et�Y<M��Y�l"L����X��O��_��,b5!9r��IX!���ɭp>� �&q�z���x����.>���x���<��k�3�dlE�c�p����
����t�P~?���m	�l/�� )�0Y�p�6�������K���>����~�EΧ�(B��k��>=�u�Vp�B��Z�)�'|�w�&�ڐ�[�oD�| uP��-(�6���W���/Q�W}��Ny�Y�,I�Yɀp{�P���5]t�ރ
v��+|Ȁr�|���HP��r���]�V���T=bt<i=ϲD����L�fw޴���vK"���'�i����'V����L�z%:/ז>l��
0y�8�D<x�Ɓ�V�j�BP[Ł�-ؤ@��ԯ:(����<����jB85B;����2 �;�w�
�h�	w�� /w�����ط���,��~/��u�rm�l��SFfJ7��ˀR7��Z:Ns9��� �j<$�Zb�j�1e����A��Y�,���������:m*�Qx�pﻡ<k?�pzHJI0�{�w����V=Ds-�EƧI��M�����uv����O�aY���í���@ �6˫���s�A��=ul�����_blo���g\�Z����ܕ`m�����B���ע֚V:)Q�&n9����0;L�f���"�w�4$���눫��c�*��U*�ݴ���������ˁ���a�Y7Ԫ��6�k,�D���e#�����.���I����2�V赟�p�A�M'V	�����z88X�T��Fϛ��/�o%�'����9:�hJ��՝p�x׿p�_�L�t�4�	+<�oQ�g�>��}�W�
�0!��Ł�LM��l��k�Π��y�d��C�m����ׯx1DQ�x�"�h�szwo8k%H-+������6]�+�O���z��z�pݳ��`����p6��a8ᦱ�YC<���uO
m*3�f���nŃ��z�mv�i��Q�����Qj���a�T�\b�2Ti��1����C9MAE��8�U�R�Kq䧧����!�ՖЮ�H\:K���lj�eJz*7�Fb���T�B<7:�V�씚Ҝ��|Ҁ��%��Q�=5j�H��x~�u��I�-��$�
E>c�gP��0�ğ4��`A"��ûS�/~��bJh��>%�:iY����8�y�9UF���^E�(�z��O��qw����r��Uf��'LBw�GS����b�d9���)����E>X�a���F�����x񐡐��������l:�֟��a9�`�j)D��@<!y��R�+�@�=�x�+|�.zz-{F�w���Y�� �D��ߑ�0.�VD�n&-��2Y��D���e�.�U�X��:�� ����FC�
e6S��!G֤�d���;S�(x�s1�x���˛��ŵa��97ݫK'\y�D0D�}Z|����a�T_1̂;�cat
H�V鳸J�ʖ2�� 8 <|���v��Img��%�p��lM�φ�kϛ��o��;�Ւ��9��!�`��G���{�OF�l�_�ٽ�����9?��7io�����!�pf�6�WB�$��Ѥ ��s'����S�$���gEJ���!�N�`<�4���xe1�A���U���@�y�E=�,��5߇�e>�'��u���#ي�+��d� ��g��˲`�6���7�sg!�Q��a�k=1���Σ���n�,!1FC�K���%hO�>����9����>�:o��/���CsCBP�6��%�E�K���������!]�a0{������F��f�y�m��&�W�ݓLK߯5�}�c���o\��x>�.�&9�.s7�F������3����g�-�����ܶ��~�M���xߢ�~:0���B)��˨G�MS�����A��ϧ���=����̆� .��h�
�ޜ4�@Zi�ݍ��T�@�Q��DJy�Q�
^(iv~q���1s��o�Ӱm0o)}t��΂S���e��?��uZ�T͹���FB�*W�ʌ�]�&�� ;��)(����Y�g�3���Q|������aE�7=���w˂�����\�������L_��2��{��~�&���kr���[1��D�����N�iA0дƎks�S���ןd�E�����s̕�MY:� ��B��z��:��"�� T�b����#�5�'�����6��Ѻ��Lr{�.�1
B��$2T{���p`������}��������J�]m��Wi/22��0����J^f���ZՒ�L���sйŌРk�=��b���z�=]P52ߠ�Cq����ei>�q)T�4�jJ��-iq@Y�WJ �$�1�o@Dʢ``z���>�=Zpږ�?�_;{E��J�OEO��u�<�����!�ͩ�8�-�p�x>�����"Qt�h:��F6�m���5�u�x�g�]�(��kw,�Y���m�
�6��r���%¬n�7l�q��s�R�\3l���|�*�J�f�1�Oe�u(e߷��Cv�0l*	��Z��K��L�ctG��
��5�6u&����J�!��u���@HBq$T�@	=�1��K�Nb��,�d��V	�(�.����v�}�0+p��:HYt��!��C+ƀ<�19i��1�#_��O�r�V,t�ja�#�)��0 `��hެ�pI�#��Є�.���Т)?]��m�|Z��z&�\x�y��	��Z��J�ο�����W&�5��f� �vt� LZ�9�u�CD
�^��>o�C�Lzg���L���A�x��s��aVq��:!�dPp��aډ��߳R��F���p�3zr6#d!��F�m����x{ծ�e�V0�B�|7��'q���r4�Q�y�V+�G,�$���	���'I;��`04uh坒/U��J1s������K���<Ϟ�K��#X���O�OI����� �]d^���-���9�%sBlR����4wDP�FLx����^/�C)���{9YZ���kV�_7E�D8�D�D*���-O�$f�@�s�;M�;�SW�oX
��B�� �=�����KL,�;*��Ӝ�2?����Va��2>�C_gz���ɩWX����\�5eӛ�B�s0\B�g]�	�\È���*�-zK��^� ���
�E�31�W1>}��bK�P$z'��PIH�7����_�I�Hʳ�+����uv�T���ǭC�[�%���J�8�:5�%�������^��� ����!�FO6�v�,�7�#�K��0��.�w�7�.~け3U���������^�'j�$���ͯ��[]��I��i0��Uo�]JN[�C_]�~Ѵ�H�x��!�����X�	B��l�,s*����,�v}[���ݼ�(��6�8�&��D�|!5��Ho����H!��Þ��v�6j(T�貿�p��-� �kJ�v�}��u;�����І4��+���1N�L	�L�<Ǭ~JYS�"�_�:���-�r�;1>��MU��T��wV{)�sl�t)P24����5��b��[��fc�_�{x��#(w��D��>o#���O�S��w��EJ�]S�]=!Ұ<Y���Iֶ_�˦��J�v�)Y�U��ߴ3lm���7a����t���@���N�K��T����\1 ��ް�zJ�Z�(
8B�ÌYƴS%
�Y^<0���m��y���e��&��ڦ٧�1I=�j͛�y�v����W�q��G��`�Ѐ��'��$
�`�ܺZ��{����5o�q�[`���8��b}j�s=`^wJ�7�ZMO�,l�Q���2�w�C�>'�(��q��#X�%�iIy�t#�c��g�NsYkp�����t�p:�zt*"���((Z�Z�\
�q�%�ڑsN������m�~Q��fU٨���F�����"�}�f^ާv���	���YoYߚ�c�����Ts���'k�;���>�w}�1;���I�>���;V�]�Ss$E*C�]�7�MhZE�rс�2 ���b�WԖ�#+�L��*;&�V9�y�Dv��O[ݫ�:q`���ڞ�}�xY���/אBe�H����c�l�AM�?�VF/P�ďm�t���m���
^��ڴ�A����4��� :͂l)�J�k��}�Za,�
[Ĵ+������G��J3�!m���<��Ư[����3k6��+xMV�����"����G�Eށג�&.J� l���K�����%}�$�>ٲ��%�#p!Gո*�$F��(��D��	�J�33<օ_物�K�O�+`e>e��zc�7�L\i��Y����y@�H�Mc{;8�0���pHm�ٽ���/j��K�T%if��T"e4���,�pJ��F�<l^D�6���1���:���C�_w�(/}���C]�{�\�������&2���+�챸�Eq�;����Vf��"�
�~d�L,��h9ι'�k5��^�DF���l��pl7�U�MrS������F�V��Kpԣ[µ��������,��J�9��5��4e	�N���;��"_�ͅ��] |o0xc>Y���R�Sۢ������k�����֖(p��@��˒�4��!b��)��#Tm�]J�eP���T^�wU�	̸uA����WW(��;����y�g�o[U;N���E~rd�{�T��X"2-K�4^��d��v���ۭ�&ÿ��׶�p8��V����+3a��|���\Rx,<�썍9�֍XS�Wb��1&��U��d���"�ff�r���:Y���g��7��@�KO'ѽ��Ivm8e�o��2w7>�x�拂��^�%���1An��s��uaK��D�#���G���Z��+]�[v ���ߏ
� {�&:�G8�9M�{e�h �m�č�cȲx�����K� ��UL�f��5{��O��p�(\��SA�P)0�u�hF�W����� ��.-]@�aT�2�%o�zD@/�1k�{Y���m]�6���fi��Yv"'�fq�`'Nd��*?�/f�fg�G�N�㋆Z���$7u������Sa-�4�P*>|q3��S�Z1D�wڦ�*)�"��5�̜0ٽ� �Y� ��j��@���k&@�4o����1�B 0��� �S��Ph��2�<s�l*�zk�{�\;�B��b����'�+r[W��&U�V��ٳj�K�~I�S�(�A;��[�V�t���zFt��4F�t�x� j�P$"�.�5�L���B*'gC�,�����J?N�db[D8����x�7H��58���#�1LNy����!nļ^}
�I����"�Dٸ�,�9LGv��HF�ڋ�I`>>!�1	j�-�:pG�>5oCY���J`�Q:��R��[�3>�ڈ�`�{���fJ�l���4J-3�fQ�	d8�0: �Q6�J��5�o��_	m�no���
�(f]G5���P��va���1*`^����B����ԃ��7E�W�7$�?N(�����$�#��W�+Dc��®�g�-�zB�#�m	é�1�-��
�����wG�:��z`jm��ے�3�`��2�]����C�Fm�:�k�G6G�aˏ�s�V�+�^ĺ��_0�6�!�j71�uUX�*y �5���_[Eʺh�z�F�F_ko&�9%�Z�|���A�V�,G��Z��
~�s��c�|~3�X��F�'c����#�x+F=y`����*z%��y�Z���Fm@�uGd��r�XCn�@v��*�!A�9���O8ƭ�,0���=�
@;8��ߜߊ���p5kߌ�� ǗA�Q:j?����ā�h
,��zět�!`i��Ϭ��}�$��'6`)&XOH{�ȿ��@�ܡ-��iH�u�I!zt4UBb�g{Xðg����_{We0NCݩ�V�V-�	?�&3�;�V����1U�a�~c�&�j;��	�/���2��̀�-�ssn���'Y8
.2���1v+����m���$!��̮֧��x��	�҅����#���)8���4N���c����'"�fmb��r� �9�8j&z��Ww���S.x,;��܅�b�C�X�%O9"i%o�ÆX�"�=��zM)3פq ow���y��1tuo�V^��'Ds�U]��=��&����7ܲ�Z�7>��[Ѥd�6�[}=-ϝ&�F��L����G�X\���ר�WiC�K�kV|���L͠��S	� �7��:��ݫ��&��}7���U]��k�pd.�76�a�R�w-�R�h}�-K�U�٠&0�"�q�ݢ�2x���¤{�d��$b�L���M��xKK��U��P<�!Il���q�� �PڃY���0͎KLc�v�Z���d��|Y�`�˄�D4AYq���{v�8rגY�*L�#��v��@�_�ֳ�q�.����q��qf�� 	ʠi��xw�񔝶�x��n��>�0t�L�_ϯA�X�f4JΚН��]9r��U�1��1R>8�$A�5w��87XF��x�sQ��Э7�h��"~B�*Y���d�����'�v!�Y��#�!'l
� tma���5�Y��	Y�h���؟����b:D��ϔu�/�R�n�7	F�P�����-qfv<���
s{���s	wm!�0g��/7/F�kfh$J{��=�{��=ג̃_�����S�	z��xv��S�����)�
H�%e�48�TV���?,���
P�)��a(l˟�i�5�nfn�����_n�����ܶ���U�qs(�S�m�7s�
I]��jY�D1J�+[�l����K��M�Y�7r\h�� ��-�i=�##� ��i]ǥ�^h9x7�"�>!���k��>��I���W��v'{��5��t_k��C�X]ȁ|l�_+C��\���e��`AV�`4y���s^^�)��p>�w5�=����S8��\���$`�Z�Q���&S��V��j4���n���as�(�z�x�?k�Mj=fi�9^��a��)a�X��A�}����8'ꙟ�R�<�i+�N�䷼�0KE%)0~�]��V��BX\Ӌ��ő�mD�TS�\]�J< N3H�R�U�u#C_���x�W��UB˵�=7����-_3��
�,�+rVfO�\�Q富�~�g-�:,I�hb�`����u��tM^��ӹ��1��0"&o:���<��֦�p�էX��DG�& (�rMPC�|<�NK?F��A�F.A(��ds>.����[s�?��ϒ�n׶]_u���s�K��,�3��Y��{=��m��Ϫ��8yh�I&�Qo@���-�j�h�,������H���B�;t��PzK�8V��a���X�'�R�*B	,�J�ұ�l�GRzK�5�l\q>�͹�
�c��nC�RFFr&�L��D�h�̿��5����@�Џ���jNUy��1_U�}0����6&6]Z���X�ˍܽ�A-g������a5OȦ=�d�I��f2O�p͍�������{h��5%��s�"02����j�x{�:n��ş��p���WI��d���6�^*�6u�Y�>�D�N����z�JJ��#�0���A�M���}d�宩4Z�"�:�a�B���<��b�NnY6ݜ)S��iA�<,Z��Z�K�f�v/1�������ƃ���
��{؞7�z���t$A�zl��83��-��P.T�Q8_e�Js�{*��vk��,�lL\��,�y ���s�%�M�C����a�A04
C\"��|��ۖ_��r:�j|Yq@�����׼�{+ǻ5������{x�Buh,p �G�\	"9Z/�u&�T�@������b�M��r� �u: 6A! �K^Dr�Q���"c�b��|�$xO�Ϝn"�}Y��0��k�UC�5�C&/yiJ�)��Y��7uv�/��TF~�@�4B/���0�Nh�1�ł�5���}]�g5�#D�7�~7H�1����9���T#YV-izQ&��b�x�m��{������#9���( �X�����~�H�����҄���eD�3j7���N`��v���mU]��zKr��� �ժ����P⑑f0o�Hk���k�l���u�*��g��U{�.]��7|�m�J5��j�Fk�'��h��/�}Ia}�XA��>uj~ҬǶ��}�1Tn+ e��g���*Yb ߍ�:�غ�$��kN:�@�?:�?R���x�����~��G�6,��6����}��'�-�o�j[�P@�g��.ز�T,�EP�bg՘�}���C�g�a�D��V m�0�߇�����o�n�$�v�k/�(�Fy���+�� ˢ`�I�cC�W��:����rmt^��s�c�ȇlވDEܵ�\��&J�%P�F�L.Pe� ��j�EM4�1�?"ћ5x.7��I 5�	�p���p�y��ĥ��_3?L��'3���FA��zT������Qڱ�cc�G�Ɗ�H��9��g�����{$5%��Á�J�>q���*��B��I�y�
�{geok]��CZy� 
d"ue�(}nl�}�g8׬�hʔE������v���Qg|��s�S��Ԑ� k�f����`y��j�Jbe 4����a����D�d���6��.���"Z�<�d��Y�S�G�
a1=Yv��ߔ!P���e�m� �H�_��J��U��)}B�+1���$�"�5�B�I��H��C���5ji*�2�%O��s:U]	�;|�)�KF����/P��ze-0/m��8r{Kz}�нf!��)��_�s��TȺ����Nk�����_��2f���V�������K��3�p �|�Ŋ�f���T�x/��(��f�f&\ε0)Qa��0�]��e�0��8]�V��`�Qp��2��-���:�4$�Cq�c�����H3�0���9xz�{㢋��4�\�l_����Z���� PǶ� ��	<�CDc�R�Of��a�O�<$2'�q�v�9���'jtǑ�$N��e{�����*�1�2E�SAw�����œ�6���v1�u"�F�� 3R�z��"RHd��W�E-���K@!�L��o��Z��c����W����ۦ�2>`E�B��ۄ�����B`�C���G��D� �+������Ds�nd��(ҳZ�KC�6f��A֦� N��K���\����	�L	��
��e�12�"&��LJ�[���:����Ҧ�b}�e���!�m�O�X-��t��46#��"�8��H����U���q��<�F|���x���(�>�3׍��$�:���B�B ����Rc����$�ގ��o��8�>���+�
^.<���0է$ # �;���*�(��9Ŵ@P�6m�#{�����)V��B�N�U#
dN,�g@]4b����ҳu+�=ݸ�sfs�0��R���^��D��Z�}��T��=����=K���� �`c���&'��帑pF�ý�/�����S��l�0J�ω���\�����7?��A WU��_O3u@�B/}2���ϐ��C��%�E�N�,:,;T�/-6۽r�x���`"������E ζ�}�\�B��ј!5� t���o�|��~%�r�>��m�Ƶ���yv�'�7q\�m���^;~���.���/�X��F{&�]t��g��mO�0�
���;S�P�? [��{T�݄��{:SY�\fj0�X���ћ��vo��qULƻ�<,j��%�{ ��"0u(�"�o�Y��SU��J� Qm[�a4Y�����,� �����b}`odٗ�?��ܾ�S��^�5VL�J��e�@J��;Cci�6�G��;i��/;������{b�u��4�E�:���n<Y3�\6�rAd.�^rɇkEc���^)��?�S�!�-�j]���U(���[���oK�D�>��&0F�����<�r�NU(��_��Β�F؍�����4�t�ނ.�p�j
M�d+5�F(����P��Dv&_ ��`1*Al�3_Y���k���l4���NO0"PR.�}�P�X��j��i��O�w{�w��.�*�;�?�cq�R���Ӏ��W=%�"IZ�Z��*FV�X547� |^�V^���ZE@G��G�g�Pw���p�0v*Mf�t$T��CK�I�s�0^��x��e�ő���ąn�̻��$6���n�`I�,�{�M�09.��WT~����\�L_�C�լ]XcR�w��+y�4&]��oM+���q%��>��@Q�a+Enh�CX�.G��?g�u���E��3���qS�J9aLv�R�6���"=�����ɟ��#�Ua�=8G��/��Bz�v*�Ov+v�:�]-<:��Ԍ��*��#��1{� ��Ukv�#E��9�7�WF:��ڇ�{��g�F��^>�;�0�Ӓ�)� _A���ihBh�A��%dÛk�?���d�IItR\�{i;�^ps��=�a��g���a��6�bI���(�o����0$�}�u, ��{$����"5�w��#��Z�l ��]�r^��9�߀������1�z�8H 7�an��j��
�x8��	�a{�.�W�{�O�+�v�}&���[��A��G<�2�O��y�70��w���y��I�?1��g8�O�Ԏ��x7-x<Y�2��lt]���i g���:�Vӷ���C�����}���ɑnC����x��ִ��8��r��as�M7;� ���c%�����rd/o~��z�d������;�=����U��P�r�3 ��d{�5�e��&O	O>*bo���n��0�Ĺ@����B09�ʋ:՞^��>�r�-[|�oN��VJ]�Y���_�=FMe�C$���L��D�ASA/�߫��'��Յ��6��£�T��]h	8I�L�5��񒙐LQީ= �@�Lz®%��(����]�:e����ׯ��#���$~�!�1#�M�y]�ꑗ���.��C�l,�H�tp?/�d �Pc9~���=q팭���; �k��X1 �y��{�(-����� ��:��J	��_��3�v K�z˺�P�}hmq��[	
]�IFe��J���Vv�<��{�|���I��i,��p
���%y���d�^�ury?]3���-�{mM�H�1��&1���8�Tk�(|?�bԔ�.n���o N8��8v"��c��1����jt$ ^:��c��_���}��!��bo	t��H1�g�e#aj	�ԣ��i���-��c�� ��^&�� �0�.�쵶�Є��Z�������"��Ɵ
[����op�����-��t2�� �HHɰ�#�H�Ya�������+X��橧oYKI�G�� k,H��.)X"��I��1�a�H�ۄ^L�aq�'l�����+�g�'�Z�g������dI���-��M@�4�P���Ӫf�/�7�|�N��X�8=�]Y�UF�A��Elr�y�!��{c�#u�J �Z�\�Ό};*F5����͠F���'�Y�2`F��G�����H"S��G+��+#b7!��ޕ��	�5hS�2�.�I� �^������FN����,��ԯ���r���/r0'���E+/�1.O��E�(�/_(����牫.�����Ʉ��H_gqx@ǩ��`�?9��X�{*\ab=�������O��<�3�y�	>��l��U��2A��?�@�����oP���y�DN��$L-����(�	)��y��|O�LX�ؕ�f�s�j� c��i�4-���y~F���I��O7{��N�ma��� �W�=Od$B�=�!|��G`7�X2h��&��#�P�-\�����J��=o�'���f��$��j�_�[�N����X�ľp7iP��v3j�����5�'`��E�_9�3q�	's�J
q�D.C��hz��gm.�;i�Y"r,�#Xx��<��>�}���_��q��c��ܴ�Xl���!�b�-��o��;������� z9��_���w8a�Q���*��?Ѣ��*�!T��]�s�l���u�n ��Fa��G�̠�����s��Ȓ�{j��&�6+�	.�T��G��fj�ׯ�J*�k�V"�1P�F.���|����mMϴ#_�O�y U=,��_+8���r3,��{Z��(��S}d��]j�v�����/ ������X�:S�8e���K���(����MQs��(��W�r��g�������|�rP8D�����>��TI�_�O��Vϛl��ni����wm��cE�Ŧ5;@�Ei\����߁K-&� l �=�� ��7���#ܤ؆�2K��P8"���P!�x.,(zr`����ua=>`*�1�4��C����t4n��g}�^��}h�v_1>w3�Zs�%��d36�TO����xy�xG72-ٗ͟i�DlBG@�n�y�R'��hm��o�8���I!��y��ެ���1�}���b+�p��6���#����o���>z���,_�g���(.�t��t�l¼S]n<~���a���G��Vr����%(+fZ��KG��kz��wT!�fF)�^.Ӟ�3mv&")��`�+��1�vA�)�<�ANG�G�t]a=
a>�3���b�[�x�W+G>���n�S ���O�3�P�eݏyک1슒YM�~���m�����4 �C�_�V"�&���}] �n�h�Z���nC��t��	�_8��cp��F� ��L�?�|]�K�@�4��G�9D%�D�>�ZŮ�W!d'���NE6��H���$�%цߴ"��4i�T���r�fI���l� -�����#+���F���ь�H6���`|��g�&�J��������N{�k�0��u7O `�{{7v��*p�zһ��FG�n�� o�^Y�.�-��$�7X/�78�҂���- �\^9�.�*M?vf���"����e�$dMFW�ѯZ;��0�(�~᪤��Ń7j<Cͷ)hF^o���؋M5�B)�����4�~L��Q汉ί34���5���C@ڦ�����r]t=��A��Y���%<e�l͟��k�'~�hiB�߮�8h���]=�&�2�?�L�#���	�Ч5
J^i���k�؜�m��{�� �c2�]S/Ы�#�kh�}J�<vz��� %<0��b��!C0Z;7�ߧ�:��x�D��	%��$8F�`l�� �0v����"���|�ѐS7��T�h�V��� ��t�R��ݺ����( ��OE�(6v�ˠ;�pJKZ���m4(�c-�`��� �i5z6%1w�B`�]��c��1������\��[�l�a��Ud���\T�L-^��+t{���%n&�i�W��Q*U���yI}J�]h�!V�	�a�?#�x}�JI����J60���8����I�4�- �D_����g�^k�i!:,݂Ŗ�"	g�x�LcLf�6��J������ݙxA�a��ظ�'���SNHE�k����-Y�t��T�K�`�|��f��=��� �P��q�!7�x�l�T�����
mE��s��<:�yE�������'�e�;�����m��д�'֦��e�é�`�J��G�ȳ���sD:�#}G�ch}�k�W\�$��c�����E!N1m=�X啊 �%"sa$T���BH�Z�)��UW#r0�Q5}E�t��|�L0����[�)&���$z,Lt�z^�vl7�z��-PcK������R�_��5&�E/l #%W���*>Nen�|�k�sp�������>���	�6!���=9FI��\�e (��;]vp��|w����%��3�}��,ϔ|����5=��߇1PP~�K�ǉl�����z��x��6g+���w���'i���*��k�(�oӲ@Ybla��f��J�� ;�]<h��ܞ���jo@���_c�X��Uq��!�x�)pod��1�dDc��D���)àc#��m[}��(/8@�T_�� ��D��iS��5��ϋړؔ0�7n����4�U_D}�W� j\�j�ŏ��B*�+��fa�֗�6��+;�n��<�,�A�H��I�SZ��d+��CIV\�����;�<�@���f��\����j I~�|�e����R �x<�R������-�X��s��Q��J�=z�M�<H+�&%��IL�d�V_�F�� ��"gDA����]^��#Vl$��^_v¡�˭+B��i{���!X4�����fK>�$���}b��&��oZ�����/���I;88w����Zp��>L�'�,�`�=�d*�p�k��s����=Q��t���;na.�v6����O9z�D�A�R���"ĢǍ.��	�"�0I(n���!�Z�Fk��LZ����x��A��C�G�(����Ǝ�9w�H�������͝D�&���T��R��y�R������y'a�7L�q�Ⱦ^�Yz+�& oܠ�\~�5Z,a��!
��M�2�p��-a�z�͋�_w��h(!�>�ƽo<��1�׷p3����]�}{j���~��켼��*����VFc��.~I!��l�H̕6N�H&"M����G��x42�8�VR�*$+��H���:���RL?!�yy8�:T �i}�|���z�Z�2'��!��h�C�m�ІA�6MN��;���ȞU�I��˱��[죛��r��Ca}+*G!=[U:�l~�K�[�'!P�]��F$5&"���4��:W֮��j@���D}p�Xz"�@�e�g6�HW@���҈!�c��C�m�Ӥ/9e�8�<e#����o|�A��Q�ɍ�9�?k�@;z�y�Iͽ�\EC����{�H�&"/1#B�p�ѣ�v��eG}/"�q��v�Ӹ�cǱʈz2W��9�Jn����nO,˓|h�^w�V����E/NX>�C���hd`\OyJ�h�ЁJ�'Ɣh��T��m0�w�o��+�&��U�^Y'����;H)DF'3�l��֯�(ܠ��Z0�ɏ����JJ-�%�].E���r8�P���љuB�����w����.���&�<��-V�0��T�P�3��ʍk�x�͡���+:qh���t%��%��^��Oa�/�M��i��6�-����/�~��\w����F��da�˥-�;n��]pi�D	����j������
�[��֛����n���v�&~0,���=%��9F���Q��KV�(Wsel�Q����CellA�����*�h+�P;�3ր�����ؤKW�R�P� �!	$ ̠2�@*��X< Atusz�0��w��K�����/s�i ���M�z.]��������+�M��d���Yn�@0~?�#��e�AɄ��`w����� ��x�5b�;/1o9p�R�qj�\l�6�Kw�({pu%��vb�eO��Ռ���߻�a5!`7(8q�0o�ǆ�"���K~;c$r��L��d�Ǹ��;�?�I<�3�	Y��t��m�H�BN������K{�,��&Ɨ�g��KP��$��}�������Q���ư��
���#.n�]��w����F�\�����|��B�Ar���L��š��?z�­��J���X�9x��r�/�v&��u H��7:Ғ��jJJT���<���(5�6�\�K�9^�r���<ct|/�È??���,�[���J��I�cS8��'��
�92n{�&����C��t2,2dHF=&&T�*�
P�{�Ɨ�J�'1����?R5I�hgK`�P֤sƪ�')�c�z���K��Z�U�������U�7I���V���7-ջǸVQ&k�3�Q4�I��.�9�V��H�z�9�L�H�핚����Np�۩(C��X��柴~'�5~�D)�tJ&�v�Mw}ٙ���K;E&�!Mi_�R;�JOֿ� ���_t�&ψ($�H�o�aZS��<k)�$ZY6Yެ����'�>�!2�(I�m��WYs���>�:VF0��2�m��G���Ē�"�$#!��Ak��>t1ߖ.(��T!���̬�ϼL�g2@��rA�d�i��q7�@}�5T�^]�W�x� }���4��R���*�<�SE�+z�Y+��g�gDs5�����rj; 22ΗF�a��:�.�{Dy��v���o�>�D������Q��i�((��Q�^غ��V͙�8ĵ\;����KLo9q���
�h]�?Ur@2_�3���M�J�߼!�|���,D�Y~`r�<�7���ujI�+�[�G���<�KL�\�v��i�L�G��&t������$_�IM`�l�h�
CBT�4��i����\h�R��[�����T�o�v xH��۩'�\������@�h7���(�ph*���ƌ	3� ���ϹbP����g�!h~�S/�XJ�
{�<V�ߖ1���E.
���2�������^t<��Չ~���0ä@�Kt��Yn�	Q�ooJf�I����w�5&|��,Q'�������R�'�oo:bi�M��,�Z�t����7�'���^��T��<��3�4׷=֕����6Jt���î5�Xw��
tl�?�P��-���[v�D6p���<��?��yy!�/F$�pE�h�Gh�����H����1ȼ{)��QU���f���Y#��<��Ccgw��9�_�F���j��~#3��Z����r|�֎-�l6�8�J�ÚB��Wf�K�S@-5g[vs�*c*@�E�|o�=J���iW_S�/#�N���`iByD��[k�]� q�:��2�?��aM��xW ��hA�ր��#�*IìR�� �-yngP�I���-�9�0sv�\w�(4��lʶWѯ3�K	�fދ���]�H�D
����B�{����U�)����N�:���2A�"?���@0���>���#}��+��=	���������ؼ��"!^���Á���nX�Xa%�-	�&��qB�)�lv���"7��
?	��4�2#��	�x�P��^��KV���W9�{V�'G6��5G��%]Y�a�eb���6�M��W�Vw�qw�x�m#�~r��Hw� P9�C���D�ueQ�M�G̈́%�Hmf��:�d�Z_�i&���iz����7����/+	~��]�t5�]�N���ڑ�� *jg3������A�Ͼ��2v�S��_����=]16�84\��C�I��m��2s��)F����=R��߹��0�L:e;+l�FZM��.�rE��� ]�f1*�QLٞ��(�7 \���m���!�Hf�-����m�\XE?����q���i��"�m}[zUG.���ܓ���X^����bh�����nZ�W5��H�f�y�v֣2��Q/	��7p�t�p�4H�C�h�wV�/t��<�n�D�Z��/�-1.~;[M�ߤ1���-���=)!P��	�X.�Vm��Hӿ^�1�ӓh;�Y 9%�gs@\�=����o����5��G�8$��T�O�)����Uܖ�o���9��N^��r��,����rT�G�^�k���@�ǣ����"/xf�	�o�D�)?�Dˤ� �
����A������C,�}�)���\�`2��dB��w�#����>uZP�/l�.��C�ō�m*/��N�?x�ȀG��ŵ&Fp��s��J�e�aӢ}qϤ�3U ��p��GX���vr��I9�H	RO>�,}O�J[��>�)�6��[+x^%����W�SXK��PJ�X��m�'�(J�I}�}��_;n8D�PjncTZ�OA�p�Þ�g<�䚆��J�`�Įx7��TwJ=��ܡ�[O�l�@m��C�ք<�� -B��;{e�/.3m���Pg�q$	���������_}�@< (����/�!Q{���iՐVK�E��3[D!�"5X�7�ci~.?Ev/=�xW��&ㄦ��'q�ĝc8
�� ��u���n���S䆳Zz�uoØ��e$��!D4K-J��n�\�v�3�yt9�X�)mZ��F�7�qfV5�[�*V��/W�J�����K���c��dJ[�] ����`�#@\��ސ$��,�혽��ǰ�M�cQ��l�Zs��p�Y�+yU��q�3	��#�Z���@͘m�WF����٘���`tjT��zN�n2��u�&�
	���F������N�!��� ��e�O�8#QE=٪%�l�W�~�0vu<��Sa�;�T��1��g�h��me��wB��%ӥSb9�{ҹ������f�	!��1��Q@O���H ϫC�?���,��V��O{�f���� ͔��ť~�:|c:s�]�#6�|�V������]�(��S2�Jg��Q���Kz&%�"/0�F}M�h��7�X[ئ�i�'����N(\���SҊ��)���W������;�֩��)'[��
\�ޠ�'@��	/ba]7�y<��+Y����@���ʢ��Ǒ�|F	��.�	0=R�`9���.`"&fTN~5�T�}�U����WKzV��!�7���Zk�RW�4��\���;;���Z�?�/��_�P�չ`�\�v,�������r�5�`|#��w�(򾑰ǵ��ý��P��*�H���ð�۵�k�ľ�6�(.�!9�ׂA��Ҙ ճ�eiie��._~.��L��~���i���F朦u,x�k��C���ф���1N���[�s�$M���P �hr�F�O�v��U6�UH���=3N�H�>��P�
�j���:tL�����z�˫���(ص�w��s���v���c��9�9����i��;�LB�jfѲ>`%{��n0�&��eܳVu�����{�v�<��J*Z�W#b���%��͡4R��r�c7�`��er_��K�R�����l�t������y%[���1���4[B��C�u�#e��6�������B��Hh��X�4W�.�b�l>��3)�����{ ��In�rS{Y�C������("i�lD��Doҁ��<(��	�+����#Դ+�
:)�d[�k�aEc�K �Y~7��7&;��S�̀*��f�Q���:��y���]�u&R?��YZjE���"�P�hY�{��dǈ��[W�b�`����p�9R�z�Cd 9ΏY-újj��ܶ]�Ų��Y�(����Knֶr� ��<aP˳����iS~�ɽ��h��� �xb�;M.912�TT�t�;�!S��~��	��ߕ��Ѯ8M���|��6K���	d�C�_��uQ��6��"���e���j��F`�(y�����oODF0A��l�D6w�sB�������dlK ����>�����,���:a`v���P�SDݱ|�;�v��6�y���&�ۻ�x���%j
����?ܘ�4q�h]��F�S��٨��7-�5z-I��r�f�V�w	�u �����E�u1��1�-c����\[d1Q��"�)�լ��xbB�硣4�0��XL��?�9�����h�������^�˸%,�y�[N��A�뾄��@�X���4�~�~�ۮ\���`Z�e�b#�AX|�,���Ey�J_g}LNy7�T�z�,�Fô��c&_I�����#b<�E,��j�@�U��~=6�*�du�0���Mt	�c��?X�����~��U�;o�<�
(��[B���[Ո����^���'�t<ߟ��#)�h��������+G;�����*��M$�^�M�w�s�W��&B�e�b��g��'�O�ͻ���~K�;��Hp�Վ)0A)�P߶eU����S���Y��7kR�2��8:�����k-�Ϲ���U������M�0m�qF~��Q)Մu�z�b�X��A�=����j�ׅ���-@��(������� ���m� Y
�2%OF�U� �ã"f���BEi�Rca��'_�H����O��F)TZ��w�l0�l�*�L�x���z�/�9��D������^y)Y���π�����U���@�O�	6[�7�,������7S��)��\;9�U�e3O�y(5'h�Z$�)ܛ��e���4�$�}�YJE����Ň��f�z�Ql��-9ˋ�PeZ��[JDI
FN.��b!��8�n��h��i[���Z<j�s@���gvڟo}�S�����;��E�x�D �ٲ��S�~������֑��G�0fQKˠlF���!<A7��)_�K��S�ӿ�CӦ�Vf-�|�f^���.�V���9�KRMsf�j�ců��<�y\
����3X4Ɂg�vx���bǖ���f�U~l�J��Y%M�!���7�lf���3�V���:Q��@P2FA{��T�~c  �5!y{Gu���huZ��HT'�"� m-�
�$���g-�M�eԘuX��ל3ݒa^r@x�R�@:�k�ٓݳ��<�9�S_A+�w�3TL��Ղv�f�ȱ^�!�n]Q���y���+9lFܺb��},�C�����|,&Mc���{k� #c�XmH:��E���2�]{��o�.�����ь=B]���X���0:�������uE���p�Q�s�\h��o�Z=0��g�B�����`��&ї�f!�Tz:4�\�fB��TMjkJz��#���˼����&���i�+CR�l:� Ĉ���[��N>��yVc��pѻ~Ì��S���� -5����Y���j+�mxM����1�,�A�B��ڠ�XB��k�7�����R.�E�M8ll���R7MA��:m-�D��-�u��ɟn�Z�*!|�UL��<Lz���t�G?@1�~23�RJ9�=δ�V����g��8N�� ���G�짉|+miU�13V3���p��p�����v�?��ݗ¢#��:��z�E�X--q-��l'�Ou�Uth���kL�0�[7��������բ�]����0��wovo�9��N�q������1��������A>�wds_�����oWO�O�KOyg��S��g�.�>z(�`����d��D(E{&l�9��݅a���+�܆�w�y�%�R�j����8bl���	#nb)䋄T��Xs�p�8��7�<d<|��[y�nk[ 0!ƽ�	D�	�0���|���x��/�O���ɫ�m-�������s=�[���,�9�'�a_��4ܭ)G�9�>�3�ǠPgw�[A��z��MEBًf�pJn[!�I"�g�W�mjHS�~��5pA��������1�:���Aߗ��B�٥!M�n�!>?�:�����g��Q��^'���=�K0�5��F���eɌ��J��~y�� Ȉ��f9��b!f�'X�+,��E��f
s�y�MPƟ[9Rlry)���ia�-�K�J�SC�5�a|����4&	��'�zEhOmD����B��0ו����)Ȯ)xՙ�(*��^���WBP�O7j��� �!g���p�́w���C��i�I��F�-�6�x��p��խ����������
�P�����؍ �?��5�~�/��x�*F�6�y�8C�A���sh]��	M61�儾��@�o�9G��hg�=HDlkp�G�v<#3A;�?���l�MrEШ��q��"���1�1@���ݰ֒m-��mmPh�eEa����֏�5Z͛EQ�❮�`|Й}�iHGX���I����4*��7���ˀ�c�� ���_���)��(�TϮ�z*=���Ң�T'�ʕ�ǉNguJQ��a���U%:HYQ��;��Y�����ha�Jƫ��{(��q��yǾM��Ɠ\:�vFj���}H#����:�釰.�]+�s{��A��3�Xh\�p�V��W�Cƙ4�U�e���>���H��0��?|z�h���sX��N^N�����u�X�J�1��򔐤x��N�KbNBNY�h�������\���txjA�<ws�tZ�+J���������$��T!�*����Jz�����%��!��P�nUd����cI��+f�8t���,.F�O�4K&��U�t��@?ƥ�<�s����p�	���G;�0$�@�g��wX���$Q�&$��?%QLFW$$�m$������D��swL6�������	,��*��~ft�� /Ѵh&��E� ����?�X��I֡Aː��Q�`���2��\z��/^�Z���}����M�e��G��������.o�4�i*�Qk/UBv�N(�U����c�<)o9�WY�� ��m1X����eC�[��	��:�?8?��!q�[:�I��2�&����2���k�B�)z���9���X���)d���:��ܮ&��d�w@�U��]�oJPv���h
����8�y�����l�}����$��������� vP1 �jRI&�8�o��̜�@!b���(�4�66fb�������䘙������A�`�������i�h�M2Veccd��s�jϴ�}�9��-���]+�t����B+�5��,;�s��X���Wx52w3��JH��sg����xd�m{�!`0�O\b��C�Q��E|��m��c�<i;R
[𡙒[�%��żյ��{�["�VQ��]��z04�-z�<����;r7�8��%��[)�hI��A9�)��<��S�h��������Sʓ��%~q����Y��l��L��a��A��m�F�
[j�j���\L��K�4��Ԯ��&��n$,h�&@]���K�C�ŌI�*�Q��p���K��3�x��_S�X����	/�T��z�la	&�th���7�d����⌶�"Kw*sSΧ�50kJmh�脩��Rp2)�G3|��z�Vp��U`}��wR�h������h[T�#:���w~�aA��n��Μ�A��N�fd{����Ϳ0$ 
��7�z��7�=d�I�PMk4���T8��l�����bc.n�� ���gޒ��)���L�/"id���m���ctp�YqԘ���hj��zDv*#�-��p����|���H�i��n�� �l	�J�G�1F��c?��Ja�<z�#;u�"�(u�pD
�7��p�
�p�^�d�Z-p����!.�G����o�*)�c��
It��1L���X��G� ª�.�{P'��ǝ�n]WL���Sw4o^�}	���H9��ѠUV�1>�٘#�����̕jUkK��9	��-#�nP��������rI���2��rx�w�G<Jw��t�l��$+�	9������:~���C�4@�����6� ȦH��f�^�3B�Ez9�p^EˣxJ��[xpW���K17�v��-s�bgcˁ[+O����s�F��o�s��}GU2�ˏ���lHz��>�̝Y)W*�Da�m��NI���%U�P����w?D��<�	���i� JQKdAg�vQIl��m�����a��Pi�Ik^􊑰���V�u��`�}~����*�I5�[�n�SatC�CQ	�:q |�`����,a��*:n��5����]ظ�����w8IZe)&����p��I_]��*����8}X".io.�Q��G��4��OuĨ�Đj�~�L��:���K��f�y�Ha��X�M��M<�j��K��o���1AZ��=נ�Z�_:OI%����6�)���m."�&h��h�Ho�p@*_����h�+u&�ۧ��/	������M�v�tՐ#�1�����\�;����cىP��V��2-i����zl������Q�x�~�s�f�>�N