��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��� ���/M�������Lӓ�_���X�ʌ�k�db�0sʏ��,��Y}�"E���u���W�v��0�~n��э'aԠ���{RT���N�o˫����X��*������(%6G��u�O�����^=�vn(��	Zz�j�s�2�Oj� �S���Q���Qy�A;�/|YtB�C���6������o]���גR�f����Ҽ:�j7P�ۿ�f�2��zq���4<KK8���M�E�ƾ� ��*��B.@8u���#]�(r,�}֮�:s��퍳��ե��XH��l(#�l^5����'�� ��lYB�;gt)����ƭ��]���m]7D'T/'������`�u�Bb΃I<�ϚX�C���Lz��}oߙ����K����AɀM	7sA�i�sl��3�:+���i����SJU�M�_\�����Q2��Ȱڹ��<�Z�E��9�,��G�I�Bѥ$l���lBx�)Ԅ�A�U��?���Z;��&0]��_��7
Ze[��Yf�	�������q�Թ�3�p��n��9���n���__��v=���*h|��@��D�#=���'\Ajb@���1��?11.��*H�S�s[Z�h���*Z4&S,��K53���y�6�@��9u�����r�Rmes��J7y-�J���d�v�W��%=9/�h���[�`V�+Gs�Wj6���ZS��D�h�+ov�yXx,^ I�.�b�$>�MѶA���. �}������zؾ��3t��;uf��!c�_*ك?�M��F�L�}2�g�p�ʸ�፻�ա��#���o1r�Eit�.��-�GI����8�l\�?е�jur�d��pA��m��!��z�N,���("&?�:h��J;l���c#7W@y���ϲ���P��sD�8�Q-=�Q��G�(9]���ǐ�/��EN��^>����#���WOq}W^��li����bM�|���ߜl=9�_+�_ʐ\[I��M��`$'�J��L2&�`iI��0V?A)�P!��{�	ٱL��][��k.����Nn�P�G�Dx�USG�gҶ��G�㠦-f��E�_�R�l��	H��_�ɳ�0 ���������tf���T��:hZ��'9�o��bƧ�8�aek�ž*�i��G�0����fq�ք)l��3w27�P}ظ9�}L|V�ˁPIO���� 4*�y����UY�1p'��0Ư*�
�� �G��5!?\9�P�#�f��"]�D�ua�lyB)�Mj��)k�L ;槁S4,y(R�i@$W?�&�[QIG d�%O���ux���m��Y�[�V���Q)jD1nQ���;K�,N��T\�.�!a������[��ظ1;5�6�0�e�6v���~�ogW����~Z0���� ��h�
y���_��v�v'��S�?	�x�J:�"���*Km�3���(Wy��Ŧ��M�N�b"m�]`��;���`;"V�(W����	�RahC��Z�&a��{�*�M	)"��18k'�/Y1o͕���c��*�P(s��5�޷����{��L�`�Α�����p�M����]*ưi, ���y��A���LS�'���Hf�t1N� �뚼#x��kRˑ�4��a�+۪��r��S��+�r���	�;�s5ɇ�x1�Ȏ���{& Oťv�
���7<'G�om���.�L�l�<�33����s�'��g��kVO���w�OS�T������*�!?uz����iZ�G��ӛ�_ú��Y^�2/ϔѡHꛜ܌�fܹc;tw���+��+c����(��3���d�z�OG�u��e�����D��0�:rʙ�N���y��flp���Єi�( n��c&�E�Ex0���W^���O�ܩ��B�,�3���3��ᓶ��	݉ƒ�%�jJLmk਩�r�gP�ٶ�K	��"-�(���:S�<��WTp�����n���������E���AT��'�z�(,�JA��[J���nŅ1������|;�EH�!��D���mH$��<`-7�����D���دoě�f��t�7�5\댪�%����S^����4�_�w�a�L�\c|4vs����ve����
X��p��q����8	�8u����zĈ���l�U/��!��_w�ҾV� -��g�V<.���h��x��������S�PHj]��`�d���f�l{xw�%��`�q/Och?(���{�x0g<�|��Z�@_�^4�^���ej$QL�@n>��R�d|Im�~�y�4F~T�3�kՎ��*�T���;>s�3ðe�&!�_����C4?E�����b��q)�>߂���!A���g�׀U�Y ��`���~O.�	�e6^������1�O'#��8�P�A��Q��uX�T~�����k�[`@���"f�VP�&p��h��s����a��,��d^Lf��_,��L�����`�,v�R��sX��=펢����7�-�
ӥȁI�.ֹ�q��_#�J�f����ʴ�z�X�l��毖�kk��B���(����ZUЄ-mn�w��d�� ��B�+p���b'�F���G�7��ېf!�%�l� �s`sru5fh¥�Rb<{Uv�<��{'c���bW<�s�����35Li�M-*�E�]��U�	t�lg[v�~ʗ��+�S�xaX�5Y�"���aH���:W�ZCvT#U>�b�Gջ�mD�>����?$�UbF&�3�K���c<�޶�i��2�lXL�Y#�M�IҦ|#�|��t%?�t�_�f�l�	�:#G����9?Y4$�	VZ2O��/�+������_�/��y��;�)O+;�ֱ�S4���ߦh�n�2������Y��uw6��O���m�{��O;�䉄]�-�b��Uj�މz�MK��ޙd����A�G��(�ڥrs�'���0�������x���3�2f�|�|������M�Ω��b
�p�F9��Q��N�w2�V���j+q읲�w^O���I4��ZB�,��!> �c,�X�く\�&��Z61LQz$�k��#f+��t�)�h��O� -�s�T���I�.)?ĝ��${�9�Z���)��B�YCl��!f��O\�u<f=�Hn�H�. ���C��4E�`����om�-NT����1 `"h�k�+7�=����\zzɂ��B�U��L[�Z�Nvg����Q��/� ��Aڝ�j����$�_��`���r�:���!���N���d=�+H��Q��ܭJ$�-���MRξ���#]��^9G]���nYaQxJ����_!���@�V�Ob�U��{�+<r��+�k)� ,X�1�\B�Diؑ�����33
��������Ǻ���]������x^��(�gO�?��[*h��}�95�O�S85�R��W�V^����?Uƶ����g���O�;7�p�;�e��J6+~�qY�/�v� �o+��I���H{AD���V�]B5f)tΞ?E]�5_�����#��2�c.�y;Q�W}��/u��V�=�se�]��7�	7p(���&防�`����4�)��u��t�p�ȫ���r�̓�ox)��1����V����3�B�.n��i��v$��E\zkQ�ٹ:�M!��7=Ͷ�h I�P`|���J�.N׫Gke�Vc���݄dlT�5በ����R��0����|��X��Ә�N����ֹB���}��,r��x�Xm�p�х��䦬(��q�2Q�1P`1� ��h�]�|究H ��I�D��K�2?c+�K�ǑxZ��N�V�H]�]f� ��،;��me)�L���H���� 
I�b��y'���
�imq����ZB��62C�PS��M���ƥ2��]�#bW��q�t�0й���"�Z%�O� `���ұ�.���-��Ab"�c�9� [nǆ�,3��&��νľ�Y�	?~v�,�W���C�C/�-'n�b�����dY�1���6�[ߝ��"}��2_�d2� ܁���������-���ԚL�c�\^in�ڗ[��0?zC\�3 69��
��+��a�Y;�a�>vzV� ;%j���w�Vd�.^��7a�}	��2?��ݥ�Kd`
�o�����4G�n�j��D��h���w�[��W���oF٠	��ܷ��'��[����Ӿ� []�S�Yjrp�#��h�{"�&K	bGH�?���� |�n2�jS0�M�jC�?���7��n'5�Tҡ��wqk�g�}l�'�^�2d�3�45�M�k[ZH/5�C��@$jt:����*AY��Щ�+yX���vt>$xV������Lb�*�#�l:�z2|���.$���5U>a���������_��*��r���e�G�L�sR����֦C��Q��͘�$ ~�8s>�)�A��f�4�[����ڽ�<�&3!@k�xSU�M�ڑ��K�H�`,O�%3|��(��>f�p�'TK�-��H�6���]
�&��9�v���ͱa��A0�I�� a��U��Gh�v38����w���x����������ӾV��F,�?�uM*�Jg.uA��aE�F�����x9Y�'��pmz�A�0Yc���*v�� ��*�I�S��W��{��QX��

��/9n��� �E�qYa�SyKڡ��np�G�AkN����6d�&XrI������o{�.�.S@B*O�s���p]�=n��o��H�~��Oh	\G$�OoP�������Q�^���>�
:'��۝�JB�i�L6;�E�kͿ
eB���F@��y �R@C�H�訓,I|�%���7J&��v���E����r�Z�E���%��8�9z�Ր}���owS�G;E�����$�9o](6Hn���s3\O쌒���0��!*+E����^
��n㽕�Q�/K��EE�p��� ��F���J\�0��7v^O�YLdP^�)�4�v�"�0]��ׇD�*�s_���iV�a'-���j�1�3�gg&gai]�A�؞_��PMK���X���97�&�Ko@A�*[�<�4h���m����>�~�i���~R�7Y�	䕖t	n�O��.�Y�2ߵ�*W���f8� )����/��8��cMB�.%����4��t-1�w�v�=��pbH��|�r��JC��5�6�
0��\?��N�N�^L�U�Qm�F+��(C���y�l>��y�R{�|�as�QW�4E��s�ڧ�Bo�_
�B\��W	G'��M��V�I�\;r����9W��[�M	�F�sC3
 �<��:�m��>��J�i���;hy�P��A�3�P��f@��@V���k��yg+G-"�/��8�|0$�s=�]�~�d#V�Wi�xLd�צW�[��":\�J�/_{�!y3:-ib�2܁{�-�ڍr�ޛ��@2ː��zG¦������k�AM�Zx����Ɩ������<��²��Juvq��~қ-����l*ϒ'&���@i�.�N�>�͐Fg���+S��v:C������,�/ht/�"��r/�>��@�P�SjGjt�1�|vf8�=!,+�48B��Y��+?���Ū���v�����f��.�LL����eVH'x{6a@$������}q����uς-�!�C�h﫳^##�|� 7� Ȕa�!i8<\��
�*�����u*��V3Q�n
�����_LH[W�V���f�~�Z�7K(�q��B��E���/�w����*�J�Pެ�A��\��>a�~��i��3�P�
[
n��G��_l2d(�(�,ĕ~�ɵ�);,ª�l��.f�Hsk��7h�w�i�ϙ$t|w�9�2>���}ʈ�lԠ��˿�+�F$lF��0AN�@kwh�?^:�;`Zu�O7,�F��3ڀqX ��+2������7�|?���v3���F��5�/Iu��,A��J�{���t�����n��� �-S��Ѿf�kOu��c�H-eRf���4��K�`�B�
,Y��y��f��a�`힝L�:�!W�
��G��#�5^~��4R���ބ�cY����E-��>Ȯ3��)��/��/���-�r��?]��y��f�Ԡu�r�3G��d�N��q���u���L|�B�S�q�D�Q)�O�c�u�G�f�
��s�$���@ϑwV���"ey�0\�z�m0�{��������Y@c���v$��� ϙq��xv�n��"������Y��s����%���[�`�02�*�߯�ØD�����N��˗BGj*w�\��A�#�W� R�(Ĉ����_F�y�����9�2ȿa��	�}?�u��/|��?�e ���ND�o
{q�ye�����ߞ��{�n�j׋__����|�{�2�=���5���'��Ѡ���͗ؠ��C�U���t��?l��L��+%���X�c�s5&4��O���¥H����p�+�8uL��ԥ�m�>���5�r��	��g�ё��H} v|������#.E�TH�^)����~�_
�"�����T�tK��v�G��-�!�޸����1�j� =cp�#���Le�j��
��]Zf�p<���֪�(���t���)Y�-�Y���,�?�ru+��r2`f�_I�|�6���&����@�}�x �y����٪olL����b��+�|*_ʾ> ���ګ"ڿk}
��}��E��M�3�nU*�YR�dp
h�a���̰�TM b�����-���f�7��@��%{��{LY�_����_����wW�j`~`���s�Z��n���5�^2�AN�����.����i��˼�JvP��Hc�L��5�W$N�({h�J?׹�V%�ͷzHy��>�,ސ7�#��J#��u�{��/���%�q�h�� �v�}dJ��n�m�Ad��=�<F�����'���ȅ��]�Xb�뚃���!�������+���&ð�
������`Ű�*��Ɗa���'����xP>~���qb%�}�'n�q%w�Gn�oٞl��p L{CY/�ׅ�s�
�T�*���l_��S���x q;�)owJ+��}W���i7�:WE/gV=ݧO�e�V�Gah�CA�Y����L�(k��p��]�c�ˉ��-�-�7�N��l��Z����x[�����jw�&�s�",�\ǽXCc�z��9_���oy_��CZ5�.�d�16C�Kyk��yx����fq�7����t�O���VsW���{� �2��ݡxπУ]O���Jr��%���t3��ͅv��t��f�Iu��a���Z1�/.�;̤�K'�� ډ76T��$p/����u�J�	�e��`�$�vf�I(�Z�4���id����@��Ρջ���*Z��{F��~��{���Y��ɟ)m�vɕV������`�W�㌼anO��NӮn�)�gV��^}�i�
����J�%x�����:ꐎ�P�/��*O�M��c���lQ���m�B�A�M+s�{6A�mk�&L7��,:="��7�^T��B�r�_s�HGD����:|��?hʞ>-�v���p�����;sT�P{�k�����p�+]J{u�q�/���x!u6�d]jJE�9V�ȩ@�-%`nwA��}[и�Lh\�hD�Y�#�/�X�&��d�P�WY*V
��3Ԧ�:�ИG�3�ܑ���Axe|�?B�>�R�@�7kW�s3��֎M��h0:����d����j	�L6�}�¢3���In���J9��l�0��ܥ"��ڶ��3�q1F�n%j�rSS5�.�Z�YT����Y�{$�	�܄e ���Ca�ňS���S������I��S���h�3����gMa2[�}Eibv�͹�u~O�^�r����F8t@{"��T��_|�`�� s��4����FdLή��z�٨y"�w�&H�BP��,.ǲpZ\d��n��E���t��P@�_1�pG�ŗaX�5/�?�yi]���X���)�U���v�͢>(��
�#b�ƫ��(���%�8�]�{Ra:��o	��z�1.�s�"���G��Y1u��^�hm�{LxdW��M%c�p�Ӿ�,Z&�hx,��l}�f4o�ےC��k02ܙ��"to3�n�S�+%"��]���'������$��a��Y�Rt��0����TQ1Ӝ}
�uH��TIgn�/�A����ک����Y��,�ek$]���sq�-�,i�����6�m�(��,��I����C89˽~p ;Ot��P�������W܇�}:�t;������f�LKC�ℓժ�X��9���3�;d��P.0Ӂ�H6T�)T��͋M�<DZ�m����N��I�R#�i��Z��)��+�݋5�Ae�<������Y���9����U�\�%� ��0��@��8�,�)M;g��f���1���?x�1m�\��N�/v`X^�r��X��e,��Zk�%��8K-�Z])f����8yŦ;��P�)�gQ�B=�*d��6�������o��j�1�VyqЌ$�]�Y�
�?���5��(���?z�e ��檟��z�u�`~���{�yrK3P~�'��6�ߥk��7P� X�F2��5	'"�w �u�du��}A?WEyU�V��Q�j�C=� ;׀�Y�������{ 9�a�3Ġbx�ȥ��M��C7x�4l�����ܿ�k���â�wb��J�AD���i�!�����b��&آ:o����6�a-�8�
�װ�ᦦ|u��$��[��jv�j ���1���g�9m�_�弣w9 ����*6q[0"�ah��ǃ	T�o�����h�?X� �v��N��W{���.j���N6H�7��b�U��x�dN���]
��	EM^#$�$�����mT�۔g��$���;1	��,�;"��(��"�
��K&�_q�b���5ҼW�+��Fx͝������9��͓�K}�Fٜ"���萫�D�vt�",�6N�jV|U�W������d�1iW�T��d����K�~LA��R�i<�p����xWl7�ȤJ֙�܅Ū�	��I ʊ0��n�kb+g�
��4q8U�"m,�϶��K �"]����:lV*F/�gWq�{wb��e����ϖ�x��L<��d4W��&5��B��ݸ���~X�4Ŏq�y��3@�c�z:��B�>�\�������T��~�V����~�s�Ξ�[�n�6��ȳ����>F-���D� ^��D�{Ht�quAV��y��	˭Kvc�5�H�L? <f�E�VO���-��d4���,��>�̢t.A�������*���:R����	q�"d??��:H��ث�D�JVD1��}�(c���@�qR��~�Ҧe��ӥ��N�0{4�R�#f�v�,�3҈i��{��4�lk�0>���ۆ-�)����N?R�k�O��t��Q��%��A��x����@ǽY����s�4��X�������$�D$�Ĥ/ln������_ƥX�M �_o��jCS5�$�SC�.�W!��3��3��\DB��m�g�Bb�=4�KU�g"Ic�;3K��d���|:� ,�E�7�r�ɅXԿ7t�]��ny��2;�6��5z~b[Ǧ� ��y�@���;�`s�`�Kܣ��d��i�iZ����Qg�7c��E�̓4M�<XKo�5M�v�s�؎du~3���"�T�,!����,�����?�>e�l�|��(�e�F��;l�����	M����pF�숧/,FXu�	M�	�g$��,.y�7�&F�2��dY?��PO�3!ls}2vW��ݛ�5��e�`�ۡ��ʃ\���L4��Fɤn@��ڛ��pKnx������ᓎ=�J۷��$���}���N)N>z��Q�p��ӈ�:�l�ئ��F7xov1�_�/�D���r�@�mN:�Iɯ,ȶ��T�G�M,h?\�r�& �%&���N���ԳA�wȴ*K��88]>��v\w��'O���c	�x�nB[WÊ����g�.v�4�Xi<�M���+O���JO�-Ҷ�����r��=�UD9�K	MV�j��|�>�!#H�V�7v=/\2��ޱo���1���L��, 3\>a&�׵9(�E:[�HPs��$��PZ+���	Qp��/,����S����l:����ܰ֠z������"�ie�&���g"�C��3�]�!�r��o�������~u�
4��i2�0��X� ��5jU����}:,i����Ԝ��dv���jgx��XrgG=`�_M��������$��[�+%�y�(P������(fmǴn /Z��vm��?����Z`�.q'�F�+�����]9.�%���(!��|J�v�pǺ's���p�{9¢�C�8��W�\	3X����) `�H��wo�4����Z�)�u�^���?���X��YyR*2Υx�9����氆Z��;���P�
�T�����dh�V^b�?���� >�r�#�C
�y�x�-�'o�n_8W%'�y.��S���ec�g;>_K����`�C����L!�$B��u2�U������!I*z���
���b(����;��1;�[D�� #��|����6쯞��K�{�b �����>K��������_�},�D�EБ�n��ӵ��~��	��P��[���(����~�c�P���SV$ׄ.�>7=w��F�MG��#-��1	M����x��U<�����]�'ӌv�+'~I�ͫW!�6�`��T�����	�ґ~h�vߞ��u� `��s1��t)]���@�{S����tZ��ǡ:J���n�� 쇆e�oD�W�P��nP}i�=�����*|o����r�l��@����)���JUP� dd-Ljvc�j��� Y��|�s�����qu�y5�-��� ;�*ul�ǖ�I�Y��&C#��3���X�-�`�����{9BՖ�j�z�m+d	�4���~��_�qK�i.eoO�^_'Ǐ�;�b�~ ����Q�'���}K��O�K�T���5�o�ِ�6�#�i	�+3ݲ��*��?�|�] Wu��V��� ��!��T���ϺEl���}j�)��`�m>`x�bB���D}=p��7ˮ����77u��l���������^��G ���_*��" ����"��d���4��ϋ�3�5�t��|�A�­@3E"<��ʙ�[���7���J*\ꩆU�#��n'�6$�J��,�>�Φ�m)�A�%I��l��k��QJ�' $&̧�B9[�����L�L#��'���wF7�S���cK�a?ZwM�[Qݏ���=��1,��{�Xf��C���[��9An���k$�_'3~F"!�$���'w'��^�3��"�H0�'��oF8ٿ?�j?�	<2���ɀ�V�EE�C� G��Mz:���;D\ܥl�0Ot��@��F�td�"�f�����_o~ͽȻ.��������U���ow��iV����FiԦ�L��	��=��6�F�峑W/�ɍ<�W8�\�˫!8�fKw(ߵ��s���?���e�,�~���1>A��Futw�̎^�G�L��)�X���P*���;ɂVÖ`��lɍ	&���R_��y���|O��\����R��Qζ)�j�c/��|���Y	���<�j#W����C��M��I����|w{�	�e�fʹ�,�\��ZGl��K��zS��6�D${��>,�->��)U��l���䁞d�wQ�J�������Fb�F#� x�B�ǡ5��8�O�z$J�`w�F���Ĳ����3�����z0�-3R�E`f�h&Y��R�`W(�@�a?�������?Չ,8�Ѻ-PE�L�\'�ǎ�
'�Y��P��t[6�n���p;|�ɾ��R�&Aɬ��D�v��'<�m��ɠPi������q���(*ح��qy�K���Qӥ#��T�ʼ.�2J�һY7��1-Jp�2��ق�;��#�^�ǼN"i;Ͳ��G@�ѓ-���,���0hE��v��:��^�˱���]ܽ��q�Tښ�� �J���O�5��/Lb�l�f�]��ꏠ��Y�+��n�)�[?�`~��Y�c��w,M��Xr:��A���m��f���@G)u`?*���ѽS�QY=�`Xϡ�q�G��l�����R旯'�c��{���[<+q)Ij=��c�s7����� �)� ���䗪�y��&�D���Y��T��\h8�ވ>�˂�|a�9�G��C%r"������F�5�S�`�r��{�( 6?�z^㡔<�����@5�����wp��O�:�L8�%���|v�Me@�2N�<,:�t��� *R+���X�&+���t�F���X^�E�1��!,������r����R#���E�um��w��^�J�%#��q{|/�Ή��&A*�cnM��i��u�W<F:��X*/ǁ���y����ڇ��$jK�w�L�� ��&>݅�xʈ�"�!.+f�&�x�k�=�2������@���E���1A��0��'if0��3W��o|��;מ�1����F/M���m�$������(Y��0��n���|D\T���]�)����
`�-�]e�t?�Ԟ\׉��t�	N(��}��*'M�
���A�Mn���,�8�E1�����-�bO�ٟ��5����52� f�{ӢBI�(��iU�3�<2����,m�60.˧�N��L������!�\F��B/��HuGwV���P^+MM�qD�Zrh��s?�,����czm�~��I VRI����wyLk�����TQ���J����k;��g�k��ɕ��^1���^��l��t���*!�_���.�U�%���tn.g������g�Y��Z�F���#�2H3�^�ۊ��]����!���7����[]��J�ctjRYd�b����/�@�V4:%R�T++��d�(�.q	��8{�jה� 4M!!�+�9ϼ[v�H��H�=,�1o]%���ju�3��*��� ��5!9LJ�". a�_�
��[]���o_my�A�]�J5b:��o9�y���K�yi�sg���3�+a��'d���~���6Gx	I�b���T�̯*W�+�գX�}=��%ξ��Ր�}��L�݃mtӑ�u��{����a�z�`D8��rx�#L.�	3{ ��3`�>{�1��Hs:��?:T�&
8@\[ݳ/1Ԡu>?�M�>0�h����_r���s_�#��.t>�<��5)�Dw*���KoW �Z<O��KÎ�yz���`���J�'BP�/( ��f��D [�2��}r���U��۴Y��Fek��kb@��(\�o�����,(\ɗGؙr$��3��^!�΀(����$���Ew�6m N§�dÅ��񕣖�I3B0N�I���J��	2l݁#!l�T���p3|=;"DB?��U4�0;HL"E\<5�g\+�B�,:�>�St�bD\7�� E���]��{��Qχw��"��m:]����o�JLP�A��󙫖��A��ޑ�j<�&�i�h�zWvC*���,�ȬU?�)�o�Ic �(�� 'GWP�B��Z�n̂�3��LzZ�٪�ؑ�n�_�:L}XuV/O9�V�y>lԨ�=�KR'g��x޼��(te��k�3�wd�G5(��9��?��ceT?@��-r��}`ŗqr_y��>YV�@������{�l���!�Q�o�e�@�1�����;:C���^7�'Ǘ@��>!T8��!Wd|�2�!��En���ۣ/�G�Q�TG4��1��Nn��2}��E21|��|���7ڎ	t�6�2V ��q@� ��^�
��w����>�6��E9a�`��	v0@u\��`�K������x#��kh�dIao]�R����OX�����U�3�1���ȴ�ԛ�[/��D}"d�N/`������/�Ly_��Z ��m�[K�|���A�<�&���$��)=�]S_���뚰h		tD�W��%ŉ[��	�t���xl���s(��M�L��q�2cIz�ӄ�Է�C�5��w:��t�6z�Y/;��.�F�Q��E��t�ꂅoi�=B]���a��IK�&Sg<2.Q8���eh�s�=wzm���e��v'�Tu�a��cΈ�"����,�>�ٲ�Y����-=ȧVC�ε���Sn����;Ὦ�O?�&�^�J"kux��u��zF/CعL��5����]��W0��vߋ�Łem��w�=�
On_�M�e����)R�e��m[[-�M�kF*����/�R��HE+)�6��ŷz�9�Uh��>�֛_�s`2��$8�+�>�ĲU��.��n��A�ʹ�[&��u�}�`���m�)#�T>c��A/)@��9c�C��C��Wyޝ�#;I�=D:�p���F��Eɋ���'��N�w�:����j�ޔӜPd��b� ���5�{Q���o�~����	C����^9�D]��K�Z���\(#�u�6��DN>�@d�REZ�^s��E{KF��Op�:��k�n!���P��)Y��|���P�c��W~6� �ɶ���������[
���*�ͪC�@��tMj��`�����Nae���"��J��)��'q�<�+,uԢeە#P�h�+~���(�H��4]63\�
�C��P�6�槏_�PYbe	ݒ�4���_.<��/����Si�<�	��Z���}W.JU$ǨH�����T����A�<\3���;�:OBO4�`n��g�v��Ԋ���e��v1���ڤ�(�a����g���ϘF�����єF�VC:�O��� w-���������;luM��0Dx?<�Z�3e�	'��[�}=���r�ԛ�h\��ח��v�D���r*��p��5�yy�S�V��&|��~�M��`�S�C�@[��ɚ�Q��F�)������դ�ѣ:���x?�� {����M�i�{KB��W��L����q6�}�+[����G/��i����~ѹa��Ж��u�݃�\�N���p�?���}�
Ë�\b/��#��z�tKs��X<@������+��#���cD�d
mC'���XΡ�ȶF�Bn#��&�_eW!������6�y�vrI�>���'�A͞�����C�՟l�7�c���'��9���+5c���c��MO��w�r���{^�e;� � ZKN-F�%�PBR�c�}�v
\�t�t����)N��l�+�&��-�5 �mF�Z�U�`�B�eֻD�K
>>���o���0ٕ�geb��W�t9b�W�uIN��3z	�ԝ!gTN5�w�Ju�es� �T ^MMQ��٠�����VO����$ QБ�[s�3H!tx�����m��?�pl�٠�a��GZ��NidQ��Y����J�Op��w�{MSO�Sa���&�4��Q�$k���ܝX�h��t�d�>�A$�n�Dĵۇ=),�V4�E�FZ3�2u��PLޒ�<س�I�4G�c!���	?���~�P@ԭ $��Eq6aPVf�����9�A*uIr���������'�US�w=�6�B7�~�q���ռ�͛y��F�&|�'K��F��-�u����lS�]Q�,+=F��-F��A6�`�=�	(@�(���[|�É���̝}�o��sK1ԝq�w�z�[+Ȼ��dn2�c/���Ej��f�o��L	!l�a��yAi��y�+n.��oGɅ�I��� 4
���O˚"��� ��}��{���V*�vx�5>v�i�D�@�* �㴴 �ܪ���������~�Wlb*�����i���M���Y�ªe��8jyހ�"��7`xȦ6��:УQ|�*V��Z�d��z"F�9�5`��.;�N��3�ކ�.Bf��|�4ͪ�L����8]3K8��3K�uTs�[E�����#V��3OI�a�7?}�� ������<��C�-�� �7?l��ؚJ��"�E�	T�%{�B�����r+J\���\5�%g})*s�c��MY�x-�t���1�	����u�K箇!�h�44�+��[�2v�'6�	I��j��RM7@g��?�D�#���-"F ���3�s8y�T����X��g1��9���Qp��YEM���ؕ������J��8D_��^Ӿ���1��.�0�vHߥ�B��[g<'n�-�����=\`��zE�|�0/�����|�Mb�^�}f�F��˽�vq:a��d��i�7�Y��0� ��������X�ɱ/�D{yN������y#c�N�/	��&�$�Ʈ;�|������6��-R�,|�f��,^�|@�0w[K0�R\8�]�31�9�ݏ���k�9�L{���2�x�3��
#/.�4ѥ�z�����S��H�o+�]d�s*oV�`Rp
�Sp]��˘��``��|I��߲'�����6�6rRm�>tU{�X��i��� �U�N8U���и���#�v�1����\�ۍ��7�%�J��}�w$����L�9Oݜ�6;�&3sSŞ�t���%�Y�SI����jr)#jF��`��H(>cKTM;q�j��|�~J�t���� �5|e���Q;tPL7|]C�!��c�����1�r��A����BG�
���X�:x�K� �y(��氯��x(�n�e�@*�^а��N2�-T�<�j�7ɽ��Z��EF�vLAT�� +<�1���3���ʶ�tX��<���t�iP@7�Ǩ�So��J��d]��_�b4\�AI��'�l���3�-��w��1�����؇f�����^�a���:��'�j\6Ҥ0pyP*R���D�vh���9����@J.z��eϦ��7���[?���g<�]'��D��O��)ø��򲳓�Y\��&M�/��1n�"j�&�GWQܟO;ɲۂ�ُ��P�3��p���~�P��&a�,t�l>2�#wl��u`��K���Ѩ�m�^ ;N�_P������,��r%}�����G�7�-�'�:���ˠ��y���/!@m��	�k���C}R�BH�X�H��OI��SɣT���R1����@��S&-�Cӷ7�'�Kv�x���N�8|��Y���_n�c��_�nq���i)�hl���v��FWm#��⹦&�c�TN��?��/�@"�w�����&� +��X��*;E�^xf��jj%%t�-�>̈́��w�BeF�	s&d� ���4��k��Ϝ��Ś���C�ޭ���
�u��$=5LeY�F]A&��.�(������(��H�}u�Sl�yeaUV���z�A}��� Fu
��d��-?c�x>��@��C� %�bU��zu�_ʦU���3��^����4�#J���M�&e��AՊ%f��7#S�HqC�faQ� ��+�Nk�P���@*�RfY>��$c���?t��]L4�N�&8}CU� u�Zy�{�����.�}�*ŭv~��AOP�ni��_�+|�/D"�G�Y~�4�I.e�v.���gې�1�%���hGԄ�b�NY�]�^�j��.���b��=6�j��#f����Or&��7G��l�6n>��2x)Ɍ�
A9f[����91�;m	�l������<���t I9�t �g7�u�(�+̘]+�-� 3���yx�Ղ7~Y=�s�/_��n�}����&���t�`�-��x��R}D�ΡX%�I�=B��]2L�$��,��{|S��=�(�\�ɂC��l\�^\����O7sˮ�?�}?<�.�>8�ay��7�s<�N$H�M�L�C���Ko�4)W���ςyT'S�����x�f!N�﵄|Nԕ�V�P�'���p�&Y�rEN��KT7<��&R�+�L�ʢ �>�=��δC<�m�y��&�����O<)��(M;r�x�$7���S	�&�sȽ
8^����c��F	5r�4�A@�B�yO/�Pu���m��X��ŧ�A�H��½���A��n/'�Hct������p��tX��UX����N�7�{�w=�sҖ=�%�o��Ϫ��i���rZ���{F�y0��U&��Lq&�t쪇Va'�D�K�<S 5^����g��!�Y��S��ي7R�>j�+�Y�O�l�%ՙ�z��`S?�MŤ��OwȮpЈ�"�g�Q��pF1�5d�Q����l���FE��@7�cK�U�K�����+u�Y�?����1���Ʋ�A�[3�Le�='�2���u�����K�0��ZtN�����7�e�d~� \�w�n#Ŀ6��l�x���D�f�=Ѧ[nFQ���M�5��0V/�I�Qz���Q�wk�5����󑋻������G	��y�n	���j>&pE��O�F�T��}v��i"llY�+��<4�eD��5%�U�U=�3�=`2q�����,L�k0���/b��nl���1����RC��#��b�]��+�a\_M�<�ã�!Xֵ��%:'Y�˪��ϩ�>�������w?���Dy�>~�{Dp��<��5I�U��*�u
�Sl����&�))˶$�3
�"�%�eQ�8��ĈRm�A�~ ����8#⇝~O��� X]�ɇ��A\���|b5*	�]��N�&�«�˓/��#؜�f��!�o>�wQa+ow/�uaz��e錡A�LI��G4N� N׾��И��DEۂ��J�E��U&������{2���A�[=�2\����\�^����U�Bƻ~���_�:hh+¬'������/�x�p�KO|��M5�9��$݅YT�k�F�;q��ϸ�ʥ
��ن~�2���g��b����y_�3�rb����Ep(�u o�97 "�4���f�B��� )�	՟{��>$�.����,ׅ���)�J���;QIP���u~�C�x��4�qt�"8=��ϼ)���{V�r���V�=���4�G=H��\d{d教��/�	77㟠�3�-��)P�7����2o���I� *-V�	�I`�G�Z�bǍv��qG�m��	���v�C���>����Xhq�/_�{�}�k���
/��%LO!�E���P���+��j��,�N��*�(�v53ڱ�T��)�iZg+�$`kC+K` ������M��@|&�v��+��q�jQ�b����E(�Fl3����b	{G,$b>�$�%�b�<�B`?���zE�Р���"cВM�á�,��`�"x�j�À�o��Jq��q_���\�4�br����8iC�u����N� �5�������y܃p-�(��{u��f�Q���Uo�KrH(�(Xb@��x�S:0�6\opձZ��dz���A|�6O�
��5��Y���V �<��m�� ����%����dE[�����R�����	L3�3��Wo��2����uMq{�)(Ċw�Y�F��ǖ3�8�I?پ� F�\��0��R��0[�Y�T�}`����޲�~v��f06�C�v�ʷ,bW5Z�n_^�_�5�B3�ԑjX���9����F�B�Y٨��&��i�ӽ�^�R�^Y�bq��Å.u||�DFP�Ub� �p/�)�>d���v
�B#�c��>�'k��[0t����j&���Q��at����cr#���򐞖0�t�O�,n�1�p#~38i?cxN����Z�^u?�Y z��ө��"w��R����I��3�����L��@ֽ�w�n�L�.a푣[�7�Kl�n����`�Z學�9N��vv q-A��.��A��3�s��cb2���sߤ�Ly5�殳���wkyIPܧ� P�;��_Э3䵹�bs����[�3+���]0oڵD�$Z8�ɼ��3�x54W
-b��YM�VbI&�Wc�g*��ֿw�Ț�緶���o ��M�*�bo���jw�G2��=:�cuC�����_�`�t����2Gv�>�L�c7���&��������{4'K��� ��ta�$��}�Y���k�e&�ո��5�D`Չ\&�(�^�~��X������wsVErr�s�;|�ˑY�6{*��d.;Y�,��Oq�����	�ҚK*�Ԧ+4�#��)�/v�k�m�Q�Ûf�sI9]�+�j2;U��[�v�H�y�hR�,d*��:~�nҧ��.򒦅��N������t�ѤF.)�qk����e��d0�3����9�����!;�q�kz��jA���kn$�A�������<�n֕� �-� %�͘���NgԒN�Z>������:@G�]{������?��x�ϫ���3�Ky�3�����V�?Lf\��o{`&��	Uv�&i
ja���������V1�[j��>¦����!ka�@����1�O! ��N?v��캌FqD�k�+�������h�m�@�5B�uv�	���Ԍ��2��4���8��5���cf��K�|t)F�w��t�6]%�eW5k���DA~	I\�˥��i�&��!��w.]���Ђ��M9w���<�<7虑,���5�3���6�A����B��~�&_Gn����۸���]��cq�ӹcW`"�?�ɤ��E����H��bj��.���i\ո����[k��+JOl��*5�|@|t�f����F�E�z��Z�`�����-�
uA����*]�͋�����G_���+a"J�(�bne9�s]�A�ܸb�'��ZA��f�xCW�Q�B�x5�¬�ٔ�YL���l�-ǎ�QOZAʕL�R��Q����)X��-�q����43��2s��%z0oW/%�Е�"N�n�Q��?���Y��M�*&��a���w"�(h������)���^��F�S�� �Y��i�-u=sj�K��t|���
�d�Gy��'},yJ�HAq��"<�iY	)N�9H�8���(�p������.N��RR.HlOؚƋ�3���J��ؓ�tlο�s�z�c=��.H�MS�j:[���#2�]&`����
Pc�[��J��t ���<����=z+.wF;�'8�p� 0�x�b�.:=�_^g%Ѯ��o��c��88FaSܭ!P\�kl���n��(噉�<�)�#uɯg��M� &�^�b/뙯+�KG��7ʆ���]LϾRW�c���i�H��19c�h�_8�%{�ĉ��}g����\����K�!}�m-/�+�L��v���-姜����¡u� q�7��`�J��	ò�3j��ĉl�h�*p}JH�#N=��t	2�bw�2��}�=������q��e�IF�Y�F���E��y)�u������τ��A���������z,��Ũ�5���b�:�?�(!)��"����uua$к$h/b�BF�4�,r��9b����vo �Y`�Z-�ޗ1� ���]�h.�Jnzp��3G��J_��ۍ�?�vW���W����ڶW`y��k���w,��2�Dr��#��ѩ�o>I��\lHyE�ړ]�kJ~�C�x������GF�<�MS��r����olc��WNA��� b)�5�E9��,-Dg�2q�0��1^�o��P�|�?�V������#v�����h�xτ4�G�Y�>#t���]�b���v��#�j_>B��ySYl���1.�[������Gp�z��/�t�vհ���ox@VANd!~ϔ� ����<�+�՗�C��1}�D�<���Qݒ� -��i�.q����}�DZ?��/e([P�8��T���c:&�j-z��w]c���O)v���{�]�b�uA~{Z؅��[<�?�Q+\Bڃ*���qG{#op&a+΂,$�8��ֱ�L��6�H���=�����}.#�pu2����E���^y��� ̠.)JmUs���-������� �
v��e�s��Jy
�W�oD3�,��x�֎������I�g��Ѭ᪌~9/撪�9�݈�p�e��W!�'	�mUT�N 3=���+3�6R#�����x�M�Dj�BM��� ̎�¬~(Hx�!��p������[��4�Ҋe���ⰡK�}��g]A\����)R�{�8���K!ζ�w�s���m���H�����t��M�$�:�5oû�֑������u��w��>��Y���j>R����rZ~��5�PYZS�P!/50��{)�+�4�(��֘����Q�{R<��2�FN��J�wmW4%.v�H�{�&M���.��M���':�C��t�+<�%b0d!��K�9
�&��~�}��{�i��#��{&ϸq�J���h�G�!�F�F�tH��7i$�qK��6��guDq�isJ(HY��k�����I� itd
��!գ�j�M�o!ݘЯ�ɤf����օ�tdFIc R��y�����J���i��rٍ����ݧ(��(F�hM�_O[��v��u T��h��%����J�wP������33�@o1X� ��}�s�L����'���8a��q�[Y��#�`~%�E#�2��-���X2��
�O��f%�eFt����U�)���%r@�UJ��F?��>H���z;aZF�:��!���²0O�~�避�- ��)�{������17��P��U,uR���pX��qb�-%<��X�N1��_M����"�����=���%;$�j\އR����CY������X�	���K��`�(�Y+��`�b��?{7�ռ��h>m�AG *X��/���ĜWiC%�ĂmF�ʬ�?�����87�z�~��Ŵi�r�DL0K��wf��C�~�w���C�O#oP�X��NM��_Z_Ys1_�X�E$�Q�Q���鳐��q��AY[E�[oK����(`���}�$-�r!'S����
�W�V4Ik\�|/'��t�sz��C��u��a�g,���J�f��=��
���'����8�קQQ?������9��6��d1�T�Rt�������� ��B=-(.�ݹ��R��U9�T��E?���y6�I�m~����a9��TsH��)؎��b)ϱ�.^��	&#ל�< ��,ꠝ|�z�x��r��y�s�{��=/�B'$��*~�֤[ކb��3<g�q�6�,~_��5I:�m�wP��	J36r��˟Y,Q���JMs��bg�|�����9��x�f�S��vё�h�F��ߵNi߳kUmw�5�&�S�2H��g���@��-
��w����`�@قs�J4���	��RI� �@���b_���^���a�ç&���`L�"\PFK����V�����<'>�@
'��-ӝDwd4I���������As��+�Ut�9���_׭�P(�3p��1�TDܠx���ɖ7��[xr��B�d�6���΄ŭ�p;���>�d��دv/�Ⱥ���\�h��n��`F�}�Z��lǟ���Y#B��dsUD�_�I�Ƥ<��3�l�rU�� �C��4Z#`w�9�V���p��n�
�7_�w����g��S��`�q����潹���B#�uK�ej��ͨ�~�*O�����x�U<�]�U��cC��\{���<��oRn䱪(�5>�ewh(���%� Ԟ�.v���/�=:"��{y��u�8YҔ�Yp������S��O�b�����I7��ա%��#�r�&���#j���PΧ�æ�Z)���BW|�~��Y΄��Vz�/��Vyq.��8"��l�F��1�!�޹�OX��u[��O���`��.��*4R&n�>\(P��+�+*���K-�fPh>���A�_mKSL0�yau�_W����|_e�]��ľ��������-@�-ȩQ�x�R�ԧM�u0Fj�Z�j�}�$�:�.T6�����9����5,`䦲��
�u��� <V��G�0�z��t5E�5���s�� [����u	�I>����r���������-�
_��>]ɁH����^��<�%H��,ʹEY��ak'��;����?!#6��YGS�K�~x��Dӄ��|]h.��Y��_����;�wti�f����~���]"���?��B�/Z�O0�R�vߝņ;n��&W����9���`/�5���?��Kq��=$g�rk4��%���GK�;o��(��qj[/�*����_W��.����H�.ƪJ2��W�uԅ�������$��ڛ?�)��aU����b�O˓~�n�2Iԫ;�⎝8�N@J.-�r��ш��ȝR�9����L	�/��H�n�B1���E�s��#H�(�B?��ҖN�7��k��B۴����~�:���$��3����_���q8�b�7���za�|�Glh�u<k���`�d��y�a#�b�3���3Pp�s�'[Z��$ڬ�-�۶�'�U��2�oiAH��_K��;�e0� �¬��:��s��.��.ϓ;c:�����*0G�
}�q3r�JN������c�y��6'}�C��F�/�YP�dc���'�l[��>��Z5d���
�K(w{��9��eBtu�ϖ?�T+�����Ƨ�ERГ�{����_����Y��l�_�0|T�]��7�fP�C�tg�؎�g��ٹ�)z�
&Ѭ�NҢ�5I|��.��=��Aeq��k�큵<7��W���=XVd��T�����19u$Y@>�H��u����|T7�ù�ݷ{1��Ώ'0�ҳ�EL6At�*ѰC�!d�Е���������y�
�(�lG�{�L���R���,/>���;�ʿvMgW�B�Ǎ)��yIH��y,n�ڛ���b�(r��݀�m�+E7P�m�H�0�M�p�����*ϣ(b�7fE�&dT{i;�<�_��an�d����W*I�D��"w������#�K5����88�N�*#��/z1���&���{��6C��,+�ij0!��R��N*:�5V�i�~���S�&!h�,����4t��ֽ]�!,��z�kdQ��l�Pk�+t��>��R��u����v*h�.����0'C�`?ϰX��2{�T��qIZk;����fعm��է%=�����ZO)�g�$���e+�H�g��3��$��0{&j/܄�,'GdbMx%���0G"�����~�>	��f�]h&�EBV��'�Lv�14����t9��yFlm�L�[�Y�(�A�g9�>8G`7(*upX+�vNZ��ǲ�+����&��"����$�N'�
�Ybg:�}L�e���?e���r0�����D~����F�\;Un�>F�F���6��:������l��{��o�'�,dq�X�Ή"�h�Q�c�=��=��{z�����~���4H�zI��T�*���&Ɖ
}!n+�O��׿܇��t�\8䡁���ַ#��K�2X!6qp�2������;(ZAM�ִ??�Zh밒
f�G���c�`XR�����^��H�+�ݔ=Ca�Dp��~�v�p*ف	�v��.@��O� %C��U���K����n�6�� "���I��[�kMKQh��j|\�����<D�����
b�(�E�}�@�Eǥ�Z�[��|�<��7-�B��!���@ I n[�A�"�>�UN����p&x\����O{�Xr��;�ZJ`�&R�Ϳ6uG3mxj(lڌ( ��|�y����0E&����1���tD�e�!�n]:L�Ѝ��5i����7��T[����?� "�_&M�_b�{��[�j�nT�'�HT���8eC��\�T?��U�oFdj��

�2c��`7w�d��ca˻���Q���3&m��
|��M����	��h�9*	ĥ��2k�,ǻ؞9̒��㭦�AC�����,�׌�WK1V��S��y7u��O�
�%��,=�G�<ՎL϶VWI���ǀBe�ߜ4�-�yHy��Z�(Y|j���ՔfCقȴ�N��|�-Aǳ��Fn(C�-��,�:a4���W� /TE-#��
\}�8�f.�gE��sF�-{��L�+���苈����]��%�RP�,��[���Gz슓��T��'dz����w����y}l�w�Fӎ'�i�{O��qmh�y>�ֵ*�] �*��oŝ��G��d����ƭ�nS�|�Q�zx�?W��zZw�4b����?ؘ�qe�����[��x�7����M�D���Ƽ>n(��} ��鱯7,RUH��H#�)���y��x��~�Ԍx;T���i`�����.�*�3�7��J⼻�� p�	�3�抈1fZ�$�<�M�o���X?��H�Nb��+1�+�J�X���i�|��c�V���,�v4P���T	�A_/J���X����3�/�m��GI�G�Y�����k�k�kC8p�8@h��4��f�MRk^��魀@NH��>h����-�)o^pI4ĸ�um;��������8�
��Z��iq?*��a�L�ts��[ن� <��7-������n��U��U�mTw��� ���N.�j'�%[�����8GNäKh��מh�-���7��n,+֘���2�����拊�l9��8v�dS�/���n4�{��1��ԕ�%��T/I���R��ݺ��>bB n�Y��E����z���y+����6@k�N$���'��>���>1�L��#,s�*Z�|�a-ࡳ�·U���+tM��p����8�L�XOl	%�6�{W��
 ��V?�������N7똣����gJmq#���K!bH�B�k�9B�	9�*;5U\	�w �e
5^X/�T�_�a5�62'xmb第
��������K�Gʣ#"���8a�����l�,��i>�-�lI�y-���N_��w�#�y� �/��W:
����Sُ�k.�>D[g�K�v#������1��'vT�〰<�%��Dі�m�O���&/i.}i��6s�����GP��eL���`;h��(cH�9Ln/ל>�.��F���ɤEȚ�a�"|�KBݷ��+؀Gr-��2B��H:	���v�p��
8�
�[z"`Nt��cN��揆��I��vڗ"�y��<��W�C�1��ⵅ�oIL�$ϡ��y�����'"�j2�՛������<�Mw-�M>��CW: �җ!7�ݥa�9��4��n��n�*oA-BTz&��b𷃷���9O�^���oj/���;0<O�|}���O$��'�o�àj����c�}����w�l�P���M�l�)�B5�w�z@�T�M�u����#D<�t��ޖ�ThʙK���͙�'�F;ҩ�2���R��<Vx,@~���[qϖ:���.q��t*3��,����AǑ5�D�d��}cy�j]~e�h�awl�$!�.�d������u�Ҩ�� �G��P��R,T#� u�Pm����mD0=����q���U��c�D�ۚs