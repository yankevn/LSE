��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+����=n� Lv���:>CQ����̛޺�/�,�]C	�/P7SkT��V���0>�܏�.� Ȩ����O���c���(�����6��ƂY-oUIx}��]d ��� �D��W^�xȚ���Ml�2�*��9�����}�$<�5��)�lY���CHM�O�1:�p��9ld��Lz��-�U� 'x�o���	��,�Q�^y�YB*�Z�1��p���}U�Y�W�8�%���(���tsuD_�SNAe���{S:|�/@e_<3FgL���|���q������f�JuY��"�i�X@]o��O�Ub�6�D�frD@{�|����#���o��g������nl2�e<7�(�L.��KLP�\�_ņ��p��:ǧo�	��'���z���x�T�����)�\�D�6���~��dKUa����]Ry��'�������h����������f�(Lw%��6�� y��C��@m��ni�y�Tm�WLc�#t�����zc��!k�Su�b�x�O�z_z��L({���hi�9�?R���?e��Z�0�w��m&��p������v1;�{|g��e�<\#�Ȏ[-gH��CR	LJ������Y��P���/Q.WR��U�KȾ����y�����P]}CAA��h��CZ矰�]�'fI�~��#e�F��`e�T�Ȏ�P�pG�(y7�KR�Gh��픓��0�e�:Zuި�R����N��[w�S��כR�_��8[���ma=�_��N翜`ѩz�v;��Y�����t���r"Y�oA���ˮ��Z0��^�Զ?���s�kV|*����,��i�f)��I�ΟF�ErlZzYP�-�P4q�Jh�3*NNʩ�`��z� ~e�G�o�j�w����2��B�>Y��A�K8��9hD�磬|'�P/�����`��������}I�������<�R7Rɟ�P��$�v���p��]J[�Y2+����K�_^���������Č9v[>�J��-�� ��S��*�G��^1�l���]��q}�C�؍侫����sZM^jp���؉��L����쀚Q.7(4>?I��w!?[,��:���g�E�QS?:
��� V�QI~�4�tv�NO�5Dx�fQ)��D~�E�F2[��SY�7��Ѕ�Q,��(�Û�N-���L9a;������`.倽�fڳv	޹�Nr3��#�����[�G�Q&�s��{�*d��"3%�G�-I`��/`m���D'7��?Ő;����I�UFOl�jsa~���$��"�բET'�,N uƐ���N~a���8HsK!CVpZ�j!�Š׸�<(S�9>�tFT����z"�܋���$�p��������a.�w�h�~:�r�)�
Ϊ"�s�	2rd��vN�_�/�D��7��^��cӂDY2}������0�u�k��	r�2�n=O%�D�#�K�&��J����u_��1�IG���i_��
S*{~��e��CVLsdT�h޴����-�jl��1���~���ӆ�i�b��;�v(�H�d�(�����4�π�/z�ѯ��|jv^�8D?���3�k��Y���Rн�=fa�0����ҁ��QW�;E�,�x��b4HV-�*5�B�Ŏ��=����g��&}S�.�'ڵ-��5��1���
O�A�
y�#�fo�?��AK�>'���ʀ�4"�&���>���̀s5��G��5��7V͐/M��i�`��}M�a��2//M��]�Y�à����1�]Dc)<u��z�J�r7�UKȮl�� �2ʎR���#�Ȥ%�E��X�Y_���5^1�s�7۔���sn�%Ĥr���1-l����c[K���n0��8�BD�db� �Q�?^�2��1�q/G2kq>�a�x;�)�j�P�vF��a�
�	?�I���l��O�K�,�5�TW��,[���z�Ɂ�Qĥ�h��m	c:2yW��H䁔�$�Z��e�����rz�m���!|fMKʢ�Z|t���\9�� �*��lS�7��h/sU{�Ea�q���q����*�&�{��͠��S��t�]�S�@QX�X������u�Ak��Q���x�i�lw@��/l��)x,�Φ{����++K�/�A�2��l��6-�Z��A��ȉ.�!6Ѷ�Bz���Xùe���
3�,��	�W�1q4�ݙ�����8�P�.a̰�� 6�q�.�i�G,I���I푋D��[�J���S�~�6&%4)�����>�A�ƣ�XGLZ�ۋ�����V�P��JOV"��g�{p�b�lڥbM��nX]���	3�������j��r���_J��9�x뤹cA߲�䑟q��,��͛9ϥ��S���v�D2�J#���,zKa`�(FD^eb��5�/��Z��X��%�x=Zɡdq�[T�ȏ��DgĒ�J?�,�W7��[����+����~v*U�K�$l�˘���, /p}<-��ge�,��&�`��Nݻ������i������bW�ӏ��ވ΃�vqg5r?�A Y�w��AtǊ�o�hDr��M ��������05�&�W��PK�3�)����)�wec���U��d1�����A�!O
��2�횑��ٟGӢ6�Z��VGYx#�mV=.�5���G��\��5�נ7�Q:
��\�J0_d�o]����O�-���)q��L�3�u�Xmt�ͬ�l��jXL4��aF�#�H��t?w�R7