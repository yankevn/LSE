��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�\|�m�2X�q�gV�^)U|e~�)6 ���zX�G���T����%��/2v�
v=A7��������ba����y�k��SL����d$WҾ��ԡ�(��D%�k�Aq�����Q>�^5'����.�G����5B�L��p�`�SΈdZ�Ӭ�90cI�d�5<��=_T����e��������iΰuRg��D}��]E�γ���P�n�LV��j�XE�hFGzljI���<A�`P�{v \�sX�m�y�7�c�t����/�~�-C(j�PR��mm++�(�S����(LNd�� �ܶ��"�!�c��F�ֹ�r]{���@�4���y���a�ˮ�v�:Q4�{�˲Y���k���S�;���P��|lm�&h�I��0w��0\�<H��|�3W=�n�,��+y����W�;���tۤKI��U�{]l�O�/&o陿�Cv?=�5��`�R�W�s����"P6��c��7��� 整2�j漢�_��b�W��%4��I�]�t���uV6�y��	���s���#�ܹ0�śP�7�9�']A�ܜNi��r���F�MQ���:F����n|Z�5�nJ�$S��y!�}�7�O��Z
z��Lw�#��T��4 >��f܋��u��ŜD��3��;�:��w�tw��C���}�B5�Z�?��-�#Ja8�^�82J!��t��}����9�']���(�wH��ZM����-�ÖG� f�*i�Kύ�>���T��=tt���>��jVnu��wl�\E�ah!����� z�VQ�όc����@	�J�7�T��Ǥ�=e�NH��a��Z����?b�h��Z�_��Y°o��" �r�f�*7n�.	����(����T�,���C�KA�M߿ ,��?�%&�ar�`����}E�C8Q�⢑�K�����]�:�5��p8�`�C�ܙY�;F�q��G��2�����'A���?��&b��MX��bv�
��i�8�gD//S[��<����
#����bjQmn���N���y@���]�`{�@�B� �YjA��
�Q��_������3s��KiA�����(l^L/�ZV�|Vg��A�4g�KD�4��@�Rm�'��6�U���a�}�UG����&<�a��yT"�XX�%^u�'�W&� �c͟�aÅF����|�4����$y�L1}u��E[>��{�#��'9n�@��D��X�k�H���Ҿ�I�t!G�k��c1�zx#�!�{�$h�qP[q@���$�g[�T�Ws�*�I�\�|Nϐ�X�΅u�t�M��`S�TO	�����z�P��3-GI%�mzC9���O�r^���T��;+��𞑸)j[�U����Tu����L��K'rFʏ�`)��b"�m�:���;s#xj�K�"����Zp⑰�{T�SF��z�N���.��f9`�C񁣉�eB@X��l��(��6�&y�����>O�V����\�+�"X��G3}y�6�|POh������F%@�j
�4�TĘ}�@��#����+�G�}��V��-�r8Y�Ҝ��L��(�ط!��'�Ryv}���57-_��d�[q���e�3=��[`�ҹA]�'Յ0-�.�\�+�-{�;7��K��tSW��ܣJ�9���l_�k�������Qٔ�I��?Z$��|�E�X��)s���A*.A���y�+��,��`�Y��q�~r�(���&G�m
�1s��2�p&ͥj�M�kӂ�� �<��xQ3���*�7�rk�X�a1�#����^q�-.28<�p�Eh���}��A���7Њ)�dZ�{%�5��M�b`||�F�2ksS���J���Р�'MǺ�\lv}�PQ��$�J�60B����~�>�<8�v4ӳ4�ʌ��U|�bчcl��Ύ�!~3��)�W�`�M��HZ���q-����B,�Z�k�c,�����.ɾ�޸b�$yk�b�:x�3пZ��cj�f���3�62��,O�>D�@��;�H�wt��{���hu�X����ST�������0b[ư5K��5Ɠ���'�uc�M3f/�U���Y�p���
���I)|Ɠnr޶��Ɯ��k�em(3��z��t�.��N�i�twLZ�������Yi\7]!�_
�[�w�b�c4�a 6D�[�B��xA9�,iW���4ev�����R��@�t�ŧ����MǲT|	�A�&�}q� Y�ˊ .ؑ�!��/���z����S��r?����Z7{�נ�2��j@�賅��YIV>���z�}��#�<��ZCV�B�f���Ŝ]��Q8�)���S^eGU���:lX�b�8P��v~�b��/%�u�{�z�&�W@�:E_g�xp�E�x�;�&�U>�lƢ�h�d,5�*�U)^u�.�P�lw��x�x�h�0��u;UVԗ��==�򍥼[��{iw���Q�Ճb{1�טf�W$�����!�v�Ng���H1�K��8�{"8��e��p�8��[M��u��/�n�����b��8+ ��w��:�w�0Y�V����������AĹ5h��	�	��WH�XP��
�}~`>s�}?[[�s)�#`BiQm]�eHJ�v��02@`g�f�m�座ǀ�%:���F��.K7���+>e�ڡ�� ��2Q��@��vp�>T��M��D�pS����ڜcª	���>k0��(��2�������*��AM��ɣC�1�bI�^�䔚�0^�BkL�V��m���f�:*�XV�FS�{�-�o>ntĻ�ƚb�7\}O�����
��r���|���+��1\��Q)>��M��n��/m.ф��ȑ@[�����־����=�ۈKݞ�YL����j�o:M�Zmuk�3 ��R� �G4�+@�\Q�E���!�,�s�3��ߗf���_d7�4[r�������*�I�y���[G�{�t�`_�����1١��6&�oqd���B���D�{�wi���J���/�����d����$�x�a��r�4	z��������/2'����Ǡ`V�-G\'����;��T��sE�<���U�!	�c��0-�n�큚���`yY��bϻD�1,0�o�B��*|"{�r�R� D�ۍ�'��X6�+w['z�8l6z���G���E?���p�/�>��ϐ#dM����&��j�&ǋ�~n�#m%x�D
Q�9(�i�����L(K1$2�� �'�!����
��g�C�%#��c:��z�������j�'�H~h me��6���J��N�:B���u#8��M�@()@�d֜�Is4b�#ō<����g�A̔Ǽ�s�X�i�|�7VW(���
�l�M�(��R��Xy�l�`4���%�f�w4�X 9 v��M6�\,�2T`�%��Kh��ۉ����N�����{p�RzŎF��XMɤZZ�k����)���*�q�����Y�7�>~��"3�i�;@�u��lO�]����W�ܐ�����X<L��8���LI+���Y��Z	��P�/���[D�Oyz��*̱*�b�:?�0�k�/��A�ɣ���G^L�?�@e���Ak>�x�h2��%�8?��V�|�vL��f�q�F�7�u�цp�?�!���bVR��d�ni�4������G�Y����-�Q��z8\��Gt�z�9���Y ō��w|?��|��t�JD���ǭ_U�v�]#i�޷��(�6������i��r΁1�7K��+��[ߪDf���
��ʵ��!�1!d9�,�!�����r�[������>T8a�9�����@�]E�_�i:�V�-`w~Q+�#vfU�/.���X���LuB�w��H�V�KZ+�0�

�n����H�Ƌ~32������Hֶ���dC51�<��Qi�=��'��H[b�I�8��aE���P�-���`/�
����=��̤8���.s^��܆I��T��Ƹh7��$�v��� ���&��ɫBY;�$�y	/�ˠ��2\�P���J/����(y���R����<���Ո����cy�+�C%��M��nJ�V�/�i�X�Ut��;��A�~b�@����z���
��c�7�F�p���B�7�U�aͳ^G!�l��M?���g�OJ�"E���=ISz�;��n�dXz���D�L����Ѣ NA]���Y�x����^oU�V��[|GG����8#Zc�B�J0���k� rec
RDJvI��Q�$r]��;dν�C�s�����������][U�Z��d��]-���)��yG�O"Kg�7�^<K�A	뇹'�T5
�n�/�w�
ʳ�>9����$����3��O�9�k�rҠD��c����i�e��5)$��sި�x��n4 J��i�Sff���w�b����v����J�ߌ\�W����/!�T������l)��U��P
�6����q�ʃ�}A	�1����M쳐���f�ź�ֱ4���6�H�5����"�@\��ύ�_�U.\<-:d@I&Ր�7��>�8 ��%!2�"��@y&_�0$��Ŷ>[�����<�������v�ʾo�;�U�(�DȽ����k~�:<[�t3l�`�K�թ<�Gk��ߟ~�A.�������XI��9�;Љ+���t�
ڔ�����K�����NB��[�s�#z���i�;�A YgY&��l;0��%��F�!�m���B��M	�tٖ·�9��q��K����@�$o���B����4��>�ך��ԭe"�\�l��ׄ�s^_.��E}���{��-���Gf_��\�:���?��Ed����mR8��$T8j=���K5�UbN���f5Ks��}��>�/P��
ׯ��KA�}t_`5�Jp� bk���h�!3�轇k5@K�^3P�$��.��N݅�%pƶ�,�w�.�������7�ԏ/��M�[+�����5J���G�(�e������Q��.�ª��{��~k^u)�	6
���"v�?��Ly���L5nr�K꿸RHI#��U^�vk���v}�đM�Ty�pX��\8����+�����kɕg�!�2�����KsH�3�����|ѕF�{c�)�����8
�����Mf�5Ɖ�cht�Ӧ2�b-S%+=�/��Mk�TF���+��4���2�H�w���zE����}f�T�澮Z+�%R�
�.�W?iF��,������iV��t�g�p�ڮ�I�[J�0G��M��+�#0����%������]���0��՟Ϛ2�y�nf�·�z�|g�/����;G��}��-Xs�y�� ��\o�v������mb��V����T!vՊD1����a9Z�f+"ϻ`r�6y�-�����p�{s*C��e���ZT'<]���|ng��7@��w�5��<'�Y� `�'K�Z%�g�v��6���~U�
% �K�|��Ǣׯ]X�3���`��м������x���r���7JH_�&���'�+O�;�I���)I.��ٛ���^P$���#r���)��	� �Q""[����ό�`�T7Z��q�V��Аn�>%w=����o�z�%��;N�+��Q��QJ��}2;��>�����L�C���/.N6�`��lx�Pmw�m���x���Y13�0|�e��Nh�?�����z����vвÖ�x����|��!l�^�jʏN���ڻcj��A�}nn5t��p)`3�,��2�&.�m�k� �q�eߎϩ�,[&#���!z�eM�[ !;��Y=u�8`�/�FŢ��Z&(�6l2�RV{�܄�>%)sfۉ�j3xP��D@Z ���̥:�v[��'��]e��V�1ߪ1�C�� �c�P"��Z�@�D$��S#�������j�?���Qޜ� �aTX<��	ǴJ�FyP-O) �K�G��|Y+�6K53���-�Ә�ܛ)HT[g���K�~��"i��D���ͥ�1<Nb�E{�VNλ���(]�k/�8GZ��JA����b����=�
�κ�H�`(9����Hbf�\�p��ej/ͧ+�([�e��w|
.��ܵ�ӷ�-��b�5�z*�Q��"K�p�L���;`�c�@���U��fI�>EO�C�9�xrC�~wSs�qR�����s����&��Hy�J�ο���
ڜ1�~�~+�c$o���7��恾�����2vlK�	";b��J�ʲ�v����c�_g������Շ&�_�J!��ր. oS~���I�a���>J�(�/*�
�>R�����x �}kė-�ڟ:e2�v(.����1�
Z�$:L0���¨/�| ��y�_��?�n��E�(�PU���y�1��T�_)9�k�pz���m�I\�}4#\�d`xB���|LyjL�0Rm\�+H[P<��3]뺂�P���/lX��!��cA"�9�s�m�.v���J#�X��J��z������^�p�\�Jd��_:>l����1��z�7���N����}��_��~��},tk���m*�p��)<:���;�JQl�g�>��?[����R�"#l�Ũ6x�֒��^�~�'�u-W�8����&5&�Fdđ2g���
�a��/|��4���bYh�(��o�G�� �QP��[A?��Cb����9�|;)�q$!�ç�����ǁH����S�(~�D����r�xnIm��u�R
É����"f��֌�'�7HA�.&��#[��n���a��")2Z�m5sŅ7�Ge5������b�����݊�`���UB��k��w)�_M#;��:�-�n�)�n=F{���"!��M0
NV���
Ѣ�T�(���}�9sm�
SF����g�l��$��r#�uq��!AB��=�O�_��@[����uT�v����:�����#��G��#z���,�ؚt��f=�ucQ
o����ˇ5�2�@�)��r�2�B�r�S�<���wu\'Ku����ϟ��*�V`:O���d^�H��)���@f� ��7T��:�ux�%�&�rvGɎ�F������jMh�3Ea\����nIgT�O�]RA����;5�.��).</U��꽫^+B��.VTؽiA e��L��'_6g�BB!��}�F�S��F̥cX��Ox������ʇ`����=�ˆ��w#���V��9j���|+�t�Q
�a�S��oq}��SiRIBJN0b!�/�MGՎg�vH�Z6�Q��3�w��;b�x��:�+>�*p�-�������61�F��$ύ['�ޜ<�6��	02��T6�VI��G�����evmZ��̮hϲ����<	
���L�*HBZ�x�.�q~m�O����WC���7���z�1Fy;[��1��e7x�������nH��"E:'�7�,h 9Ҏ�J#�?�PӅ9}fU`�Re6L��~.h���d�tn:�")�2�آ@�����1Ⱦ���	s_R&nc(t�1hIE1�2�F�@��C��E8���p�Ҧ.���h�Քq3�_��ՙ��+i`�ٟr+��K$��p�S����X努��6�9��R#}�Bl�Ӻ��\'����-�S���d��g�.�u�}�D�J��$_(��Xe ����y��+x,���P���IMf��d�8��Y�_�i�s5�w�I7+��Ζ�N�4^�l�*�����D��'C����@�sd�m0Q��$/(��e�Z�E�y-B���%�JDS������o���_��i��p��O��m�ФâbrN�`���NnN�S�R.�N�s���� �*��sުԩ>�@B �!K�~��Mzi6S�)-U�@��ٗ�VY!���n��1�s�n5�7`D�cϲhB�?��<��[�![&�X���fkZ�k�kfe���mm3��9�dQD��#���M�E#�]�z�W*�����o��AX��Gv�#�r�e���Y�=[Q�Kxu"#�7i���e��7L�O�` ��;�b	����
���ƛ�X����À��P��2���Z��o��F�T��@d"����C
䍼5�̜}�}�Py�$ }A ZL��t�д��=���Tm3Ɨ�Fs�Ƒs�z�I���P�)�ŋ���	O�:��!i�q�
�G�#�B��^{j�&��
C�L%=T0d3<Ø���CD�au�ֵ:�u�+CDL4qI�v5�Km�t�2��G���v&йj��lK�`C�W޶���{�(�Xk����wCt8+��ܻ�%���s��|So~C0~g2XѤ&uqI���&&dO�����[��]��zk�D>��J��ٌ�#bW6I�$q�<aN��4��d���� 'z��+r�3|����9��'bA�[��D�1Iq-�Cu-�����ڛmky�?꽇�E>�M
@���������ͩ���:���+Ȩ�e<A�wޢ�?Gz%��WG=��1Db;cal��R�U�ø6��$�����9��_F#�޿���A��9�!���9�֣+�,�%��>;�@�;���@�6U�D9.X�ׂս��U�ƪ�#�9��U������6��Q�Yd�-"\V������☩���$_���V����Fb���<��T0)�ܒ1��^�YۼԨ�-n2���uSk�j�h���b� u���c�����7&����W'���ٜ`��l�7Ҧ��6�
]���c���k��tSe���-I�	�R{��M#�cFk|�B���W?�0\&6I5������L�S�׊�Rv��VZ���٤O�+�߸[Zy)(`�/���b�A�,��Z��/Z��T�Â�X��?�y��׹,���?�����L
V��zgضi|�$�u^Y�䰊Dr�����$|{�uX�n�L��	h'H��!��8���?���Z�>w�[?�Z6�^T7���E>�'��|Ab,��,��^)�Z-9�����E��~5Z��J���ч�?�K��_.���t�>��i���������"S��7��5���v���"��ꂰٻ*���AC���r��c �X�x��]w���g^zL]3-�?�;2Oe�Z�=��%�=��='��(��1���}�)��~-VX����̛�1Ϩ��6ei1�׺���A�&z�,�L�a4ۊ��^�w�����h�JB	6��K}�f[����)�N	4�{�����ZG��䈋o��/���E���k�p>΄����䈟�ɰ�w��s݆%��4=�*3/=�b'FT�Z0AtM��!�Ċ׭]��7��k9C�Ƥ�W:���6��V����_���ﵴ�\6髥n����r_ ��	�t5��ٹ�� ����ߥ��Xk4sF�gم���b�"�ۥ�L�b�e��%GmwHҫխ=Ο��(�Z�RU�c��8�#1"�i��_o`x�qĒrN^�g`4)��HinC�����7*v��[��is�a,ѳ.�����j���O���b�\�k����g�[1�w>����8��!�{�<��W�>�Q���	����]P��ob��k����v?9����^��ٝ��.3��崔�M2h$�-�͍��rJ����0h_�Əe�s\mI��)������7�l�1�E���Gt��`�2ޖ��JE �Ŷ��zJG���|�U����Rt d`��2o�� 	ʑU����]ەǓ�.����,�<([��|ɻ�<�������A̵�c��t�W�>���j��������Ċ��+���	�����I~�� �1N��[��0M4�M{�b���(G��?��1⥶np5P�Z�6�N��={p���H߷���-�΁$�+�v��b��DE��	a(_�ŚO�L�,-{)���S��y�$O����L�#���vSF"�Hfõ�}!fZ���~7�1�f�m&��E�|c%����O�M_�7��	�:ax-3���@'O�fFG�
F�W4��ޓ߂�-�8ѫE�#�?.iQ>1�$;�������.�:�������,b���҉uerS*k?^�X�Xt��2��~os�� ��b�w�� 7��� �!���&߼dﮂJ_�M�x!n�{6�\Es��o����j ���������}��x$�~����ԏxk�Zf�#4*c��̳�����u�?�o9k}�=,X���΅��[+`8 1���qQ��ʹ�2|GG5�BE)�Xg}n5�~��Qk5,3>�*6��^�J.L���y�$Fؖ��M7ƅ�I��ߪ<.�x?�g��v�5��G��C� �yXj�\��u��.�ԏܿ;v\�^�ұV��4��hd�o�\�3 �4W�Ӕo"�4���ω��.�k�wh�\"��b6��Zfr�D��g�ɼ�·����+.�N��i� �&Z��M��BI���;L��oy[v�#Y���=7O5��O�l�i���"��Ct*�,K�p�6[��qs��%���b!4��7�H�s�g[�� ��+�p#��n]���y�^1�Ŋ/��8� %P���\��γy�B��������62Zu����T��"���b��:N�b����l�5�)�w��[`Y�����[��*Ft/҅/$�a ]�/�N��|�%㠡-��3�p^l�߼�S��#�'�
"���mW�p.�+�l�Q�O4<h���:=nn��;�_נG˫����E_�|�1�X;&o�bi�N�G�d>�������Vã�@���}g�]*���;�����K��k<"�nb�y�w{���e����ݮ��O�{�h��^yY�B����Ѕ�`� ��8e���j8�R�V �TF�ڿ��oY�&[���_�A�P�ڡYe�N�D'����w���զS<I�Ȥ��rzZ�O�]��l��u���^���d,~����xF!!�@���~g���g9�w h�B{�Hr�w[��\7�G H�nrk�M-��%��ǘ�+Vf�GQ�(�W0��p ���{�h�@��E�@�ý���