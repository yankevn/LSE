��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��?�I�J���6�oe�"�<��dZ�d2��
���!�b��s�~#��-�- ��S�K�S?
���2�T �.�X*Q8��=kH�cl��f���h������$��pl�u��mW��Y���1!��d�>��X<�ݱ(�z��R�M�@ڃ)Y�Jg�p���Y�/7��ΛZC�oX�`h6���	�h<S���2~�{su;"-zb璌Q-MT�${�J_	������u��ׅ?}&�,��(B��� ��-�TiAӎ�?ָ�Z�I���LN��'r�c���X��u�G%eWPьrG��B��5�t*�T�5�Jh����T�b`_��x�:ǃ�g�as��CY������#�BF�5)�2,Y���(�z����=L��%M�jYWa�"M����|H=���Y=��A�dK����p���h/���I��AY�i9%�;FX)2�z�M��{!�ь���<�;���p�,�)�f�C��t'i��.��X�Iq�o��?�:�ya�m�.�0�����[k�j_(`�PaU�jˡ�e)18����(=��,3��щ(]۹��s�=���n/k������+_{��?gV-;b�,�[l~�>��~'�;^.s��>��qJR�ĝ��P�>4x��gm�ϋ8�}kt��S�;�%�d_�#�j�V����v��;X���_�-*?8��z���>ђfe'D
Px��٬pm�q���~�(�L����X��v����'>���,�0>M��p��Z�M�F���;M���E"�� ��Ea���#�)e����l0���V"{�]v{�Ź���	fJ��k�[$�74���Y�a�E����L�m���9bŀ�����J��&������e<�$(5��7{܂6ؓ��XT'�_��k��9Z��;��4��
.J]:��'��P��:?E��#F�[�D9�U�A�T�AI�lI�_2��[l�!j��r�2߹(Ĩ�]����0�T�ȥ� ���s��t�k_�r<����0tMx�V
!���
iD�#,�J�U����l����L�g�V��jk���\��g9,h������OA<i%ꩱ�߉���IM�>��W<�u�-z1�K������Ng8����g��?�P��eF<�wJ��A��AVδ��L�ӻ9\������UdL���>$�1�Z�ךd�z׹j+ɯh��,W���*:/��"�|��V/e�=VO�����e��O���͉⮸��K��0C�K��L۽�3���	����(DV3��i���//���e��{~f$c�8��e]��T�����<G�D�-T#�&�f0�ټ~C0"�!�PSD	���JR|���@BY�l�]���*D�4�d�;�
P�2�2y��@J�kq̺|f���[}�ɵ��<���Fm2�j���DG/��O���7��'�5e �r�CP�n���,�nף��7�dT���;���vAb�������ȋ��Y��M�at/: 0��X��y�d�R��=l������E�J�e��x����֏�Mlƻ|[4fMJcdqB.}o�]�n6ә ��K�h~��S���p2�����:�vj�&�S+��I���=n�f-2���P��a�Y�'�SIc���ш��x(<���2>�;?R1;[�ԛb��Lrw���iO�5Ȍ#����|Kq�C���rj�x��s�Yb!��jQW1�����o�s�-�����]U{�o�یO|�$���<n�h��2D���~�K+�Y�i�Xz~h���36} ���� �ۂ�r,QUأ�(�����Ѥۺ<w����5
c�A)3a�D�}�F¶�
��$Z�`QEV�Қ]���;��}ܦ���K0��3Q4˯,f�F��rLK�w֦h*<�.�(EKř/��M�`F��������5O�6n�,av�x��L$��
.�QLv�G�0_܆W�?*9WN���ѝ���ăe�p�H���{�;t�D��(�ɟc�o�N��(Ps{+p� ]ǊP��?Y�i!{8�)}#���� !�
;�+ϐ�Ԅ�0��mFdd��5f���x���m�e̷��İ6u��$u�R��`�W�λ���h��x��}?<n6�S���R�����⁧�̋����A����7�鎽�Y���/>�=<�[���y3<���(j~����ɖ���6�����з�ǟ��]�P�9��*�k��Uc���!d-	2����c<Z�ANqvjy���S쎋��_�(t��o\��`Kj�;7��pn�;�#�F��?_�-�.g����0�u�+1c������[�[�K�<�+*T�e7��@b�>�vNMsh�KR���IG[
�{���#��a�9��D)%���G����/ȂP�$�(��wy�3U���{�A�<qk���e��@���m�K, b���9���-�m�8��E�ߢ,>���m����Ƹ2��JI��[�=)�4��c&�
ry3��DV.Km��LS��ʨ�7�N�A&=�T�񥐦_�w]�� ��T���h@����:i�Ë�`*&��'KͲ	�]!�d�.Ҕ�2҆O9�j~��o§�M'���/��# �X2�*�#a\�Y����za�T��8Ї?�,�F�po�f�#��1�\r��|�QQ���x�dXS�� s��	���^�q�CG	�)�߾����D� �qBmD+�ɟAw�H*��@
C�=���<[bt��E�k���R;�k�#�<C�(��1X�h���-�y޶�tA>�â��6z��������5:U#���Z�w��<�l�n.�}xor���V�ZaOKV�_1�/ɱ�z7��_4��hr'��A[��qT���B�l#{cɪ��XZŽϺs��*]�E�^[���G_딿���v��.��|J�w.�Q՘�����Q?W5����@F�"SV���u�v��TyŚ$�&�2<"�����q��tW���^����e��JA��+R*�ŀӴOH�����R��H�2ܡF���%�M��Bv��#o���s��s�r�So��D����K�d�6�#0E{t� 0J��s�Ej(�N?V=�m��T��]EМ5�B�߱wK)�~��5��ț��:��F�sA%����(�	.$�����=4LMW������ȍ���i;�%����E�FBjs��u���y?ʅ��"�K�l�	aE)�i}�V��ݖLt)Y3�zi1	O�v�(Y��9�O���٧u���^	o�Z����J@Nd�KWb�� ח�^�[��kB��|<��lF��/~1��$ԫ�ڻ?�^�?�~�	��W�l�;/�2Eg3�rr={�TaV���������,E�����:!�<8f��"{0c��61�Y���SS�gB�i��������ޮ]�]3���=�o�z����W�U7��m���L~�  Gp�k�� :#F5}~��8� �g����N!Ú�_y�V���X��3v����}�E<�*A�>'��9�5{��G���Z�L眻!J��z0(<�A�Ř�d���Q~ɱ��%��j�A�v�c�0��8t���ëTeS���3X�9��̴,���[0>is�)dn2��	�}�(����dƁ8�ki2g����O֔�8S����v�R�+�
�Z�ﵯ�pNdj�(�Sge��|�Ҍ�qHʀP��46����M3T��≬@]�&N�9�ͻm׆�H(�\��Dr�d�O�vП���*���)U-��@��LY�m��G�����zQ��zcI�-xh���g�	ǝ��*a.o�xu=�wO�cjA*lk���E�C��Ri�$X�#�>��P�:붏�$$�vжI� �a�	Z~�����><*��)mV1�\�*�:m�Zu���%d't����4�e�[H�&�c�Uڽf�����j"<�F����"7�]̷rn�7���D�ھ��O�F	UYf����OC����r���KK$/���gh�~��\�&�c�_-��n��L�
��^t
�#���^i�^y�е�N�$3O��R���+��XFG?X�o&�t�}���� p*�@�	��ESU�����~oZ��|��A`z�ǰV�z���g��I3���0������N����I�igR�wQ��r����&�ap������a5�Fh�+L'mh��r�B�\�D�8<��Y\���a�u����a��'�����	L�b���2`����oJT��1�Ӆd����t���$�G���{E����'A��7@�X�b�eJ ��������-}!�E#R��ůp�a ˤ"�N���zu1vT� ����=&wȈ����.��Df�����$���hpډK�ﵥ���0r��ذ=�d���<���B�c�\!ݐ��>�L�IDkr� E�7gH!���e�&�1�����.G������)����ȡ�����)���K2�*��ס��>�E$_Įu��҈Y`�W0���jR�r#-H�7˂�$��{U^G�1v�_F��tg�v�Ҹ�C*��!oޕ��Ǡͦ��9�+j��N'�Ma�J�dK����\; �����*�f��$Կ����Q݇ڽ��/�=��>��#t`s��*����� ���+��ʺ�t4�J�5mzy1�D=S��2�*��LFn��_� ��4��[��G�N�] �M����>�� �p�t*�<WX��x@�����>�nP� �<˿�_�1�8L���%���LuQR&��V8�Za<�d2�OS����hw���C�������'_.�uS���<y[G->*� jZ9V�K͢Am�y9��#?��3�j�#�9���z�!����5��Cv���1�m�$2]2K=� .�����d~Ao�ps��+�vy��*N.�y�<�O����:&�( `o�2�q�1��O%T��|A�s�!LV�Q1� dp0���Z�z� �Q��%���%���@S�@ICjV-O�=���ph���� 4��Q*�Ď����	^�B�NE�?Y����K��b�>��/N���BO���I���ϗal�W��9@�k��!8<�Q����,��Yl�fZ̃d����' h��j�țXTM
��Fg����.������3V2l�<¯���/�$<M�UM�)�]�B�uRX�b����i��&���Hb�� A>�]�A}���_�m���1F�6 �<���0�#W�;@wP��>
�q���5��Ml!��������g�D[z�e�N�$ ����Iw��AA4�SlURm��n�e�L��[6�m����]��:�^����p`(���O��ۏ��ƿK����9��f}DA�,ʂ�C�T�X��N+�^0��f W���'"o��8�:�[�Nd*���>+�!5�r������ϕ��q���(#�[A���A<�1቙�쩘��!��d ��r&�֛��\�AkZq�rȏJѺ4�"���Zlv?)CP����j�C�M_F�˞9liIR��翾	@�6b�Vw0�d�&�͚;)�KÜ��U��_ԏ2��#��ҭP?�ܡ�!���ɋFk}�y.��z����;�B72�ݘ#AŴ ?�Ӭs�:ѽf�s\h�e#���G�!��1l�m���!���{%��+�W�.�k�4�nvl���p=���,�Ȭ(X��cb�	�B䞃�v���;Ќ*j #�W__��:T����Y!Q�3�l�hpW��w�51��%���3�}�ߑ�����&
�k]�)��#��>>3n��n�[��s�Uo״��v��Ȧ�ǺE��a|]Ȧ�e
a�k«̭���;�����{�����du9k9���VU�2}�+ͅ|�/�d^��sb?����v���ʁ]���8���ґX"��B�mXV�a[���8?3���L�e����2�`y8���{I���	]�Şb�[����H�{�)a�.f
	�H��{�̽ C��]�s�(s�"��S�u��+��/������U�N�@��?�y 5;PG��f3H�lP���ǀ����.V���v�r�\=��y4�(�,8�<r?�kj�j��й{��b/�V��u�t�Fi���u}.����UXT�6�X.��':Q���J;n7�~��&~���ma	����2�N�`��н�{^p?�������c�2���G����6�IZ]k�/|H��H�p��|;	��3�>���h]:.���K��o57�H��m,mP4Ibʁ*�E�X7��S�H�5��4���}��
�Or ���q�N%�a�����ux�p=�f���	�>�{�Y��]�&��j�<�K���_��	�4LA��t��Ir����sX�M�il��'�	-u�ao+;����]/~A$��&"�/�K�_�v(7Y9��<�����s��^h����H�����l�������G���n�[zwi���Oe��e�-[죿"cat���2r�7Y�����[�<����Le��oy�" �]vxrX��#
O�|���h�r��_$Y9i~F<��4�[FQ���
��sg�FS�8;��!ء�T��*�/��})�ʶ�qf�&q�HH�DI �;�?��59�?}k�݇����ﴱ�1T��@XQ�/�r���9J=�����~6;
Z9l8E���^�:�B9�*�T^'�n�w��L�A����I��x�#�
�!>��=mԮ��.@p"�u��^�z���]t����^�W�2�BC��zoڑ���rh�7L:�B^�Rk����dOJ8��%H�S��G]�����n��]��5_X�Ķ;�ܯ`4?n�}\��_��pL��O�U��P������v.��7��f
���j�c���x���L��%�P�L��W�=�~���IlbZ1N�Q�襒j_�9�\�Ƌ�%#�P����~j��H޷]���V����A��>�6�=W����6�B��_�&M�i :["�[�"Z`��q+��%2��J�|����=2عUlK�[���o�*�Z���}�ǦP�'�#��X��m���6	�S����;�;��y�9�@��Q2"6 �ݖ�~����X�;A�6���Zw�WB�;䅟�R�h#�dB�}#:9Z-ߏ�,�r����M�!=�IO�L�8U
��\�u�K�ؼ�s�soa�8N��b�H�w��3���T�ն��������;��q�a���M?�:;�D�o�a��z����gg.:uQ�m�P$ͫ��"�TJ�0���c���l��0�W�7W���}�q"hw�u�]7J�둝`@����`j�@>���.��63�.�!��Ŏy��UOw�FJ�$�#P���\v�EEa'��`��C�S��N;*�1E�)A�c��o�y���E�v�����f֪����~�d�m�" �a p�6$�Y o���n{p�1~���N1��@��Z�B���RPL������Iw�>P�������ߠ�_Z�s�w�\Wb�k�؃�-X�!d��P��8w�Ŀ�O} U���3�]��y��"k͏hil��+<�+����Gq�����wh8����A�#��|���&3���lqȔ��L�U@: -��=��ߴt\�$I�и�,Ic�����4��UzFG¿��I���#D��&����O=�6�feٞ�\>���r��T�D�K!	w�H����F�1Ђ��F�\�!t4�󵲼W�خ~(��#Znx����͹R��x�����(J# Ev��ʍ�l�R�`�P�����4[���;)t{�D�<D;GdI�2��q�p�,ۇ]�,�`0�؏�%�,�4kǪ�}5��סg�W輪��7��C6\�?�_�<X9��@��yN1.$�N
�b3��>�B,�P�tJ��!�{+��:�B�H� ��1	��ǻ�`*2G�3�:����XX`Ȕ������q�{ZST3|P��q��2�ߌwUu��WM���סpL|c�.aG9���y���&cs�Wj.s"�{pŔ�|����C)i.d5�������.���D�γn�3�MMA�H@Y.���Q�����t�'_Re֏R�Ш�"0�XF?(^niO1_2q�X�3%��Ǝd�?�LĴd8��}r���A�0\�E�Z���a�A)��b�j�%�bm�c��N�׊�]Xi�dՖ.����^�@�܋	��z[����U]����Q�v�7z���[���F+�fR��g�G��^�Z{/�Bֻ2�����6 q6���L��#�ݫ�5
 �wk��	rK�~�g��������@fO~�j|�b�>�t&����P�z�,)5�0KY��'��>���%��=���>��?q�&8��@�͹���	��T��?ؕ3,F��F�Qv��������q�6��7tS���� �!7�9<�5$�m���B6�U�o�5�?�L�y�v��I�j��J�niho`|b�Ft�ʉZ�0c���ԛm��҈	�T�a�mxvj;H7{�q��I���u�Cq�X?;��6��?g}�K��!��O-h����J���ae�F����^"Z���R��ZB'f�&�Yt xf�}#�i�7�%!G^P�m"9��pb�0/�4��p?>1O��&ZvY��&3��f���a��b��hk"�)�j|Ӷ˥�C�(#� �!x��1<د�&ܢ )�R���tyad�8k��t-�~\{f��?�v�Z�Tq���t~�@��	��ǋ��(�a����u!ң.�'�6'�E� ����N؝���^�����$�W7%���|7.��En���&em�W�/kZ�����Md,u��1Ҷ�,�H��2�������i�h��6�P�t�䳲�:�ٸ�_��>,x�Z@��;�3~iȐ��:�����*p-�j�T:@ng��PP�8�ς�=Q|4�X���{��.4�Jf@G�e�k}wS��!����J��5b��Ī�#m��͹!V$���2�0��Z��Of�%~-�p�h�1�m��la�<M =b�\�Գ��o�������8��S|���_���s�9��1�7m�WޮW���5v���_�.�����y�L���i[
S��D��"���fa�ޥf��$�E�H@�2)� �9�
�%��{/�ͅG��K*]4d�<���M���,l綏��:�$q6䠣kU��'t٦�ʩ���A���\޾�<�O-����TbJI�+�(�i[�K�Ayn�X�����1�'��rh�ǘ�����A�Q9H�/��\9׊�q
[�Ó��{gk�,r��g�*x����R�N=���Q���]�����y�'i��o�EF���^c�t;�u�	�.� i7[ֶ_1�дP�s̞+�@�M��;�fz���f!f����I��u��ۜ�5-��e��6��,w�h����� ��Ҧ������ʎ I����+�,�_�zS�i+��T�F�- �<�u����N���ﻗx��tk+�1�u��3X�]�����Ɉc�K\�I5V\�Ԗ�=ՠ��A�ҢC��In���t`Ƶ�xG(���њ.lݒ�Ҕ�zA�K��+���t�A�����y�:t�4�c�#�����F=�A�G�E:�V���^�.Op�+(d�(ʪ�,?�Ji�|�z��廱�mZN����s�2jfe�ל��ɩ%�ޟ��H\�Lo܎/���&p����1EuD��2Ϩ��#�A�Ї7�5���1D�L��z<���Kc��j��� �u�g�������/A*�v|'�(�m�O���6#�t�Nϐx��U��;<���`�H�Jy�Pj0n��Ԇ'��D�Tr��c)	��횙Ν�~*��Ք�>�?�W��b����n��<kFZ�鍟�|����d����_�������E�VHAm���/ShBy~rوy�$d��z�>���$sK]��W��h���kG�5 �i�Jsr���؁A��,��G�(� ��[��u򂨍ȇbg���0�4�)������ɽ#����P��L�TG����^nep��9R�:��Y��:Z]�[uj�}��HJ 򦯘ͤe8�'J�9C�<�H�Τ�u�#џ�2�)�:(�crS�P��NMDI��(T�������2h9�@��t�Ni�x|Z��D�L���DY3 �_��:%>Ռ�?
�ܖi�V݇l����,�������ʡ!̝H?Β�1Y����nsG��Ȍc���u%��9�B:�J��Fs,�
�Щ!kW�)�BX�yg�b�Q�99vZp
��<�:&�+Sj)�녭H���&�d��z��A+�T�Zȼ�I��5�܈Gº��%��g��I�(ԇ3�\(,I�td�T�{>�u�[ ����u�����j���AJ2XԹ:�([i��s4]_eR��Vg�wˏ�}ԋ&r/w �cFD��l�Պo��E� ��A� a��QI�Ԏ�TMŃP�Z��]����sc����ė���RA��3��)1���bhL��V�`N���`P��Oj��jk��I�ڈ���'z<��
	�8�]�tc��[�a&�!K!�#��Q� l�o>E��3�>ʣ��P>�E����OJ��#@�� ���	`�v�=��Z;J��o����swQ��}sI˜�lwU�Two7��eg���+�1�t��5�� s�������\���9�v�Ա���f����]lB�Z���쇧	O�Ҏty\n �M1^�y��+H�ɫ�ʪ��aB����֫�F6*C���/�)%s"�<�����z��g�Tx�Y�	[��^exmel��F�.���6.!�@���Z������~�a���Ցv�;�O�?�>C����Ew�n�\"M����;a'���UN��`�)���f<�qlc��"V2ysЇ��,��#�r	��5����x�I�c�z_��H8��h�}ߏ(�57���(D6l���%.����xy��9"#��}m�m��R��.]{��e3���_����P�2����/�`?1�\����N(�I��������c?	% ��e�QY9�����m��b)�cΡ�{3J�]W�U۾ۋC��r�B������"#5���/,�uX譧���"�_������J;��˭{5���d�n�̜2�� �H;���_�x�Y|���I0 M:]Vҍ���}&I<,X�
�$[�T�9��Z%S�����O�z�!�pO2���J|2 ͈�;g,�8���5�y�o!L}����<���+�f�/�[�A.��i�_6d�D�|҉�4f:�ԫ�nkb����r�3H9
����w�i\_���MR�>!'0#zN2v5�8����$��(?����Mv��7���"�Ł(��Ï���4]�HO����L��=�� �>��P>.æKT��rή�����į���Q?�팹��G�OՌ����.�j�5v��N4�ș|	Mv{��5e^N.2�2��.$,i��^=| ��
�sI ��O֮�?p\ő��J�Bp��㉷��F��!�:3�?>EF$x��:�6l�b����losw?��?�y��x�0�]���]�����cN4�<@"�@�pS��k)@�����)$+��;��I���|�|�� "�,��W#qX���A\��S���򀒿,�lAYZ|�$9����O� ��������[G�TfT	�C�T{���T�J��.���IL���u����MGd�bD@���rڃ����祺+6���ė��/������b��Ĕ���E��� ��I�� 槹�m?a�[?����Ϻ��=�ifXv
�Yr9��m*��$P��0edq��?�C�,Ư�8$�p�oZi��#s�z-���&����18[�X�~9|�'�0]o�s��"����$6ߦ��\F�>7n�z�i$%s	U%*���8ҏy)��t@B\gH����U4a�4@���,�g����,R��V�3�v�OZ9�:���!��a��+�PP�fr��/��Kދ�v���������L���X�������{ �bZ����pu{`3�e����9��(�h��6}�!�#�c"m@r���c��*C�O�����<�*R��P�j�/;io��Kv�y�g���`I���)�{����K����M(o�����ϞK�fF��y�#VP�� ��e�C�H��)�^x/N�L���3b�QG�����ߊ��G���qvZ� �K?�c�!��;&!�{Gny���ʖ��;P�+̀��o�K�7g���0�g�����D���\%F�%��؆ +1LÜpigA)6	
��"��g�� 6Q=3u���X�I��NĮe�Z��X3/�l8ߪ~{Li��H���e�����K����h��;l'3,���'��ϔ4���vX,��x�f�t�6�(9SZfNM<�sX�k-0�]Ǘ������,:h�Z���d;�z�i�����������{�B��D���%<�������`���gW�f5���<�o��˽�#e�aR�3��1�FE�ѳ�~fG��%\:���b!묣Ot�)�-����E��<����_���'7��BP��Q橢��_R�*�e��z���\��lЉS�k}�_8���Z��� 	WK������_$�W�����ق�Yr������|�< 
iW(E+��B#WP]��tU*�W�A�7�Uӟc�}l�r�m�֤���Va//y ���~ȇ�bY�ۚ*s ���v=ν���.6q��z�6:�֒|���BX�>����A����~�*Q �V%%-����s�i��Korh*���uk*�F��a���dE����(�` �a�������W��h:����ey��r���G4��|����o�1-B[����A�C��4`����(���6�`�戚����$�o�>���'\Mt��8f�@�Uٝ�?�1l3�7j ��䩤�T�E����(4��Yv��0�2@r,� ���-2J7��������Y{*�@�O3����
�(�Z�jV��=�X|�	J�>ưf�i��g�-��l�G��ig����ۋ��-��k�����NB@`X\���tkoa�*��)��oRE�,�/���(������>R8�HlJݸ4�C"+����S<`�Hʥ4p�p��핓f����@-/��4��G���C��]��z��fg���	�O5b�C�ev:w3���m�}���~�c����tF[.�ۜ��V���|�� Kq�%Q��1�����'�$#opWG��I�A�U�Py�3�@�]~�N�"��@���r����;�fJu6)�,�ʐ� ���Y[S��XC��F�D9��cL����t�1k0'�3�R���(�Q�oͶ~��!{Mժ�:���46�֕yH
�|�|�������v�R�6}!m�⡋0�y&�K:Ư�i�-���9"r_4����m��o�����Q��}���A �a)�����r�&�&v�@��&�KG�F����Mbp8KS�O�z��0�he����N��-�9jHV�J$��:S�4VԪ�~�ѫ�z��]Nx�����D�g��ޅε��ѻ9�7C��&�vxݞ�%��ڥ�^�@���ϝ����NЫ�ƶ���W��Wϩ W7DY�B� Cd���;#�A�P8���97�"�P�:�r��
����N����*�sn8��2���"n^�0:�*�S���w�v�!d�����0˹�h9���"j��b��AA(�;Y\k�����\7�}�.���9�|����*�R���~�+�+���{)V�m�:ky���f��W졅�kO��?��j����q瞎�&A*}�L_�k��3�<9$T�,��U�<��.O�T,Yj���}:���gԮ�4}t�x;�l`S!�x��o.Ҭ�&L�N�f�gi��h�2�:�O��=D<.}�3��~B��)�b����J��R��n�[wz
���]��aI"xJ	2�!��$hgw��fo�,J<;�8��[��f�h!�T�[�p-ub��\,9�W�Dv@��Y��KC%O��z�k[�b����x�(��=D�w�v:�v��k��@��t�-d�n�R^��D��I�j[�^ܹca~�X8O o*.�c1FbL��D����I�\G$j�$7��;Qģ)�Կ��Ш��>+7-&�6a��*,@8WA���KkJE߽\��vz��r�	�֭Y7Ψ!t��܊���sf1ξx,�1,rk���%�E����E�\�����SRztb_ȖLX��5w�a�
e�&�Va��!�eIK�/Rp,����'vx�������"���:���K
�o���G�U�)G��N�PH��ܻ��c���0�K/��.����fh�c9�݁Kl}��E$��3@z����׭-a��Y^b�jx�`%;�{pL���%$�f@{�1���������}� @���Ž�� �%��a$rK���I�bK�"��٣�GƺS�'m[����K�3["\F��>�w�3(o��h�:�0�Ǣ1������3l� �ŀ�O{-2�(�t�����q�5�Zq����(EȬ;:�&�w�}�.&��$'Rk ?���0����R+8~ LJlk�hY^�F���ȯ]�t	��������M/�*$&��2/u�;>�[�gХ�F�T!ƈ>Hf�/��B�����B)��N�S�S��N���v��E@�]b��*��muۉ�(���T�ߛ��"#
��y�����x?��a1+��qce�T���xyt+/Dl��x���L�
gOlh�(�n�-%Z�����YM�R�4�N{c��A� ƾ��}2����A&L�A;�%�l��5���F���cΔ㍐aTdE7�>)�cI�ڄ;����(�H�QH�6�H3��� �U�1ˉ�w�ƾ2Ak��X����+����X�^\��<��U`Y�>����Ba!HA[���L���/Zs-��{D�X�V����pH��ϴ=�H�)������ـo9����(�'���Tdd����"���ű�˵@�J�F+�f�/F ? ���lN!u �(����lp��v�x+�g�yO��,�@Ƒ&?�cT,���fBJ��l- ��-�/�\��w�����V
�Fo���td%�z�u�/���S�c~��}8��E���C!c���%g�%������5'�]�����e�W>��S$h�cgo��:��Ow�W��;�Ùᜊ��V$��㎱0v$Qq?Q��,,JO�$�3��%`[���h*�X��i��d3����4
c\Z`J�H����h̕�L�2Y�7��.�Ff<�U1;K9��G���st�U<l�z�=���j�5�=YLԺ� ����C��4�c��S�P�jݙ��ek��A�A�`!�3ą�����!7������=���� �#i�T�� μ?c����AX2�F�E�6j��|�Hl��UjCwN�������Q?���x�EQ2+mAƜ�,*#��+��5�cƮ���iO>�t�&��~)�1��Ş���c��J�C�
D1��{��DcZE2��d  f�̞r]�J��W�ev��yRVC-���&g�d>��%�r���p��g����'�#�>˾=�
���/\Q��5S����[D�N�=�$V��V�B|׊4��~��yb���ό�du��(Y�C`ق��zJ�}�R�6�4���	�|*#��r�X�E���T����]�'��||K��P�,��]6_t����Z��kU+@l����+@����E��������L��O�#
����-�TF7d��	����ce�ٞ��zw"�Gc'=��t�ubZ�d�2HYǙ���ߜd���8�B9	av��?��:������
oËKX�a�l���&d�b���b����Y:�5��)4�=��<_�����g�S����Ԙ��_c� jz6r",!'-�-�����$%aSgHA��V9N&�f��|�F����R�[��b��	���QϹ��)�3Yb��g�O�_�^L/�=K�t�4���Yg���xOTXyn r����SCݫ�4J��"���d{p�d�Π��H��Q���I[���A���8��h�mI�}wB�����4���R��;��y�$b�������n �Z����(�3]���Fn����b�E��j{�!�h4�:��³3��z�qQ��_�%\�@s"��l�*Jkv;���[�t��~en���Ƹy�w<k�C2a�aQ����(2�#��K���3�1�.xU� ��3'3��N9��2ǽ���d�h
W�#�/g	�_F�`ݓp��p��3c��>�GQ�J�YY)����3��P�� ��2+���,<���06<I�{Ё��PP|�����ºD��viJtKcZ*�P_ku@��k,*d��[�QKA)S�	$J���Ku�c�F4���d	:n"O����@ĕ�����>��S;T�������E���"����<#�O`��K�e=K�>){�	�Y#-��9�/.�]%ͷ>��|���G�4.�y�������%MR��Ri_7H"��1�<o�s�j� �%b���8�-�TZ� �U�C3�$.z������1ߍ��	s��U�K��;FB�B�X�*��,x#D��&R1��j;�T
	�]��3K����G��n7�៘iV�I��~�qnv�n�5�/{T�x9۔�{+�wf;�Z1�~[t�3t~��}��H��՞J�;��{��I���Q�d`��j3^�o��d[w������,��%��>�������{ ͫcv��ۭ�R$��,*1�/���y�2�$[��:;��;W�������|_�g��]ÈrF<�X�[��9�!�ȇ�ܠKˋ]�?Z��&,�$���%@T���������_g�x-�a����G[<۱Vᇜ�C�i��y>$ a�3��bY��H�=��!�Ae.���4X���G�ˌω�{�[�AA�C�Z�N���ɷ9.�ռCR��qU��9�7\
�t�r��[�%�ޠ�34���c�'&���F��:km���@%��Yov��h��ᔅ���O�-���ޕ0��39�n�(�j��IK}MQX�]����Q"�����
�އrզ% ���n�I�V휰�轢�J���Y}�f������r\̅O$4"܉͂H�;�q�[F޿o5�N}Y����w��/~�e����Q���S��/ވ6�v<1����V��l����j�N��Nߤ�LAUcf�r��
Ӑq�\K��;��cf���0_�j*�/j%0���$"�	�۷��$p��g��V�4dT��S��xk���Nl��������H�
qz�Y�]���x,F�P
��a�pg�?x�¯�,�_��e�(?�'iP6���e��(.��b9{�j�[\�a�����+��XQ˨���I���i��)�XM�{��!��lK�a0�օX%`bj%w�W�(��T���yNm� PUxJ�
��?4��2]3?���(TPT��f�N�¼��l�n�������'�
r_�F� .!	ۏ����6�d �[��0���%g:%��~-1��4���g�FR?=�ZY�`�Ű����������`��8}ߧ�~�6���[WЬ �/��fBA��AдsJ�8�N��bN�f��+�1$�=��6Y��pY�&�S�7.���$�q_�B�G��&�EQ�^��݊��H;"�.4Z4��܊�k��<:s��]t�o����\�H�QaO�N�K��\o�S���[e�Y�E��̙�=~��bvU:&0���;̟��q�I�ƨ�M�Bi�,�j}���9G��G9q��Dq����P�
(_�����bqH|J%9��k�qz�����ڧQ�\�+�\�� �e7��I��ct�r�Hd�c66�A��L^Ub!�<O��;�p/<����О6�C:@i(a`<k?���y�<�n�ƭ��ոyZ3�^q�h�]�*��D�54	1ؗ;F6N:�V���c+�.�7O!M�����H�tC��Fg�0����_�vb�L��m�����BvC��e �r^`]�ѳ��/E��-:�~���r;��y�p�[z\\뙛E�+��O~�1�
���6g��$�s�y�`�{}	q;�[;+T��}�sU��k(��?Fz�?�c :�/M��.�#�v��!����I��p��,����g�eLg���T�B����2�?\�7>L�Uv��?�N�m�=U݀��]T�S}��1�q#�'*����la��~J��L;?�0}���D$nQ$����-T�T��eu���h�����[ڏܲ�� �9<Ԣ�*n�x�Br��7��auV�-�l���:��o�s�i���$g����ۆ�9� v��H���X��WQ�Ap���J�˔�6��D�C�\��qg�z��(F�U>�<-�������;lV��S.xrs�1��Z|כF������:/ �57��W��\�Ap��C����)p(�LX����I4�p1SZb������Л��~F&�ȖF^�� v�O� ��`�j�+3F����`za �j�"��[?g�&����O8,Q"\��2�֔�IY֒(������jF�m �E�e��O���'�U�+]^�4p����0���]I������[f�̍�6Խ��ԥ:7Je�i�S�K�)1��ݣ�~��6�&�y	��I��v�-1?T�����3D�c��9�Ig�Li���B�]+�2� �|�317�n��*�j�DX��l���zȞ{�BM���6�tbY��k*����o�k��;���0����B<���aK�L�>��Ц��02����c�k�6�x�gwS���8��Q���M	'*uǸNE����XD426x~���jk������4=�>D+ؓ~W��P��/dȜh���n����^��z�V����L��-B� #vOb-i`w��|�� (�Pzw9��8���R�{F��i�����KЗ1�7~}^"�7$8_U�ke�_�SBU�4�m}cN8�QNk4�eeϱˤ$��s8���@�|��[��wF.�����h)���6o��+�1�~�_m�.��c9�L5+���FKîC(��MlW~�@�T4���k�<P��׳��K�j��Vp�p������4��+@2�^�h"jsW����3����'�(`|�lo��VA�����d�i����æO�ī�En𔼬�R2d��ߔ�5>�ֳG�����O�w��v��eJ��LA��|� �O	I�y���9�:wʱk2�-Iu��7�1M~
�� �U�`��M�O�}(/��=>���1��P_�G7zP[��z��6Y��hN.0�����D�����{Ȃ�&Q�"���at��m����Sc�;|S��ӗ�P/NW��(z�t���͉F{YJe�٧�%-���|H�66��W�tj�$S�0#]pc\uLA_��sά�IQ���p�߶���Y[R�蘩�1���5U9���[ +��v�}��r��|�4�<-�l� i�A;<���3��pZ%�)�2h?���ǁ�?jp�v9,�	A � y����zg��D����1��n>���E3��	1ּ�� ʂg�`Q��:�y��A=w�#3=��7N��N 6�'M��8Ȋ�u\Ff~��G��̈́r&\*��e�t�&k�Mh�rԸ��m��p�d|��χ��c�d�V���*��k�k�������Ĳ���(TaC�H�pݒ�T~����k���K{}�ޘ%Q�S޺��9Ǻ����8Ky�v/��5�^��sx�qa9��#߳+ff%.��D����9)���藌���Im��
$����!A�ީ7��Ү~�Z��Z�eg��ش���"�� �y�S�؍a�=���� Gc��x����S�ħ�7�� �����tS;q�����gy��3��������a��Ւ��-U�@K24�#������B�=��Gk�='�J�л�*�r�I�rdO�l�{�:�nNF'�h?�h#TFF9lWC���f�֪k�"f�7X��,���M�Q�jh�,;� �7�rrؔ_�`��������"�#��[��!ҧa�r XS��(+�f�� .~*3��F�u�+X��s����x�'�棨'wdmjC�Vq� 7��i��3�}��s���UV� ��-�������\oR"0��֨���X++��t�j�[��ߝ�&�mB&+^[�͚�h�T��كE2�4�`ۘ"e]\'�������HT�=����B#�hjY�J4��|�N��&�s�ȉ)*�#@��`%õ�bKH/��lNS�~�XD�l�!��#<���K�؜�3�$RF�hM��4��H�M�|�:�5*j�q�=x/�y�q���L�7�#��<�q9qth7W�Y���yu4��O�m�Ҫʺ�a%b7���+�roM���z���Ewt�Pd@�vD-sV�\��>P0X��t���l���uo����߲����[O�ɀ�)�k�v����0������@�q�����V�x�E���� 6�.�[��י=�$hs6S�BJ.}�����m�7���}�X�]�;��RW�eb�|����6��3ˣ��f�L��������cZ�-��܁���|�i��t��ʾIw\��M��b	k60%�
|���-�f�br��T�_����>�		���r9�	0��ι)�Pȑ�5����XJV����e�Sf�j�7����_�����^[��c(F��B���
���ӟ��JT�"���w����dv� ϗH}�rb��)�����ϩ��w����i%�
wʿϒl3��A����_FC9Dx�v	�F�Msl뭅�m��\q>�V�2Ъ]`��M���s���V���j������^A�
G�`0Ri�����;�~G���h�lt��T��i��W%����˾���@�Щ[��5�������LmdO�8����{ D���y����_?K���(���ip}l
h�����f"[��v#o�M�gҩ�)�R��4�����tA�n���&2a*�5&$
�L7��ɺ!N�Tr�D� '0u���q�89�K'��`�}.�F}��h�Ns�F� i��[��#��=��3�O�O/@��X�Kf����ސ��f3O)����>�2wq�$~/	��?�%B/�5�4wc!QNbgƎq�W�OP^#��r3괏ت��,T{�2��^Tۀ����(БeZK������`�)�������[�Ke�6�&F���S˝`���5�/���h��� �N[��6�@��geSq �?H��IH8�ZA��h��SZ��I��c�� ېD�����1ԭ�H.ݟ�* :��pm���[�슇>��03@p�F0}�Py 2u�}���#��S ܰ�}*D|vx�����~�>�V#��a�8�����ץE��3�#����Ȭ������d����3�	^�F_�eg-f�����ܷ,g�}��a=~o����1��9]�J�-M%�����b<L	�C:"����u�?#��Q$8���1�i�� r�R��ڵ��i�����c�;n!
LrdĬ2��h�]Z̍�+���4�$Æ)����{��T���@�e��P`���7���yA`����e���
,��U����2�|ڦ�6�K���/
cUQrJ��JP��^�捪B�wM-F�b��2��#y[wO�dF�� e���?��l\�Bd��Oi�!H���su.=G������¿dA+�*8Dy�����Tٺg����|ڼ->C?�Ǆ�����fp&:H
�ԉEH��������tS�uM=L���R!B���-���X�yq��Oy��z�$ϔ?[\�1�%w	�O�O����<^���p���R���ȍ'Ft�I�rWkB�\�/�ލu���a���uܗ)s����.:��K˅<{|m����d����<�!�-v����,R6]#�t����=�����	7�i������]���D̄:�I��k^�#C�o�����!�ҙ�T��)j3��zA'�pg>��3��u��V�
]F�b�����Vf���5,��]#s��Z<	iu���?����]���^	֡�-�O��@B�6��7s�F8����d���N�1?����j�U�mפs>$�&Z�S�Vn���M9�BӁ���ɂԎ�U������L �sq�B�k��Ϯe�Ֆ'Ql}��XiGu��?����Q[,���z&��!�JN.���f�q����5���O�L�8��"�f�i�Ө����0{1$���SPSl�N�<:S4�;�mw�v0�%��UBA+�r��c'C�_�_sڤ�8�2~
ل���W,��C���G�U����@�',f���!$w�jN٣>;)���k�z/�J��̊��Aϙ�kƚ$-���&WE���)��O��ڝ@�g?��sf���Ji��Q�E������m��r&�rm����]5,��ԸѬ`�𑝁�#U(f�9l��Xu�(-���7
y+����y�'�����x�GsE��� ��%	nPΜ���A�30��4�A���^��>���n�ăO5��".�
4��9��/<��m��Z��L��m�%L��q_^��B�����(���~m�����<�j:�n���9��:�%��^�G�G�oJa�7f%�:i��h�S�@꾒����;%F'��i�Y���Ih�Tn
�_q��$|t�11��"���[�o�q��/9��Iq�34{r"D�9-�<�`���
�ܭA�Nv��~�T������MCd�"Dnv������a���
�RmQ	E���ڙf:u������$V�=y����j�C`bN+�NERbv�W�T_�cϤA
.�5�M!�܅W��KP���a[UB�$UȐ����>
u��VL�JM�rs|ⵗ!�d��܍�fi׳��_�7�̓E�"������`�!�� �9���n�|�~��A\�K`�F����L���8!Y�{�����ݎ���s�%_�gF�Ue"V}\s/��x`r-���,� ��LL��mZ�6\���(Y3����_��Gk�s>���3�-n�����0�G:&�>���#?�Z�l�<$(s��Q� ]���~�����w�
�T��0�ʉ�F>וT�5p4� ��#(��pW�z%����~0���u3A{{J����)$��y�E�<�K��-����l�m���9�f�e�׻p�, ��Bm�0t��
9W�{�k���dZ�F�jdl�yjG��Vf�D�LJg�-׻�`W��c>�Vg!*?�Z��_���m}���xe��a�F��������G�l�rUR�5�L��l0ȥ�&0V��s7�1^�~�bJ:ɨ��Ꞝ#H[oC�'�uy&�ls��_81If��F�~s�u(pቸ�M��5C3�Uo�Hb��-�����'�#q�}0��K���T�՛l����cYl=��j����!Sr��;�k:��F��p�FY�O ���î��,����S�@����S�"QQ��7��l
�,�j�l4O3l�dLW�Tp3t�V�2��9W.��\w��}N`�4��K���C��d�&�	�b8��Y������g��~��sWf?�ߥu�;yn4}����S���C�[����a���s��"��Ndg�=�7*<$�����=�qj�l��ѝRG4�EV�5/��b'E��.F�#,��bEu�WB8����s�xe�70�����,M�u�;�n�������}�a����ڗ�`q���{�1�#�<p�2j
�Ȑb����N^6���Cߖ���K#��ӧ�C��� #N륜t�L��Ẹͣ�s��ᕸ|%����;^C;A��Ǻ?���DG#���%�`㯸�t����}ݘ.���*%>����'xj�"�X�.�&�/���=*
E���[D�^�q���͙ăJR�N��(T�	��p@�kʤ� �Iw��j��)�uZ+�F;�7B���m���h7�X�ͩ��U�ȶP�tŏ��Hd̜YC��6��E?l;n~�m�[����D�KoCT	'���j5���ڴ�^6��k��H���8ы���+���$��}Mt��չ4��%��ڝt�n�"��$6�bA�9�5m�ލ����#�?
0�Z,ԋf��M,D�nF���uy�	��E��(�с)�6��o'H��,�j��`1ݚ�mZ>c�p��$z.�)�p�%�Caĕ�к;�B���ǪP�~�DkN��)򸩏�t���
h�2�,(��y��v�vx.MMl�w��R�)�17i��)]% � `�#��|������	�_hC���u�2o�{.-zf}�s3�
����i��/5B�0)a���9�9��\5�}!��-�>��`�z����H���2Կw|����t����%���˱�L]8c��&f��<L�_t�d����{�#Ĳ�����7��<�9ւwl�Տ嗙'^��98�5;?*�>�3~8�pr�T�<S��n�VI(�v ���Kzn�
�k־H�&uN�Xzi�7�!�/�ۡv��ڼ�ˍ�C�E8Њ�~_c�x~[�@8!�u2�t�Ƞ�28�x��^�
�SZ�f'm�;A�9۲���x8/\ΑU�v�R��(7(�����j��l�ț�Td�yZ����^"�!?�Vq�O\�#qfs^��Q��b*â�ר��P4�z%��*�p���O�L��y;-si-��if������kFwx7%r�GU�FN,;�z�X�kL���Ӎ	O���6� e�W�$�(�c����V&�Ƥ}=��Q֬�ׅ��H���3�B�u�8��w����׵$�`nu8�H*��TdJdTبud��!�kS/�� �;���O�J�-^{/��#w��y7';!@����/ۨ��w|}�ND�+m�~G�L��L.x���(����*)t&h y�9��r9�C. ��pA/�N�_�c��uZa��̎H��r�k
�cG��>4�^eA=an}��DLH�`X���ik�#i�e�:��a����U��/5=�}�������ӓ�6A���*�\iZ���2����r�͝��!�	���
afm��2N`aC�Zd�n<�����/���q<,����܆�<��Z��p^�v	e؁�B\$���=�3}�/�K:�yXZo�7e�Κhn
������ZQ�n�m�<�=����-������|�Q9�_��}-���l۞��2��[G�*��)Ir������~�U�1��	���c\�!&�S�Ky{Pz	��4���;s�����9׎�$Wt�o��?(��O�P���7:Ҁ��ۃ���A��2P>�s����<��֮%�c������:
`ؚ];�y F�On��y,�V�`�=�>gǄ@���|P�B� ̀9�"0�5s��:������>��52s݆|�ag�䕟�FfL�%������}Q0��[�Wdr�,�.��7Ҿ��)Ȓ������q�%�����pGi t�'���ˍ{_�G��1��۫s� AZ�>o��]T�>Em����|��̀�?��18�]	�����&G)�����V0cG~f��5�A[�B&蒛��+MD�6/b����L��D	F�z�h�i�b�Ϲ^m��/d�����-���f�1��������4@h�&y-��P̡2�"3�|�gj��N��(����iɇ��fN��
E�8���xEy������Hʯ}��2#,�$~8z<�2��[XI�M�� VV���V��{�ޱ^H�/O5jx�v,�Ic
p��u�W����̒�E|�1Η�J=��o��In��2Ѯ��X�Ӆ�jTiK-n�B��U��Q�0�R:��>�w�%:��m^��e|�eT�D	�C�F�|5���LO��KzD�v�7���e_9�)�%��� ��b9铕�)�L��x[t�@���ϤV��$G:b���V�8��g�3�"V�2���w���\$�隀v��%�j�04"�L�ַ� �//�� o�7&��5p�\���}/�x��En��mZ�����s�]# b�2+y)fy�Q~O	7����S��V��:�¯����T+�M�e��T'���.t˥�G�5
�_�9�EuL �O��y_�A���T,6Ǖ^�����c���4
UG�"ƴT��7A����;{��w�u	��]DFD=������rξ�O׷ݯBQJX���7D1�3�����1u,��I�h�6�N5�kT�`�n����?^*=W���kS�:�ߥ���gb�+��M0LܚR�ǃ���}(ـ����	�+@B��8[������l�7�w�3�!F����q)sR�Q�H��h��*�l��3�n[�{��\���B!'�����s��CpjF&"j�x<u��Z�!FJ�������ɺ���|�5�ȴ35�n��(iVYrx�F\4w]{?W�߈B��-m�
JRD����1��JZ<~�>�?�0#��F��'~�}Rv�/I�Ӏ%����K�r|zA1��J#�i�Q��0�Zv9�ۀܫab3��	V�xK�f��e)�m�kM���6��EC�{�2L��",�����S9=`�>�z���T��r(��a5��G�I����V�\H���M~:&�rA8�=����d���~�%�� 46��W��:���=�����}"1�aq��8�A��饐�SY�o�[`GL�6/_-LƵMި��o��RC�B�����g�r}��PL��wA�	u��N��a�lEB^��}Py���_��
@Y�X *�KŨ�5��I`�+;ߛ>]�����nو<�0+/4 /�ȉ�68��cz?���Y�����[OE��Ե��C��s��iGㆇ��3,�C�,d�L�Sls���֟������t�t�=�n�ג|fc��� ��@ !��M���D
�Q%��8*��,u~�ߔ�=�d�[���el+�>�`�l����
��j�/��Y�hA��b���1�jL�߸��V~�ƶ���q]8!��p�g��wrX�Ӱ�$8ӥ��l����@[U5����p���T_�)b�ؿ��j�,�/̫�N���i�l�D�g�k�� �B67�����H�z	�&a���O�M
����]a�jMY:�(-��Uz�}��h��U��ƺ����9l]��\O;��)�EE�;Q.@)q�g�#A�hs�_a�Ԯ����0q��`#�0�ܰF��`�$CG�l����������p�A�V-Z�:1�)��V}�v6]��T7�Tf+�Pf'{q�1��t��Q�ڙx��3�nx��M&δ߼�9>�����ڽ=W����W�O���^g�HH�v~�R�J���l��oUh���ћ{X~-�
�R}�Hu ���Jnt��}G� JN���}fCwx�����]{��3&3���������[ß�6���Ri;��#mB�(���$G�؊=k���H@ ����$��h�|E�*P��!�6�7ئ�j;:l��m�Rn�Z�(�����J�[f��h�H��kc����a�-_~o��?c�ֱʒ=0��G�{�eV�֗��#�j��4���$���6QrrX�&Q�OvA{�T��n7 ҽ 4���&�E_��~���UԳ�Vλ����c)��'�[������Xs�u7⤊��v?y$e6��J��z�"��v�5���xI$�@^�Q#!�LF�.Uc�BnD_�-OO�t��.�9��m�g�c�S���sk����W
��}і3E!�l�]fY�M��xuWU�{I*:���l4[��U"j`���Pe0/��s8M��	���f��~��`l<��;����B��*R^d�q��:�?�l{��%�X���Q��)|�%]��4쬌ѨT� ��"r��n��L��ѱo��Ɓŝ ��p-ϵx������nފ#:�/�qFti4O��Y#=3�5-L���?��%~:ebi����\���+mW�y�<`鶙R�1'C[�1f'��wk�O�n���{IT]￘��\)z��\K����OQ5�0:�N���n�+F���~Z���_���ѷݕ������7̅t�g�5tNi����<	YIn��;�'7�J�#�j�#�Ti���6�]��
�=�MG0i����2���V�����,���Kf�6��@��nQ)��_Ư��j���z�f�l���E0�q���?������ħ�yPX��tB_�L[ߝV`%��ʈ��66EK8�����9��G�C�A/Lóۍ ��J�4�
{�F�V���S��%F�j-�o���1�|��g�y��;͗���Mw �}��Mp�Csʾ ��G�j,&[��W�F �W����o�!���ҙ��~GZ��|�ǝ�:�j�'�5ed.�#8�M��M��+�F�J�Oi|��@�Ʉ�1ɗa �щ��c����w�ٳ;�+�N��B��[jm/^�*�w::H���.�bݘ���x7w�V��!�A��=1a�12����K<P�s���+e^.J�O��u.�\��t���Xc𩧥Ҙk�{w�-6�%H���&'m̀����������,t��۾�-�W�[ ��$�w8
���:=�n�FQ��Oǅ^f'�߈��%	'Bny�����rS�a��M�����%�����\�P��	��
�E�"�/c}k���@���'ɑ�6��̮U�� �k�|L^��Ԩ�
�.�56��3���H�~�.:>�5�[�b�������}��I�+7}�w�
rEfddi�ڢ�~|)�D�Ċ��h��/�u�7|�KrO*"��㪞��a#���?�A�~�Vˀ�^\Q�;C}�,����6�	��0M�*��"�=��g����Yޱyt��&NЕ~�<>*��#T��ke}���J�L�=�"9l���ذ�~ p���f�y���ģ^
�9�\o�)������ߪ厑[�L��9>Yt�p���{�I�.�7�A���Fwò�(�g{	����x�� �����Q[�oa���ć�#�ܻ��z	�����3J���Ji߸��6i7O�y%c��Z�����Y�����q�n�4�s���S��3��*_R���,��m='�+�[8��J6ٱ�3"ɢO�%� �<�CP�y'Dm���qI�S��*��<%��"�,��5����b��}��eұ��f��V�d�]����6�5핆.�BN=
�������#=� p��U=SaU>֋/��u�����_���e�1Ӵ��	jh�/��5�rǂ�kصJ�x�h����n`��o\�������˨�:G$�Ki��(�v���-.�h�T�!�jn��a1*��h��|�L���0^S3O���ߐy�a)��b]���[P������Y�z1�*�d����3��ܺr~c��H7��mf�IM�3A#N��S���_ao]�#�J;R��O���b�+U�-��}o!�
��K���OO�_���A9��^T��M��lR�I��N.Ce���DW_t���k��{X�������Qq��b��WF�X��Ɨm9z�%^����&� n��'��tz*!,�� 2�f�}5�A�ͪ�o���g-|�0䟲Dm*w]	����d}��>|Hu6T��A&��Qe��N���vuO*��`qy�Ɛ��/
�4���K`M���(�if���0�"����R��ҙ/� �| Yd�+�=��7*���4y.��Ic,�<�9�u.b�X���A9Ab���NՈX��a��N:��A�����%g͸�-�P��oS��ܧ��pjt%�l�{�����d^DI k^DY�}7,��<��2�/o��uylA#L7z��$�;��_�	x�b'~o�U�q&B-*; ��y�;I'D�JeOa����BƼ��'Ѡ��ǉv�\��τ|�H�p�@J�#<�@�'��N�;��x]�*��Gs(J�
.I,�]�o�gv�Awk>�1��ye��D�ٶ�����W��n���#�הQ�О�%���{#h��Ng��$|I`�?�T�Zq=�%�ț�/���I��'�����g�+�(��Ç*6~���}����2@�<�uMj��~��Qח�j���O|u��.����|��}0NDp�s*����Cx��p������(c���:o�=�֯��ۛ� �[�^dc�'����z׃��O��0��˥m6ܖ�_�`�_�(a $B�&Dd�	�A� MT��^�_�%�WyӅ I&��f�m/�q���<3Qy��m��\�~�o��Y�Tz=bΘ�V����G�;��
}�u���^
����DQQC���k��`�U^Yfp�ۭ�8���^�\,w�_�iLs�6|��hca�8�9�͸bs���!!ɶ҄�M�\Zr�]�oL?�Ҫ,�[�d�Xݎ
΁P�9K���ϭ�+��ES�{�{�ԅ�2�87$�F@�o�7�L���JzN�`d^�c����w��(<�(�~ma���آ@ z�D&P��;���Z%����,��������ab�O�$v��aT����$r���\�
��h]�����*6 O��u�柡l�h��B ���x�K� �H5�F0$�x�ix�?kHQ���F���fn�LqL�����ņn|�Iϒ�t6��7���$����Uq���ՂM����nw�dan�RW���.5����6�Wx��J���ucG�\l`�6/2����+�6V2yҷz�H+���2L�Q<K�r�T��O�����3�%�� �a�9ٌ�6�P�_�c�fv�����`���3�h�K��=�`	a�D� i��|��P��b�\�Ɍ�ŏrB�cɃ_�B7E,�����@�_��Dp/��m(�o��S2� ���/�i}��#��s:�W�qҤ��{Ap߈�T6%�*���k㩇��}x�w���YM�*�@ۊA���8��Q�X>�20/W^�F٠�&]�M_ˌ�@��k\A?+�/�M�8Tq37Vr�71N�.���U�˱S=+��W�:9���Ei��=�x5Au5(HgA>5ڍ[���S�B]��
Y��dT�u���ݨ�v~��9�#-��ޏt1�Z8rI��#�l4���`�����_R*|�:Z
��`؎WE��a��o�c����j�h���fC��#,��|W���+,���$�Z���D\A\�U��M���Ǻ<�Ľw�2�}��������h�\2n��&�/����h@ҋ����y]�>u��	�A%];0I�.p��������v�ˆm�PؼQB)/����V3x��5���>s���y�X�}��h�81.�U���P,Z�x��y���.g�O3v)\cᦹ�~��UUC<�%�^��w�����3�(�y(�x~��p���;��&? ٪���ǦR'DX3�_��怊�j��:���O���(�+���,�+�S&�<kLJH#�Bفڰ��%'�ߢ��2bP�MY�&�(j��L��D�Ê�1*)��4�GfK���KN#��=�N&ns�~�P�K�5���Œ�t��^5}Ũ��9 >��hX��Z$_B�
�}�E��1��(<��pc�#>�����v�����S�m	�F_-\��W�v���lN#�̹2aU'�#�gEr펎}�(L��'��r����Ag�%�Я���s�Qm�ʼ7?�	K� oM>���q�%a�=�ً=�q��P�m>�����-��%&:P{;�.���G[W��V��%M��C�LC�&ۘ����AB���c��)���8EK�EF��� ڴg3|����u�6���G-*�m�׆��N_�ʍ�S�[��o>�X�DC�!V�znWub 1�]���ﰖ�����uns8��iq� =�/O92|���N@<�&�(6F� $�[E�%-4+�A��h�n�G��#��^�xj�U�.Au����zQx�ݍ�GU���c~���"��@�9bxq��P6�3jt�K�o('��Ԯ�� 0EIw_�,�:չ��B]X�Nh~�]�PK�MPȧ��Β	G�J>�_'.���k�I.��u��(tyg2y����]
�FJ�J�vGWhx.����׭��ǽ�A�JB�c��4V�D�(^O-ɦ�bKx P���<�c����_�%���,�ɋ˚�P+ ��"Sh>,飀��8�bC��钻C�`��IU �����[��H����!���na�3�f�D�i�I1V)o}�L�P��PI�h�wj�<���)��˩������,)bi��i��)��q�Ó{�a���b�>�ԟK%��h{���NS�c�IEX����	E���yo���.�y-������+Q�����I'�}������ܲ0Ln(Wt�ѓ� �=J�#�b�lk*��<�e=�������_PLd��^dS�Fϟc��	���@�;9,���8�*]��ʟ��N�R�6��NS޽P_�$��^��f�v8Gj����KƄ�q��9���Y�M��~<�2��KH|�1V[��I��ݔ����[�9�x�P1~�EG�?�ᯞ�&�~�!��{�o\3���)|�][��Ɓ�Q�,��d�vIKZ�]�&�6�Ύ.���jB�-��p�+�����=������9��@Vk�˄���m�>���E.D#�H�.@��O8�B�<����ޛs0,���?$ݪߊK��l��l��7��V1��g(��Wk�ls񵴚�ݕv���ܰ�ȿ�m$�.�DEm#�ϦBS&����"��&���\֎�F#�#(��K]t�{��̒������]�ӘF�(<$��`������s#Ky=I�"O��A�蔢� ���@s'+�@�nX2�{��E���D'�F�����'Rda�^��Q є�<��S�H�j{C�?F��hp-A�h��!�ɽ�|-0
�Q�\�R���dD�(��K��Q�!++G�Dm
���W�r@&c�2�B9<�8aK}F��,s�net�V�L����	c�<�aa�om�����H��-n묙Ӟ@s���x��Y�f3l1�ʽ����l�c.yrs��{�/�z�b�1Y�4��� ���`���W[�ˠ�v�8jKgy��FC�E�� \�*98s�I��G �C��p���$��-Lt�5AJ�6__�&�.�R��䦎���58M�d���%�ɤ���f�Dd�C�@����x}՜��DSu�r.W������HY:�+U��l����ǎ�Rr�8B�j}hW�?�|R��#Hh�It�e%c�W��yG5��d-���shN�Y��6�0}��L-�oJڻ���N�3�~�6L2I>���n�!a^�xh���L�u���$��@��2�4��6L��4��p��Disz:�m�?�����F<�w]�_�B����u�+��l�����huH:FL�1�������U~����t}�	/����5 �'� ��_41|�.~�.+pb.�+_`Z?�LQ>�t*�R�n��Bb3iX��.�8����f':?l�9C�Q�+Y��S2���E~)��9��7D��N�KW�����Ij���@#-q��ʒ�h{k��/*$���+d��l�[�R���
Ȗ�$ct��l�M$�'��:��g!���b���]t-�ڻrٽ�Pz,[�J�m� �������)B+�&��T�:2�r��π8~Af��"JLi�	@0�+����ɸ#�l*��k[ f�P*�:f�Z%0V|��(�'Ӱ^#�k�`�u<�"/5��=#= ���hs�YH0�k�'� �|.d���t�bDw���~Ɉ�չ6y�Xƾ���G�uO���I�J����"�Z��O�ߋeZ�&�~�yK��4�J�8R#.^�8/�*�j�c�����8h��-Ć�~:O��`�'L��c������!%�]/�1vRLN�to��Z�o	)'*{�#���xT-<��#�Yh��c��-��P�i��	���.<1�	W����B:B��
���i!�/*�}�;'XD�d�P��Sѽ���|����Ϙx����aR����ϘO�8�Y���/z(��UI��w���d�9�5@�9���{����)�����i�B̞��+C>d�23.Db'������c��5�;�6��ܤ��ǫS�ɼ��0�"z|U4�`�$Z�$� Iz�K�����I��H!P('�gr 4o[���&���v�v�`'�w�N��|��+�����a)�2�@^�,�����Ԙ����8��1�$8�K o��B�cb=��u�I���*�m�Yy�ZCd^LC���.��D�"[�@*�h&r�J�-�kW�ԘI�Ե)~�4j�V"6)��0Y��mֽs����U("u�Eb��	�2Uh�����[m+�6�jȠ��m,�+0�����fw�Y��B��e�Z?zj�6&����?�:_o�}������<���S�������M⋕𼂝/{�F[���Ú���o���ȫ$��UJ���2.xX��,�A�|P�܁�kRS8�u(.�n�N�מ��K��#	/�@��3��:z����&�XE»�e+�Z��}��������n5|�a��6�7��s{$�C��ƈ��&�ʌ�l����w�¸h}��Y`���I����������L�QiT�)jN(h0�C�s�=��6ED��+����$Ey~Xz/S���5;0��J+���>��|f3��s�<��A4���?�d�eN#ߵz�I�'�m�:���_X��I��-%�(s�&�}V�	Gg��Zw�u]�Y{�z=���L��p�{k��'�|�t��pE��~.p���Bw�)�Ѳ;����.k2.P�̓�\C)�1D��no�O֜%U^��p��򼰂�������&+=�U��k%<���=A�U����j%[��9Ɖ���MgJ1`��$m�}#��%�A��+
z��f�r-5����*�{7��7���0Fԡ#�$���L�&����ʟ�4�a��ٯ���=� P�(���>0/6�,�l�D�`�E�X���OM4c#ۘ	7 ���F�~��nv�_.2M��<����2��H:Q�90+����8�F/bߑ|6���� �w�v���m|=����:g+#����8l�x������1���PہFI�9#��b>C}!f��Ń���#P��f�^l�]X	��.u� ����%2zmde�S|�����DU��:�T�M���1���S�}��!<U0��u�St��?�c=�B�l��*���|iP'h��i2(�~_��]�Zs��J�1÷̈MSf��J6�hN�����^>��A	��Hs������������NI�\A��P��d�K�
c����n�W(����dmHH�-~O�~��+DL>S6�8w���w�vA��7�K�fWxh!�&�|�_�]��#,`���:��L�Zhg�Y�eswԬt��ܟJ�R��v�l�'N@��~��!ǩ���;�r��xx���iՙR����}��+�ۦ�A���ٍ�Fy�a{�(�iKjr*(i��d�'�̕6Atǫy�p	��EG��k"=��x�����$G�݁A/�ª,��}T2�kb��*���Y6/�Q� cڄ5��T4_�w��a<�[�A�^��!ע�����7R�axIz ���e�j�����z�s͌L�r���GY�5���%��"b�Y3�
��:�[L��U�saC�ͺ�/��U������
`g����^���E������Vp�U��XB>K��ԣh���3E ,NZ$9~�Ѝ ��[�"�sk$�hG��V1=k�nci�:���,C4�X?W��
�g#�����H���^w��N�R����q;�#f��� �p/�%!>�����k�ֳ���@�|Ҧ/:�Tk8#(�f��m�:�m6sO��c��S�?��ȼ�B0z�yP�WL`&��g3���eM�RT�ı���OZ�9�����s�k�RM�Ҷjד���PP]�w�Cv�*_�M��B w�fa��qC"���������~Jp��
J�U��@�2~�ŁkȆ�<�u�W�	|�0T�IEYO�cm:>��K6!^͉h�98���k�V��L�w�d�J�Ϥ���06��"��姰l!�	Lޕ*k�[ТQ���# }��r�)`{�8n�"�,j��bg��m$
�iCu����-�����܃4r�cG������ea�V$MZ/��-%袻��b����G�
�끬���p��?�Ǜ��a�>In��x��g�'�����񊐕����E������.�g@�o���е.-�d{&� �up&��,"���4}Ŭ�2`1����pݩ=��fhK;��ov�J�u:�p �ת���B�Q0q�+cy���C$E�}�h�x�{x95��:�y����9g!`
�)�рq�ie�Z��K��+�Y㴚��7���&���tL^�#x?Y�?���縤��)�ܨ����:(��|Q"�L����Ns��]/<�O}`��>��ƀgF(��� g��zA�nF3�|s_r�*�����W����h��kB����ja��cG
�.��D����+���%���v9JiY� -/w��.����!Z�"/�.�R�wTy(� g���r����c�N~�uW�Kc/Æ��Zx�g�I��h����
�[��B�Ė�����VP�sk !tPu[t��L j&���g��@!�H���
Em�fQD,3υߋ�=��
_{�R��J�[�y��>�jɌO��h�4�;S&���-J,�j����6�;�X�9;��d�SB&�n*f�TM~V�EcIˊ =��:�����P!XQ�� �!�}�.JC]k*�;�J�v[�:�h�;�FA<_����Kˊ*}��;����rvQѴ� D#�g�}~|rS1 z1�#TC��R#/-�L�5���{�x�ٽ|�C�\LTy�4���r��=iI)��Zr��
{���X��)2�Xw����Z�^�1H?��GDO�,�7$���i~�][{��h;����dQP>��e�-��Ky�OV\��2�u�nH����!�گ�M�FQ.Z ĺ'q��h��S����|�Ĳpؙw��,˼�s��XD�?�D/�aڣ�ǒؿz�2��/���R�H�c�ˡɱ���p�(�djA��`�i+)c�o%� ����ɾjAlƊ>�&R���G۟�(�kd�J� �7�ߒ�8�e4�\o
Ҥ#�j�;t�͝�����Q������_��`Df�I�/��u*��{����.[�M��s�<'�x���h����f��ka�������R�G���.,�H��P�뫷�ь),I�d�:����˗[�;���45��D���c ޶ы�>Q�2�1q�����`m�R)$h^�t���B�UOMč�L!�
WX�~���F�Y*A��e�yn��	�񳷲y����X�V��yX=�9�O�U ��w�ʫ	�t�'�G�|�-P^��))�"�.��N�6�ZT����kW�G|�3���#v�'pq�/.;A	��Z�\�A�A�O �E1Ė��Ё���NO����wm�ײ@g�2Ĥ��Q�۬�t�aIF�'�:�O�lA]��2I ��ojtQ�$��ך{�eĤ:�h��Fϣ�����)3K�2�I�}�j�m2�`�Lҧ��4Y��{�ɗ�7�=�V�՛|�ƴvQ���OR8�	4���n����;�̕��6���s���d]?��U�y3�5+���R[��\�&8�/[ڋf
;���vUT���o��u�I S�]�#���c�nA7?�[%E{`_z���1px:��oX,�놓�84ȉDڻ�bS�\�<H����ʋ�?�E*�����c��'x n��`�P�<SH&] �I��]v-���!��,J�����Ү��q�	���h9=o�7   ����P��R'D��Gn���5��tw��B_��NU%��u�D5�L��e�W���t?`>�K��F��������p������w]K�a�����R���D��;���4�{���,�B��T�l�=�,6�E3+������~��4��?]����lf@ňF؋�b�y�y�5�a����Oa>�h��C�.}q0�&��Df�:gz8 �	�sy�JҜ��� .=:�6>c�gp9���Z�y�d���,�_=\�;�R�ܿ%�\�g1�M叏�^R��!^X)�D���Ҝ��b͏>g��`�vuj��p�P[-׳Gh��ȧ��8{g��8�L`q�T�dV�Z�|
g�A'��	H���0j3�S�j(fެ���6 7d���NG,�s2�;@��5$�>����T��l1]�B�[��/��<��fd�O��B�8�&�S$�jR9�Y��+�/��jF�߲�KLCh���)zX�C��iS~C X�<�9b�j�_������ٙ��F�d��J���]"X�w���6�|uA_�ܻ���ੲ\��˵:���(&��r�v$�1+�N)/���U��5)g)�e����~��$m��)�����)�Y�����u1�&�ys3ғ�7���˖��k��<\Zq�ݤp�G��M͇���	j��r�<b�N�+(�9S��^7��j�?_�p_���u�z,�� tOٽš�Dt-�.�6�̃y��&L�+��f�r���)f#����m����JS{x�E�a�
||`F���8	n��ιB�����7u�r�)R*.k���̜9x�i��y+�Ey��;'r��[�<�t�z�	\㷔��Ej&A�R�Tw=C��/f��d�h3O:�I��u3vNLa�l�y@Vsm�u�($^�Z�y�kvDj�݄曮���Q_ѣu��&��"�-��ML~�(����oڸf�1�E�#.�I��*:������~�_�@������g!��������R�΃�x*��^�b�-��L����ϸv�d�}}B���kv�<�y���y��T����E��֝8�;:�"$�oP�5�����W�6�n.��Q�� �%o��J	�M�a���	�\󛲀��|�p��@L�g��{�@��-��ԋ㐜@�Ü,����s� N]��/��EK�b���8�~L��^`-����Dy�e+�w�.davw%���M0�D	TW"��:�e�@E�/��,s��_`nt��-J�C1Q���{eL �tA��[cS�<ٯ����Q�����h�q��!������� ��3K�%�?�{%�nJ��"M����/�$yO=7F
�2}.�H�&x͕�-����F\$�����[��z`0x�qa�P�����B�]f�� 㩒4�Ǜm�X���m�9g{�Db%l��F<�%Xra�-r�%4�m�vE+K��f4�}��iҕpt:��gG{�i��2�2�H�<�?9�C0�&4�pB�%=�y�hT�7~��p/<uw�B�AdS�E#�F��>�ϟ�P�i�ͮ�2ۄ��i�l�P�lj������]�+j
n�w7xt5��BQ�g�;��b����
v���'�X�gT���C8+XQ��h�������'����k(Is��+g��IF�B��rp
t8�X��p#��1���_�wI�'�R�Yz�c+Ac�����i���7�C�Yh�l�ФU&�F��n~���or%�!�d�˱ꝉ8����4�P�����&BML >�Oc�A��p�-�S�-:ᆜ��̆$����i�=y�4�ق�aG-�����b�%�Ќ�Q1VI�V�귄�ª��؁�EN����r��>��g��3�ڃ^s�ڏ��j�{��q�	��7c���X�p������)�O�c��gE��K��q'�X"�:�V��\�\u�D�!����ZP�U�����ü^ƪ[m?�suK�6W+8�Z�)�a�K�wu徕��D{�gP�Ӏy�i��=�lJ�^t�ּ������7�6�B�-M%h������O�S�{�)m�=�]QB�t`�������U�O��^�j;�tJ�
��n4m�jAj�D�q��$���ں�DST�$����c�� t�r�Q�/8Eb���� �z�?2��9Ɗ��߇n57^��c�0gg�@�?�t�iAnT�G�qfPY�V��'�CdR��]F�N^ɲ��M���=N�EӾ�Yy�j���-��P(m-dg#�":w���Bk���4W�we��k���E!�>N�Z�9�?�MS�r�ʹ�'���56EW.�
��>�S�N���UZ��h�q�$UN�Au�h�|\�� ��9z;_�8� �ۑN'E������	�6�}�I/�c&5Un�_Mb\��:v�|�}�*�N���͙�0���`3�x�Y7b2���,c՝�<����p�-���3�2Xt�~��z8�ބ��#jZ)�0�Q����T_��=��p~��o."�
��1�������v/)5%,�du�G	ޤ�zm��o�߁y��J[�|w���a����lq����QX>��l2#)�9�B9C��pp���\*'Y����
(��G�ʮ^�@W/���WKN������[v��YF��g���m�f'!nF�^����ɞc��i��Ԗ��2���|����z��,��pI�+OT-������ђS�k�u5/A,o��Z���X�����a�ᅡE��/$�H�LM/�1D�/�a����ψ4|�Y	�w^��� ��֎�C5��N���#�nB�K�v�ݽ��[�9�$��	*�Y��b�sw���ۥh����}��*f"M ��K�;���&�{�����5�1�ʜ�ŋ�M.0�%��ua�������vI�&�g#��e��OHZĬ�(}�}���d��dc4φ98�i�D��_(y^��'�n=�(.wc�Y��?pj?����t]U򐆢�t��w�	$�B�o�����S��>[��A�x$8ȗ��%a��S;�ڡ�������k�[�S}�K�Ȱ�Mټ�fm�*1�\:�XV���J������H�m8��X��w�O'ň��,��o�����v�����K��Cx=���K�Z��6��N��5"��{D�~Q�"�'�(jy��p���"�/���� ��qW�\2ǆ�Ⱥ�?��M���7A�(n�<� k�v�X��/�����="IyH�P�=��1�i(���G�/40�j�v�ӎ�r(���m��l�GA�$�� �?;&A1���z���f��s�- Ve��֔6�s��bgWJ���_��������z� �������[8V���_���Nmu⚪��-�:�&�	�{���E�����p|���@��Ա�X%8H��AP�O�K�򷦿|��c;�uAGH{�dS)Z��kTKZ�&ɮ\~�ڡ'���	*YTŬ>�Ԭ?���݊��Q�H�����-�p�nNe#�]��v#[�|,U�J�����v��#��d����d�q��DƧ��u5<H?��/���u`ܳ@/ޏa�)M�P�%��vB0��8
Aքj���d=)����ܛ�6x��������9;��^l�I��NP�a�l��adaG.���,���JB�������
�b�����a�G�#������S�v�Or�&�)ٙk�xw����@����R�]u��f��Q5�d��ߌ����XO|o��e��l�����l���r��j�iuOn~�BP�|\����7RC���^8 tA�xܔ������ݰEh-e�C=2�J3=ί�2��?�mP��}H��4Of�:��5C�bC�5�W&>� QR#j��� �w>������e{>QcHک�l��X�f�&p*�2�\_����������^hGA�Q�'�g!���}"L���RH��ܨ�P@4�ø�lNs��W��oKBe:.��/ZuL˓8w��Ԓ�\��C��#�<3�'�y`ҶtǆQҤգ^=n�D��z�J�
�Ч���U�nz�Q�#w��Ӡ8���;&�޶���7��7�V�=�fIBi��S�ĳ׮���`�J���*��*��Cs�,���<��u�w4�h0SW���;u��W�A�7����6�5��[�yʢm|RL�E��W8y�{S�pX���0RY�}
zˎ�6�r�3,�p�v�PJ,A�,�WI@C�`�3^�*�w�К�^��a�lLY)�{�?�rW��h�����H��0���J�d���ʘ7A�A%s^�4J��>:[d�V�fz����>2sJAP�K�Z�n΄�'��.���c�k�����Vn��}xR��(I�>YT���ӹUv3YD;�;�a�pβY���Y�C��&Z��ox<bq3=�.��5s���}X+f0v���N���\K;F	6��+V�a"�(9��P�����"� ��L7��vJ|p��p�|Qk�X �2s�;��I�\�S�~Ĝ�h� ^B�Q��D�6&�T�V��еQ���K*�������,\� �ߜI~�=@\����h�:=?�ʹ�x�z�2� �,e�	#�oa��k�?`�:���N���0�7y�����1���������a	�.���B@�JM���p�jn�d�6���a]F�*+�Х`I�U�n��-4�/Wr�G��uȹ��X����}Пpl�j* � ��0dc�T��o(X�i'&�"L����*ID[��ؚ��� ���x�pӃ�q�り��h
X�m�� $�8�m81/E�"���k�q6�b*�gR�P]�d��?'�&B�/\4��x9�z�pRh�0�2��a��,�$�獋o
��_��ł̛��V!�a���SkoV�)}ʸ�Ja~H=d��Q<��l�D�E�F5�_�A- �Cؿg�L �h=2pF|�eM{i|����
[2�]����/��bYL[��l��/M���u�dH��Z���.7��2��.��3gq���LKU������;X
}��1bR0^4���糺�Pv��[���$���t_q#��CvT�Z�qT\�L�;��������XK#���P˄�T1,/�C�m�#���ߢ�x�$��2��o��,���A4�R�j����k����o����3|�E#�}�lh���/_�$�ן#1Z��XM¼<�z �H"���LڕP<!����v-�z_3o?.�7ʴ���.hx�AO��:(\=��l�y��s��C��7���8����!]i	N��I�p症�7�
�����J���p�p���Arvc��$�*������wvO)�͖]׮��w���GH�L��b�6L�B����|����#)��7�����dtR[�.Za�q���'QS����� OB��I��7{?��D�>�!V"�-�T�
9�5YJw���D������!�s�?\b�����JA��m�<������-���������N,��Q��ф��A�/�t��������!�Q��Ŏ��������%��%F��!P����6_h&���AZ1�z!��c�G���fmi�hy!�tL�t�U>r<��ЋW;�ߙ��r=�-��ȭ�_�����<���غ(ԓݯ�";��l�-��+)��`��*CL�V���I-.y�`�T�^� ��詁mX�n�^��UJ�VO �2�u���	��4w�(�E��ic$�	��G�&�F��T�2.;�巚�VA�Ebq��L5bk����0�{!3Я�L�D m���ZD��d?�����
�J����ǔ;�����9&��\�
�c�	�	�/b��(Z�#�@i�����C7�v���Ԁ.�L�ξh�z�HYu��`�U/�I�]�dm��"�#��v�%Z�mG����2� 8P�Q����~X����:�g��`��4d�Bhו}���ߙv�<Y� ����$��p��>[ј�y�{|_��k��t5YJ�F�yh5X@�5*7}�@HǴx�t�z�������܀��O�[]Ԍ�l��Z�fE�]W���1l�HtS\$U��k[��+���.� ���(����X�W����C��+�b�/Z7ֹ�j��������PT�+�J:����"��8��&Ky����ipp�(�Iz�t�r���+�O�g�grN�54�^�F�k��g�i��罘�_�h�`�`@�H�/�b���Jt=o��(�?4�պ�[��3d��S���0�����`�2��().b�p���DAH+8aK2�Af�9d���AԠ���o�N�w6G�L���.�%}��ژ"�؈���}e�ۨ�Ҧ�����~;��6�^4��u`���i@�j{�z&��	>s���2�S���6Z$�x{b� �Qn�߽s~��5BE�������dc�Y��*�:�`���1ٰ��}qd��r�Ĺ׮�%���x���1��F���uᗊ��c����E�1ü02��O�s���Y<f�0l�eХ�#�\xF��u��<��_�r���H����<�����}�SO���sʏ�=rA�"��Ty�-�v���iɵ=ST����5��V%������t-���t��pRo���$�'�c������Na��i�������\�qy٤�l۠̒qt1��m֛��Z�dT�K�z��OP�~S��@���ʲ��i�x�}Qya�Jué\��:Q'�.�|M�.T�4��1+f<����%�Q�)R��YA4��0_��+�����[,\�^��8$���8���{;+O��s��|���9�|�b��Z���9T����L𪄏���$$5�"=���9:*����k�Q=h9�N7B�&~Qr�iΚ���V�ɱ�Ҳ��)��h�ɤ!�s��b�pX�bw�57���ީý)�ف[�첤��J��^���C�cJ��S�zg,��Y�X�D�:�6Wͤ�<v�Msn�H#� Xn��9×�/��Z�zn��~Ry:�M��?م�E��p�Ds��߭RX H^����y����%�R]��|^oq�Ŀ�F��0O�,�g�tM���ϛ�.m��I@yи��V��mpdU�:]�5wS��8m����
�pd�~.�J�344	�Y]�X�)ʽ	p�����,��1���as�D�,�˟�`�=O��5�O|�~A͎F������dͪО5ί�Oc���K���rA��� [ȵ�߆�D=�;1ܔPW"��;GD���ݚ*�d3��P��K�z��=�� mI�o8��,��+��ٔI�iq3�Zd�+O,�zu�)�
^��8J�x�2e�0���^���ЗD�N�7���	��"�D���#1B��你����C�8F����72Z_����j��sO-u(�EK��ҩ|4?A������-���rͳ�BD�V�WlU�>�@ĺk���a��c��s]{��_R�r�	Zf�ev����A�х��A�糖Z�O�µ�i,���\A�&D�S{8�e.�8Le,ޠ�S���k�`���gK���0K��2�y��G�~M�o6z�R������8���R�eQ��̠⁳�<e�?|��D���,-7I.�#�s��@J>%�x���j�>\��Q�R�v�?|��������<�ץ-W��r��3/�������LH��x8ZF��<'���
�R�ʹ7�
\?�$U��(���ȡRлG�<t�f<�_ҹ�~��-���sQ���$���m��_m
��U�h�m��kgzŠ&-�U��ä�K*@'Cw>�3���&zΆ��b�q�~>���Ǟe]#@��6�L=ed�	cڰ�<]�Q^�	qB���N�'�0F-3q.�T��;3|ZE͚&踂�@�� /	�2��-V�VP9c���w6���y�Y�db��P����!P�����Rl�.�/�/r#f6��("`�^^2#��u�!�g�z�c���Nή�9�Z�Jx��>�F��	N�t�����$����BQZ�X��Y��*� R� 4��/���Ё[9���)���\�l��<��t����[^On?%@w��^N�F@Ъx
������ӯ�StF�+�� mΔ)W	{�8_5�yg=__��?z��o�P�������m>�W���^<�鈽�~�f��Bk�	�Kļ�h��%��<gV�3%�0���ښ���y�QJ-�uWrT��#OVӥ�C-i�M2+C�$�d� ��1�����2�#��P�)�Tj�W1A����������`�#i�a�����:���Nlh�ֳLLs�F��^�X��=2�8�(p-��c�cxJ��KT����C��]�[�|�6��XmmE�YO�Ou�0� �Be�½�u���]��vaw���z�ZG�c���d2���(���@���҈�2R^�i�@'m�7��E����{�F���<~�[7�TX��O��Ȥ^9Pw ��>�?SB�/^��ن���c-�>2�[��sZMWK��x�U� �k*^��M�Z��:��P���2]=�*�jP��S	T�m�`/��0Y���k!.:Ӳm�>7�H�Ҙc����Lĥ�ag��-��J_G��B��	}���'���|5�Fxb��{Ķ@��X�*����_�fI��O��j�6��Z��3��	l��6f�2��x�R�Ø7��U�*��A�Y�ƴ���%�?�0�ud�`���}���r�(?j�����w���0iDM#tŷ~P�a����h_�Kl���=`�4�.��ۯt]�����yCq�		�v�Ǹ��X���՚����.�^W¦�����[WI�z� 䆉��,Fiƾ���0XēHŜ�p��8��D�U(D
��Zւ�.i/�M��e=��������%�2�u����x���ܽ���[e/��cd�%�E��X�7�Q��H�� @  [y/�MJRp��I}�����T�u#��9�sխ��Q�GRk���xT�`0�Q�xi�l .��i�آ��d1��L�Χ+�%)�-H�5!����qx�F.�Hهu�T\\8$UR
�Ք�o�+R���*����B�.֛�=XH��ΛL���� ��G{�Ό5�"41�j��_eS�d�f��ek���	b�~��6�����b_�P��ͣ9>Y�(�_�3D�{��~�<�qg�ͻ6���;�D,=���(��Nk�#�Ű�R��S�-ہ�Ƌ
��V�	w1�Ҙ]Մ�����ym�%��0[Xr��۱F��z*D�r֓���J�L��mV��G��]w���j��3�v��CY�,K�G +�n��7Ϝ����]�W���>���� ٧Ϣ���M/i�)�5���F���&�)��q�?�}��@!бv��k}	,���X�>���Z��:f�(a>���S������#�� ����>Ƶ�=�/�IS�|wo6O�s�B��^���o۳o	k�ݷ��QzĐ��9P���~�k�r��H����2��4���N�}Y��3�3��{�z|��n��\�ն+��z�L��D�`�8EaC�ĲP��������I"Y��Y5bɭ����&�~���@ޣ��n9d�.�̙&?G���v���9d���]�9F��ac�y�f��Zn@�p�������'�x�z�&��!8���b�>Q��$_%�B]�u�é{�#D8�_�\;))ks�0�"1}-�Z����SfX��������س��ژ�9��*8�YU��65�EŖԦ�6#8u��U�[�����/�߶?&����N��:yH�1�x��]��+�Ѓ����K�2�v
?�+u"�"�b�5��?�Q%h./�#���^�]�swx���s�4{��?1�^f'��)[ΪT�{��l5�D����	�a4��j	;�,i-q�����>&�?�R@�`��"2v{�� pGp���V��9YM#�1RF鍉�
�њ�� f�B=y����\���A�⽐��޶��\���9�ΉA�%w���[YH���l��[VאL�Z�u����r��Tz��/�3����y�ܤ��L�c�g�̨� q�r�{��H���쳓o��p2۾pB�v�D����[���&KU�T��x�o����W*��zAyX�筎"H\�i��k�ŉ}�Q��y�x�ܱ|�U�ΩsW >h-BG�W@����e��c�.��'^#[O���2��΄�e.�&B&��,�5#C�����=	S.K���4~�/�K��_���fA�0��9���սI:�5e�No(݅��F=�e\J/#1���c.�ۯ��4��h)������hX)��g�'��`�_mP�B�^ծ�:�	�L(�mѥ_5���/��I�w�pOj<DSQ��+�K[B�`�zajU#`M@��ue�NN���깠,�
}W��6W=2��z���z��6�������n��%�����ݼ7+8����뭕�x��&�]"�!���X��`ZE�
Sd�~���1�#ʐ=E*�S�tC�ޙ����E9��fz��%β2�
��Q�iU��(���t���+A���S�7=�+�k�8�b�.��CB���&¨��
�;�ln�݉&$z�.ށ�Gf��q�\)���!�6��	� U��a��[N5���H�K����F$B�/�?˳e_�M#�O��F�s:K"~�!�f+6x���=�uӌ�Bbn���|n>��=�(>ѱ[�����������[���\� �)6�n*ɿ�V��Z��xP�@��0���N*/#������Ƥb_Q��U����Ҧ��x~!3�А�z�n�7D;6�WR�Bmª�K��t�I#}k��l{ٵ',?�OE���L�Ow�� �Nr����:ٶ�3� 1�lK�c�-�*�J�@6DF=�N?��� ֮�Ms����#r�LȮ�a¾B����x�}�zS������osq�_���e6'�vf��_б�I�6ʭ��(%�K4����J=�Z�+��%K��;n���o҃��c��vb��1QY+�=kD=��2h�|������ 8����sBZ��/K�����A:�p�4��4WN��y�jnW)�4dn��]�ȯv�L���~l�`6�� 䴠�Xb�f�B�1�N�0��z��͐�GDot�I?���+��P�������S�T%�|.�b�-:���t�[�HK7*�������7}�ֲ)Ɉ�:j�Ӊœ���s5�3~����]<ex)Y�Y��{��&�G��J��>��xZQV7axW	<������'2n�&'HK
� ��nC�9���E'�s��^ mf�hqE�n<�ڡO�E
A�p��s�OK����{��x��19�����s�(���.^���n+\�ȗ�d��dąo빌Ü6��Z�p+�?D�4_N
?b�'K���׍u|������z/�dW�>��yܓc�[PAp#�����q��^���W�)�K�*�-DU��b3Gպ���_W�m-�m����(~�k>Ie�0�X[g˝=��4��b���e��~e�ZS���h	O;X)�z����ٱ�fJMn����GG�v�,<���?�%Ĥ8��c�"=��׌�5���Z'��*�)�ו����X��DG�h4}����+ˀe�o2�����4��.�y	Є�\3�!� �xG	=�
�ŕ*�[����zA/ ���~�ؤ� �k{�/9��q��%�D����	O��#���-�����S"j������9���Ɛ	̐��u/D��53[&��n���z���>�j4 �d��t�L�тz������⚾�>� {@� ^\�"�0*.��t��ѵ�V&՗���>"�Ta-ۉd2���'�}�W�����lV������=ÈIm�ETL�N�"HB��	�k�bi;���-r����g���#��k�zVB������֏��_WW�e�-n�3���+�|뾖�S4��cV*O�7@B�ҕ
�L��o���c�-hϭrW�1��3�RgRĮ��3�k�Ր�aѨ����؁*D�k8��-*9��d&,�e��PD�I>o_D��G���|�<۳�`�ާp�' !�BF�|�Ֆ/�&�#B��_���_uX����~B��ϯϬe4C�I�#Y�ˏ�kzd�Ib����o���=�qŜE`�F��4�O:�T�6��%w3m�Q�3vS8G˳�Ø3��Oݛ4$�ۍ8ŋ��ҕ]���ߎ�K���h�'��c`T�  �l�Њ�u�,�Ά�E%~m�� ���������KlA1C|L=�rzy���`�Th���gif]ʉ��-xo�JX��0'U�[6��:���|����-N�}���g}G�^@Ԡ��^~2��:ɐ�3�t]��xu|��:Ѐ;�'%���l�2��X��k'�HL:��eR��Ơ�9R������i�ǖ8���9*��̙�U�>R�,pKB%�ò̘0�R;��.���W�N�3R1��f��$AQ�d�>F�ۧ�&<D�o�'j�`�h��/�N@���P�����8>'\f�Ȱ��#����M�+��n -i\�z+>;F;�$�'C*
�ɐ�xD2�'vv<��A\�����T�豷��B-[5�k��f)���غ��,2A��-����_��N ��b��(�e`	��" �<k�G���cM#��i�a���&1zJ���ʏ�a!�b�E�N�l�z2��`ƬS]��时��+Ҷ�"�_8��V��|	���20}t����^D4��1�=QXN�"�N�gFS�%�j��5�	`�b�����o p��<0���k�K�\>:"���Wn%��.��_��K�(�N�u�wf���-�4W�P�f�/�f��W \Ҹ�����rhr__��w�^�c��%=m�̛�cu��^)"jy{��<�}Cfk60�
vr�������ݡU�0�綔��l�?hsB%�I�3v�}��ʺ��.�:�ih����'ᵪ��9�� �:T�o�d��t��4@ط��$��2��P���ߨ�W��ھX�
$��	5�a�>�M{�'\d�>%P���R���y��[�'_�`1�9"����`sF#j�J�O�(�F�XB�	��$Ϫsf���R%}I���!_���+X~H�"�Qy�
��5�ϰ��I��'�@�%_�wb��E����Ҕ��*b�u �,��T����A��A$�D�����*z��k�Hf��g�~��g�c*;�U��^iEk�$��Q�#4w��v�$2 �[���"ZEq��~@�_�R�A��4��k$����1r
��`�q�U�1��#��7�3]Q���&�5�����u8?����Á�O��R�6�� �2Z�G�����1�;��_��ڄ��v �%����Ȁ��y�eǩ��9�)��&(x[���G�cd���*sPvd�mt[�n�Rr'��AζK.� ō2��Xq����-� �[��G�g]� �~U?�ݜwޯcR�&Y=p@P0�u~䲩5)tx�"��+G Y�>�^���
�����[�(� 7�I�4�\1��%� Ah���9.�;��'4������<�l~9*����҅I=�!�n����9� c�엠u�ĸf�ㅴ3I�nZzL��f|eJ����B�$*s	Ju:��W����ev�t^b��Q���G��B2?˯��6�������f��j$��n0�+��T����� !��~ĒwR9ĳkyf� \�a>aթ��^�n0͸�a-8�ē�a_[�)�{5� Wf���p���yh�X�*��)��/����݀�6 i:���g-i=8�&h�N\T���&�Z�Re���t_��c�������>���DA\-l�~G��OE/J����$r��asfE��xt�s���`���[0!%�㗺�M"���-�P��ԓ���µ�zm|�H��_ܥ�5�������d�ْ�PT"
I��`k�Z�rB��-��nSm.'���
��tV<�.��%��}h��ZN�֫>��hAi����Q��J�����)��������Q��g���%<$���T�gC��	u�Dq�����R&:�
��ڑ_�[��L�$�}d?v��qk�b7�0_r�6%��H%�v��a�j��3S|�T��,��0f�i��ث<.F��U�7�|$:��3�#�V������q�*u�����ho�-/D����Ī{h�s�7#I�o���"?�����
�l)	m�Ky��g��f�V.-h4T!3g$�ܖ�����%���iihB�]����U����ƾ���O|U?u��@�M����K������׶�7�	#��G�\�D]�(�o/�o����TP��9��J�
�^�N��r�{�Y#�E�:���𵆹8�b�0r�1#+�FT��F��SUĲ%�i������oĲ���7ʄX��A=���7��!ܰ�%����q��`���w�������s(���/5k�BHM9��ڭ��7M�|���(x����c���l0��ރ�7Oq���с�%;i�xȡ7L^�nZ(��,N��}�w�
���!���G�k[~�F��D�`�TG�g/��[L���UyH'e�F��ųX}\����b��ąc����|&�w�S�%P�*�P!G'���М�q������KT$U��x�t·�!�Ӣ�t~vG�a�u����.N�o�r	BE�"�¥�����qm�@	Yp!���#/�A3nDt8`��QZ֔����l������e�Ց,���ٝ�)�P��x6V3V�C�A��]�B�(�[J�$6��B����Y`��D�|���)�',w�б�뷉a�X�@хClm-:���G�7y �i�|!F'�w�"�b�����4���Fºa|'+���?ݣ���h���9�@���䎐��T9�' ��z�Iȋx$c%7Փ�/�5�����Ɖ��{�__$�t�Ur��\g����J�Z����"^Õ�����}�{Wc�5�����G�����Ҏ�}τ���',����U1,��'�z]*��Tg�N�	T�B^�o�[�a7��H\Y��K0~�AȢ�jII `���� �&J��i}1,^$\d��N:�T��%�x�w�ڢQbG]pA��o'���$l�o�.�HZ�'q��
wC�ԑ�tF����'�ȣ��� ���k�.!�Ϸ�����5�`�T����s�5(S�P~���/s54_^�Ҋ�7ْ����nX���-8u=%�7Ϊ�y�*�B]�T*"6gK��uU<��u��AF�z�R�������1{)Z�`�-��(רp�è��Y�Ư!-�9D56�>����s{�=�a�|�=
����Rw7�AS�t�)�_���C;��<�F��5b�|�ɴ�u�;�눎.$��+𭍤Pڨ(�$�ɋ�	^"��S��!�����P'��#���V�*+�c�^�?|@�Ӟ���6o��:d;DX6r}w�Ŷ�6�j�/�� ���(��0�mN8�	���5�q-c�^�����$��Z�L9�.v�ݼh�ۓ���4{^�*�T�u$�=oFR�I�����ǰkm⳦@|��q�&>�>q4>uq3yQ���W�<�
���u�=	��̢���5[��4������|Ƞǥ�9���90��x,�]�J!]Af���REK0ڠ�<BH�x��\�93�w�vv�ŕܱ����c������=�����7�wp'���,�5VPe�[�i��|���+������l!b�H���2kT��d�����{^c+�:���a�0ѧ�|*�8렄�?�H#wr�W�:�P��H4aۤ?������8*K$-����&��l@ԻI\~ˡ`��i?�X���ǩV�1�|��f�8���0�qu�#00����e��'Z���<\�$�����O�����0�. �7��
��R+
)�AN��`�T�����"��T;ז�'-�8?{�b}��G����%x#���2C��9��9G	�t����i�G�{f�x)Hi:��+��׀,�ܖɋz��8qA�
��u��޷0��@�bBKʶ4�i���k_�=-�D�e���pZE��-B$4�,�J�k,��Q9�Z�5gp7�Pr^~�:	qz;���}���	{t$�ZI7�l'�ٰ��
��͠��f?7͎p�:����e��o�u�bI��ͫ���=������f�L�zW��Zx��<OYP�{keb�-��ɽ�\���р���K����c�z�YW::}+��E��APg�XB�8w�D͸ş��?ЏL�P;~� �e�4zI%_�'��ە�����MQ��OY�q)k�V0}�bL#?&�7"&]�k����:A�����p���T���^\� nYI��Ƙ?.Z Q��Ё�qߑT_4���r�y�R�8[�����Qǡ<�@����� ��b��7���՚���n����o�}[z�E��ޯ���Ya�N��l��D�q���왨@ڕ����h9c��y)l��*��1�uT6���[���k�,{'�����8PT6t�`㔧�~F0ax���D��]�ʭ|�N��9@����BN:)�e��"+?(��N�-�E�t�����D���?�AX3P7qv��PS�Ď9��0-
]j$�̮���`�ͅ[���]2m�����X�Uf��zX�e��V�����.JSL��ʄ�Af����c*�A���h��bə7�+ T��r1r��B���*x=ӑ�o���\��58�+�.m��p�,J���c���)N;���르�"ւ��|�����څ��pܿ�l�
^�5�	��e�Ⱦ��n�Rt��v�*Q/��,�.��������}��ߨ��ue����
��5�~�׭�3�]^�}�PكU)����~�C���]姎��u�Γ���,�#<����l�>
ZFU���Z�%DQ���Dy(�� �&}w�����\�M�h���t9S6�4�˷"9�3М{6��S��a�c�	��b�;�D	�#���wUx�|��j����D<���o�|^,��a0��,8A��֩�+�P�% ����$&���v�օQ�z�E��p����vT*�O���I�WW��t�	����D]^��w��H���&�r&�.uvn�1��L��K��*�2YV��G��Qv�jX4^�Z`�1�p	�G��������4�1��{�y�Y��d�c UӾ�VB����ރ� �j��OZ�z�w��֓}sH�}Kz��zpO��IŗKYd&f�7V����!���T�؊����*��9IH�7�9�a4���f�V-��aK~ ��:̡GJk6F�ex/����Y���)a@�'�S�̼��}b�)��9�2(7�c���F%��|0��ؙ�&�n$)+�zJ�Jxn���⾟e��dG͉���>1�i�gm�u�g' `���G ߘEPXj�FP���3&{�Y��k��$>��:�����[��R���ё|��U�T~��z��1� 1��t"~��� ���r�@֡� �F�c�*�l�����D�nx]�Hڜ]jRJ[9��K�F�rM�X��G�(���a,�x.*ӊ����B]D��Ҍrfʿy~Kt���g��í&ʷr7����3ȜoB��/��ȩ-���D��7��r]��K.��l�ӹ��k>mu���,J��JG73ƅ2k����ѷ�\��D)���p��X/@ak�ܜ]v}�%NHg4�>�3W�J�D�e� f\�=]֌���_�+w�	�'�uO:�x��$��] �ʅk���~�c���I}]�y�6�z"w�FֱL
��L'YCJ�]�]�����|G5�����fz�_ip4�&���S��Q�:՘���Y��_�u�0A@���Hsy��G�^~��f����.�.1��Z��t������\if���5�MUC��IM�YF�>�
����*h�}u�#夒�/VM��~�zc	ˑ+U1-�K	��}��U�E��C�+����m:-˭pqf��f��೉�}�)_u�݀]���t�%MQq�V� apI<��*�E
٨^�V[%���Ͷ!���d�t���- J�P��n�7�L��9������B�i�Kć$%�re���{h��)���y[�������u���D��S����ni�����Ԟ�Ld�&�p�vzS8T��t�/YC%f�
��J�;$���Igċ��O�@��b�@3fֲ���� K!�V{��Du��t������}�T�mj�]�ے�WY"��W��A��0����>���N�&p�C%����,U1�2��}�9$4�|��2y�ɎUUo����!��B�|�����G�AE`��5L�Z���~�����=w����G�����xǷ�T��\��a�Q�Z�.�ul8��S�R�F\"is@�;"u��-���,b��+���q���qdS�q�$�)A���Dv�#k\�\
�f����9�Ⱥ��6F�EYs�ǧ�s
��:ا�)�
`���r���8�+k�ZI��J�(�� ���yd[;�:_��*���P�/#د�m�����"�o�x�w�6���(6�f=��g��`>QE��b�5�V�q��Eq����H�Ռ��f��`$Q����Y��YY�A(�`V��MG1�?��C��6�tdq�Y�L��7��9�Ҭ����,�Oq5��"�%���Ã=��G���6��iխ��#��=��+�هj��V�#k��d[��z�B��c���/6L-�ghh���K��	����<�aЧ��P�,eS{�ܮ0��W�3$.����d5�m�ԥ&���Ӏ�W���Un{5U%�$��I�es0�E�!�#ԑX0l�>y����_ fCC%+j�8�������_��`i�Q��(:"V��Q����&�S��x�}N�T�hl�i#�ܓ*CDy���s���g��&w�KY�Q���Y���+X4AK>@��SR����?��P�C��]d.ʸ����0�����~ǃ��7��!�S�6���ߎ � ���{�!��4�G 6&N@�� 
�gf%zw$�d3�E���ҩ�b?�d>�\A?���c\ �������bP��Rd!(�e�{#�V��G���H�`j��p��,��`g����`�@��gH����,�sG���	���>'���>i��[���Ń1��Zɓ���qеfl_�����?���6n�B� 6�@LAi� e��|WJ˟���͌��O�"���n0������9-��M<�?�5���Eh܏�����{�^MI�j��I*.^��;Ki]c�� *�BX�P#GB��) OӉ����[)[�i�a�[ݥ�#&��-I���؞��yJ�һT(I%̻~8�m���.�����ݒT�{���g�ϼWB�x�81��*��r��_�Z�����2��jTD�ѭf�%�iX"GSS�xȲ���V�I��7O`꩓Zw݁��	\�
��t���c�Y`��G$��:�]]��nF���Y�`�}μ_������r=ث_\Wߕk�S���t�	P�֞�-�*������n#���g����D�4�����y��Ǖ��8��׽�u�ũc�wJ�\2��ڜ!��J`���W�55�x��H�K�b]�
}A�����|�)�xI�`�W'7�#�ɝlh�ݔD�bT�5F��h}����_=R��M7Bȱ�0i@�>�g�za�*��?(����:E%�E�Z��J`<��V��� 7�]o���[�;�ƞ�9=����/4o�̪x��h'� �tZ�f^� �Z�P�R������mW�]��^��hT`X8t����I��y�� v!�Þ��'e�u8�p�9�?\{D���
K���z���n�`��a�p��-j�)�9/�~/pNY�]>Ew�<��m���6o��� ˘���< 1M��e���w��Y��������9�H9x��F�=�E���6%�${i��P�V?�ӵА�:�](p���w�&��Y�L�ߺkX��W)b[��=uǡ:��,�� ��wU�6n�X�(���b�y���������6To�=�����	QECR�ԗL	�'Q��)�� ��B*���r���[�A�����
i3L���>�hy������*l��ߚ����ȼ�7������Of��u#B�a�X�;��x��y��4Z�4g{�_��P�o��%��A�r���-�e���u�4��Z�]u~ %��:��\�r����"F��C}#���~�@=����z�<��%5"΁��J��;�H�]�S�F]VB<�`��r��	Llz�/�~kaZE��|��H����j�I	쾨�ք�x$4��G�ֻm�B��P^:f����D��=�4��7�"w06��=���{�!�m�Pv�D4�(�:B��͝5r;���;�-ۢ}�5�k{J�P���&���$1��V�S/@���`b�	Œ�mZw�t��᝷���l>w�Q%�y��KH��ۘ������dςh3���q�̗�xz�@�yL%�S�n�$BMd���V�w?�����0�E�D��]��{�OA����I"���	??f��S4e�j��U��No�Ol��h�ra���.G���ܮ���"�YFI?B��i�5^��At�3w�M�L���w�f�;��ro���ih��Lu����9.��{�����H���@�TR�xCo�(/��/}�J�HL�����.G����k�s��<�"��X��j���;W�t�|� ������JAQE �F`L�T�h�]��4�G8+�g��1T�\���#�h�3��$����Ef�U�	�g���з�[��ژ��4��h�U|�r"p2ǹ>�{��4$�L־M�4#?bs����#�tM��D�p�s�o�_�ϑ��[�5�7��8SaQ�S5��{����,t8�Y!J�����9�,�r�ֶ�rɼ9Y.��G�	}R�%�1c3@�~�}U��>^ �5��e���qM9[���)?o�j���q�@4��h ������g���Y��g��L��%�Yꆈk�V�[
}����$I�*R�~=�/��O#>&S�W����)���C89'�Q�(������n��s�4�G�	5�C<���W��;1�����_�1�Ϫ�(ޥC%N֯H�p�`�|��n�xW�J7uT [���[�ue�Є�vy�ӡ+�
�AD��-���ﰭ?�э���^�<�JK-�Z����W�RnhMH��U�,.���!�Y<N�G �OٽK^�8��d��V ��}k�)ӗ�eK����}ı�dwF���F"�ڑ#��
�;9��Q�/<`��{�
�k)���:[�lqg#� ��c'�:_Ф>34ϛ>���j�8
]�ߗLFs3�qjm��M���K�Z��#	�I��>�6��q�pLT &nW0ƫɍ���aH9Ǐg�4���pFf���ͪ��ߢveF|q�=;����*��d���W7ʬ�'U����}%DH�6� "�2�$b��S�����q���`I�;R�c-Tq�vR�e����-ZS�#e�t��a�)ڮ8'0a9�������1�'}��������_k��'�"��@�f|�&a	�Mb��Iq)�K`Yc�K�n�����t�����-�"��("]_`��aMʇ��4WѺiߚ���)�5��A��!� �?Z��Wu��D�z�|J*�$]l��ti�=l�j�?clgP��l+����L�0I�LW�tmB�?��
'�e��ƎV�Ł��ivΤ�c�e��y�nF��r�H+��n���v�a�ʠ�)V��(��� M���4H(��al��F��ק�n�K��R��^�f��:˶��V<!�c5X"�{�-zv�4�T��?A��Hi�p���g�5�e9eغ����3'��c�� -ז�W��Y車!>]�C������q(�ϱ. <��.}/	��|�@��ok��xI�]�t�cn1��֑��S�sqt�u֌�E&ϢLnjT��t���/m��?�d_s�ԄM���UX�QJSי���Ѫ,�9�(F���L�����Ց���*�L��r:�˶}b���u�v;7e%Nd,ضT	־�-dw<�]CӃ6��	?���2�3�&/�)I%��E
/�/�pW>�[�/�����a�,r���R$Gܭ�H��s��y��λ���}+&��6z���_{�$U�x2*����p����(B�Y����;\�	�龯o�F�3?�	.j␂����6v�-��ep����N(Y��ݹpuB�cI�#E�&���ET=��d�U.І��u5J���:�Ej�k�%�Q�F��μ�Ġ�Z�au�y-K�WZ�R�6�Z(�c~�i'��I�ٓKu��1���V�91>��e�(��!����;�:G��2g4Cz�{V�.T)��4VVb���Ũ͞�m�.]+����r������z����H�B��̚��������iEЕ[�����A�\�9<�I�3 �B#a�$�\_O�"0��A��Yɞ�P�C ����D��Kh��s&�u�v�c�ձC@̭�Ïք:��s�.h* �n?��eᗊ*��@O�3�#�i��t?%@�eٻ\�c
���� �F�4�� S�4J��R���
�?hmA�ԍw?�U~�p����
0��MF˞�p�%AR�@�1z��I;�~䠬7}c���fC?�XB�k��&��t����?�.�X)Md��d2�mL���mV�)'p�8ɛ"�Yg_�)� ���-�#�䙩�)4��b�S�f����T�l�ݺ,s�ʀK�|e �Ke�
i�8���}a
���v"x�$�a�V���	���\�3S��= ��C�ϻV��1�j}}o6]xn�y�h�����B�)�\�N�M�>z��<6����P1jD�'�&�^u޺��J3��#ȵ��F�Q�r�`�&3��1���sO]����7�fA�>iH(�3��QT���U�c�01�_I�2ԟ�h)�2��f��A���I�..��ԛ��e�ď�z�J���d�� ٯ<A�M�+�:�*��i�6��x%��泱���RAJ��ِqt���Z��c�Be���g���N�]A�@M���2Qeul��_F��ް���1`��W��CY� @�O	Ϯ��M�%%�o��V#!��n@������}�ќ.P5m�3�@���`JKB�k��734+����h�c���W�M
U�A�����W16�V�ژ/?�1��zB�+�3A3�&�����Щ��j� ֝����Ӽ��{tsM:)�[D����WT�gO�Cw2+ȧ����2وXF`%�lמ6+2�P��)��rM|��^�`��)�8�hxn�9������L;��J��w�8���C>��A����%(�8،��\t�I��_�-
���vUS��}#��<��b��U:_��	���K�\!��v�L���ŗ�~�"c�p鷭���k挨_��*�P洫L��lf�Í�t�{�v6�ĝ�L����eJNG��ӻE���׼�^*�5B�L<h�� T}(8M�
y?����p�k{Pj�[i���*���{��PIF\5>UK�U�0F����eZ��A:��%Î��.�X�]ڛ�}塇p�X�&�M��t�a)��4zaӌ�D�>L�!�����jȆ|���_��P��Du��N�^���Z����]a�Z�lQ[�fs��5�����
hտ�U�m�n��);H�sM�'y��t�Ʀo��!��!�8J�}�����)/9��6�9k�͹t��-�u�I�
[3j�e�k�!TZ�j��l�X�!ac�����;�n��^B}`�x��S��iŸ@+N���3�B�B��\] �-���(�^u�L:��6Mq��9^%�.���o��=��ni,N�3�Ry{森Ӧ9���ą���ЩS�T��7-*������)��8���rxj��W$�-Nӹ:&+2M��M�����\���uFu�7|^�-)�"h��,�auB��vY����>��\�f����N�\�������{���ƞJ��#�n�%;ݝ�{���
K�l729f�x�F8�x�k�n���!|�&��7��GH���n*�à�Z�GB�bX�*n�[\)�� ei��q��E&���J�P���N1�ٓ�U
��W�b�9�~$[�T�����ɰ
��:�_�A��C\���3���i\�5����g�PwX�c���z�Ѡw.^��%m2��Nh̻���Q���
�Xr8�R�/c}|��.�F�$"�p}�"3�|���$���۳	~�Dzt�h5Se�$�7q"��}LI��嘣Ҫ�F�>�xu��M�ę��ɉ��D�K��e�=�VCͧ6Х��"�A+-v���I�����FP��jHHZ"��H������'*���+{Dw�$�ۼI����b�Hx�n�H��]�1� =���K���]��SM)^~��/�FC�pК�OcD�A�a�
��3o�Et�l��n[
/�!Pb\r)�=�v�R�%�g�hO�XX��-���;�8!T���Ab�,���-���!l�  :0�	�9��xR�E�U�d_U&�z�����=��[��j��]����n������&3��6�I�2_0�?OJ���-�Sp��PlȘy�"�])�H��-W��A-PuVru)�&���#$/��U���王��p�|?��P)^���P������6Tߏ�KI��2����DP�*��*b�/��?��H��+�R�fe�_�8P�	�*��h,C���c����v4?�����-��kL�*Y��_�G<kSr�{l>^t��������<��.��Kg�JK�V��� �
o��@Rm?���?��Rx�s��qH�H�'��ݘ~��:�\��A��v0��еRIw9F��N3�����](v��L�><�d$O(rs�	��gPS�]ۣ����D�3�L�r����f�<\�7�J$'�����=�~�懀�l�j�Nϯ���>(�ڛ�݇�1�la�C�:.ϲ	�@�bӗs5�)w����"�dH����`�31��6#1��D��3XmavI3=T�;��=�a�uB�^�7媷���½�>�:�i��V�0��X����_��+�H��e�(0ve$0�NoO��j���vwC9��//���RE�\�ˋO����gp�P��a��@�}Kx=�][nn���x�X��i��)�}�1�`�����
����������^�!h{��!��[�2����{kk?)*�--�
��v;"��<T��,}�U�T�MN�n�t�t��5kJx�/��to�q|�䂦�i�[%�B.��뼤R7��<�]�,@�h�s?
��`�N�T]>"�E�|{Ƿ�G(�pPC:Gg�����(���pD8P[�S�g�ǘ���)�`���FB��_Q�M��Џ�B��&w��q��o�NQ�;�y2;a�aC*�H䏊�)��(|>ܹjv�z�o {'u�H�n�]i���_���7B�OIOO@��i'o�q,0�����RWEn��(�8�*�+3�L.o���7�|h�ݘ��󧦅�X��"��sc�2;�:w��홳J�Ь5�:T(H��e|`�Qft�����z�hC0,x�V�r`�	�D̓�[ޫ��A<H�w{����H��ӧ���L|S4��Q�DN���'�����_H5��4Wo	������#>v>篰ɯ'?��igTp������ s��|h����y�s���	�os�����|��>��'�[�'�ɂ7�Am"N�u�tF���>�EZ
�d����$�KVsp&b�6���$4�&ƌu0p]�̊8��漘JL��{�WTo߯t��Z���D��	������3�P��m��P�h��$T4ߜ ]=�����쨣@�[�����T���7��+��9��Z>���aq�v�s�@�ќG�<�>i��;�Σe�)�]~Ǚ��y�4��_ߕZ��o�1\[}�Eh�� �Ú�%)#:�3j�l _�C������1V٪jCi�ŭ؉��|jT6�F�}xqJ��������W�@Y�&�X�T�P�4oCD��3+[�Fp<��|��W�?��7�}�q����cu^S
����@#SK�I����D�i2���$K��.���9�vu�k"��%�v4��r~���Lڅx��C��+ LO�+�h�
�S�{݁՗Ů�.��#�nj[V3E����*��@���`��§ɸ�E�D�2��Sī��x+�
�p�d.	c�Į�T"#��mrΕ��h�j���O�A[r_��R��=Uy0v���a������������V�X��N�s��Zq�0�L �\�Y&�y��܀�.�9��d3뀑���נVeey}���(.�����~�K}��)�DN�AJ�;BF~�R棆_�n�H结xLi��#M�i/����3U�`��tDmodCR��x���(�"�E��q<��fn��*Ǚ���n>�T�m[Frl�$ˣ��D�_�Mv���S������A���Y��.��n��-)F��OF֙ʶ���؉p��	q#b��Sj5ҵ�����[A�}rC�$�&�XAOҗ��B�j�F[����j%� -ի���5�]G-"���1�Q��֟�m��tЮ�O2��D F���0.���X�sAHD���<���e�_�F��)�����oY�8�]��CszyQ�.]�6����K����o�`, ������ah�dL|��ߴ=J}�.MF�ha%ٕS����F"ѡm̵d�� ٚ?\�h1�1�����|��͜��qae���>�.dS�����JR��k�髜�u�HuE��I���nC�����^z�)U(���[����� ���A�o����j�MDZ�KQ��)L�P]��-����?,T����!ԁ��9z�H�Km9�^A�8)A�E�#�L[�E���S/9����gf��c���PF���F"L��[�(�.�
�rv���ѐ�
���Nz���!�m����^�vA�ܶ���Ty�H) �vB<�PcOG��.�F���[(���g��Ӌ�y������m�5H/!l&'�>�PtU~�9��4+�"!5&ǈ�O�qb��_8�v�`�`�J/`:}�a�m���R�+��je��'�Θ`#��T	����������u�n�7k�9�D�ܱH�}��]h������A@�T^!�o���e�4vw������8��}W���kz��xX���m��l�������)<S��Y4Q'yZ�_"�CwI��z�I�t&�Y�9�$b���6ڭ���WG>���8��tM�`��_�1��U��>�n����&hF�)>\�Ѣ
����zY�+'󸑪F�Y�%�+'Z�~ �V~�{�l�Þ0��G@mD����%��^O�DK���O�d(1:?jS��%�?�>q��1x�}�k��W�z�B�^78Hk�A���ӣd6h���d�v�#vK%���N��f���I�$�I�-H�7�+��Al�mмpGS� g�5k�W;u���_��PR�Q�;��NLȂQ8{)N��r5�����L(��(����S�F��[�`0��r�{K{H�[I�*��}&��O��`E͈7���m�,�<3};M7�*�l�PL��U�-��t��v]��W���jXj�T��1���������p�^��j�O�0�x*ݡ~	)��W�6]j�0�CK��J��S<�a]��JA�V��޲X7�E�������m�;v�\0�u���s�F����I�_�^������m�ʃL�-����M)b� �c qL�0���ҽ����NLH�g*���D������@���D��p9,��DN�����<MQ�^H��!��wao�7y�Qa�;�¤����LNS��@�}E�Ղ�i����,��MŎk@?6N�,��!"/^��c�Ϙڇ%]cuVlG�W�mS��`�0�R�^�?�g(LkǺuRe��	�ӭ�|w�R��b��i1gIsF> ]��l+Hn&�[�W���O�T�5)��\"x�'����i�Q@���i�ŷ4J���螓� 2҆Z���<Қb�hY���Ə��Y�!����n&��&�F�8@�D��lu��n�Z�=��F��>y�Z��|�rf����G�'*k���43�L��D<���~��lM�\���"�^J����&�� �+����|��}�Xv��!+�;u9����6b9�o�-�$���#hG0�����Zp[�ɏ�3��nW�K2[K|��q�8�g}��Ռ
'��~���!�J�l2��%��٤ZV(m7�N��V�,D�(�|a|��%z��h�ǘ�nCWoW�*{c��\ذ 99�'����?Б=^�1��jbu�ߴL��l����&�S�wMz�� �ļ;)����x^S��.�qg�W�$��R�d*��LL2����^: <Wqq~�`!��t+"�O��p=WL�l\�b6����6KǊK�VL��ۗ�"�'+3�Ȁ�L|��~gc$���d=��ߩ8�B1�sK�><�n�����'���&��i3��!b9��b�6�v��*����풜���\�l)��NָUf�3�f�P=����h C׹:I�����W�7uM�a[���%��*�y��Bc�i�Hj�V��}u�Cݵ�B�\�7w��SI`�y%������A#ɐ��ݹ�#R�X�*���&RuhH	ho�h��V�0��Y[/g�#2Ȯ1&��m�u	Ϩ�����|4�� f��u{��4|��B��u'�3�ef��4E1��2�i���N���Pn�� ��H��C���j��4τ�u��й�����gT�otO��|~V%\7��P�:�b�$b.G�7�S��r���Z��0&Ӈ�Q�?�yu20�ӛ�:@|4��.�b�όa���;���@���4\�[�rf��2"m�p�S�"�B��C[Mч�L �̭�MRC��\V�\E� ���:4߉˜to�ڹ�ٷ��ap��7��(�����F�j?�V��+&��}��������l�>�����~lO?d�$���r���j�z���k���7]�n��f(�鏘$P�e�/�R�c�Z�O֝Ë%�"4��_�@��3��a*#�ѝe������Hҕu����T,��{���a�ڲl�p �7LC��� ��`Q���)ʓ�p4.� �d&�+1Z`]j�.�=c���c��І��ǩ�ls�.ׁ��^�l�