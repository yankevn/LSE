��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��� ���/M��ƨ��s�K�Lq�"4=z�ѷJ���VYO�i�jhKM�/�j�z��O��S u*��o�1k��������W��;��T��r���Ylxu1�'�׆FzX�qgx89*}��#������L�ܽ�Fg$G���������"����k���� }2�?󍶔��3+a���@�_�4s���,���l��v�C�.f���d0��%�C�Wv�l�{�n���J��������b��r7��kZPP�$��т��z����{��N,�2�HF'�`�_h�S�y��/#;"F� ql�: ��c��t`�e�2d�oPQ^�и��;4��y��x�Z.�뿢�w2М����z�#7_ٷF�����Vx�R�h]S:��c�3M���zW̸�T��5�Ճ��Azs��ߤ3-� i��F�f�R�+m�j3&C�W����
�\xd�kf�s�H�nub0uUO4�h��u�7-c򠕗%�R-O2<�ק������\놧�oD�΅QT�W����_]q�&C���d����=�Y�[�������]�%�7 w���I���J��yi�|s����qX�M�G��3�ģ���q�p�#E	F�P�|GG衍�E� >��(���)R( G���&>V��������=�!NH�(d��/Ĵc�@�h��K�5B1��`	^�0a���Hܰ�$
�6�P3ĪH���!�s���6W��b:q���j<��0�*4~�"{.�Y��aGn�.j`_ �M1[.ȏ�U�x
	z�X��)$����g(s�Bu�Hw����]�81�8��q�V;M��2�Y%@��jH�
&��!" �0]��U��)��QR�9�6�9*ub�_k�P������ST��_��*��9����Y�]$ll�l&=#?6*�`�$��.NZ�!5�I�썌��ݑ�68���G2_*�ӽ����jci�o�[7�8[.<����>k&��lRcX�.|�O~m}�3
���w�V��Lh��`2�����Ѐ�RxTM�jV%\��8��y�Ҁ)��oީ���i&�Dk�q찀�W4{��iGuŠ����wi���Fޠ��#k���Jg�`��wN3=k&�����	�QWt�. x`��X��,S�E�}'�JG��lG�0!A�0P�,8꧌6���\TD�W��*n�g�����`/�[�
i6l����(�������,D��w�e6��qŰ�S���O�.FШ8�4^�SI�xD��{ƽ�
�&��֔}7�5i?>��uo��a�B};��Aѷ=dP9�y��EIqo�<CZG�>M\#�:`���^�h����C�X�CVV�T8��X����:)��ʆcH��L`����"k݁f³�L(2q�f�w���<����5Z{ yvB�	V�T��5�ª@�6�p�4L�s�%�9����QS��'��<a�k5���R�z��>���J+�i��~��d���U��F�������	J�e�g�m�s*a���6k�ݼ�hr #n��Yh�:�A�	2��|Y���*�B�ªК��y����1�|{@ɤ[��T����76;�C(�F7I��I�%^C�~w�?`�zj�N�/ǆ�7�6K5���S���?5��BL�O��& .�%~:%���K^�RE��(F jz=#?Ea���s���"�k�d6~ ���ٴbm��
O�7�u����TH��pp<���?MS�v�^aC��Zg���&_�����3U�s��6�b?����Q�xhȩr�}�<�팻rk�Bωմ�z|U���)W�Pq��#�C7�5R����xN�g����*ڪ���em^:��$��0g�^�J!@�H��3����s?�IU����m�ĕ�2���R���D;evs�@��fPu�}rI���Yc,ٻY�����W<T�g�9��r����Ɔ�`S��?A�y������W�?��ۼ��u��v�|�5#��#߭��n6�Cn���HɈp����zP	.���0�G�����Ť-�z�g�����w�oέ�B'�:_���I..K�	�\�t�>e�?�van�eu�i}�����W!�k��Rq�k��d����g�KJ��3�g�ӝ&�W����.���
c�/��r�(::	��,�L��\X�\�@�g��픰��O�\9�rC�@�j�u��@��~$s\3�U x���Ɵ��L#�;�6�H�OP�qcK�}{��
!����V�˱�A�Y
�{Ǖ�J�r��hxl���)��u�K�h���W�7 �'���Xr���T"E� ��� &��(
Ӈ��=��rP�1s鴒�u�h�	2>]d8��*p�,��bf�d+�&u+�����=V-2sp�|�C���f���ة��*E��Y98���:�d
4f������f�0��2�$R��}� ��M9vBH�|	��%N�T6:qP��a`TLCQI�m��^����+5����c�o�(No��׻�87:���XO������Pټ��Z<�,�v��G�v�^�����o{��;��]E��
p�Gl����+�������+���R_��."XB�ȍ���8󏹼�w���BP+�Eh���.�sqA0���o^��ЊE]w�Zh�մ%���iZ��p���9�r��g��1��ʧ!9���yK>\h�<ow�������.%ُ�� S�)k�/<���� x�F�*;��Zp��:���*��FP�>�"[|��eY�r>��<�`\���� #h6g��o�Y����u������˩�b�N��!۳�.�H<�js�;
~'~W\���=I6!y�~t���V��ѻ�l,�j@���[{@�YBc�D���������މ�L��/z#�9Lf�]`���wb����s�q#w_�];�S�⮌h��"b���g�2<_(]�� �ϊ¢�^Ƅ�/��mFi�04�({�֦�j��9)i���`8�~���~�L������y/Ja��'��ڼ]_�|�uL)��J{�HpU�a(���=m��F����&ܯL���>�;6���C�B��o{��wu4̐2�v*K���"��	�^�L�B~�>�m���K�c�:�b��JU9}�(z"<�b�����S�[�Q�+�Y.w�#�g~쥐z��/��5-�|����U1��U��hEYSN��K�V���f[�X����7�5�����B�������8�E�����֞�H�ʴ��*7-�jwG�w��Us^%+Fk*'Qz�e�p�9��x��|��x�np�U󍨉:�7<(�9����?P�O��M�j��{���p����uz��k_	�������Q��9���}
��C��Sѽ_�b��g-v�)j!��I�`~�ʙ6��ZK�l-�)�A�K��(p�x=�"�"��ȅ�vB%Ġ���B�e���ދ�j�h��X�ߙ/�L�+�5u���>*�O��x2,�\ȗ�]�A��n�]t�ؐC�_����P�_�!��i�=6Q�^�ꊃ��mu�'7��&o옝�R�����C��A^�t���5���漆�Y\Kf ��:;�M}:�tgl�|,d+��b�?.��p�ƥ>H�i]��O���������	�Ip�~�/�3�ڱ9�����i�7#�Y�o��7��߯������k�c��Vܨ����~��'�rC��Vb"��Y8�l�����sq��ڢVDʱ��{���I~�DѴ�ԛ� �|e��G��Ȅ.ji\@t�W ��9ny�ۋ���6�522ivX�\k���C�ۜ����r��.�': >��a6���6\����%���}�)MCf���Q�oC���\Y�����e��o���"l&GjW�&<��nl?6+�I��n8�r�X��[q>�ʷ3?*�2J��ly_�3���db�"Pl�n�PƉ�q�<����T (N�vV"�>�ԕ���9��ZK��a�{�qX�탟�J[��Ǳv�l�k�R���؉Dvo�/�˪���9G~�!$��m�V#Rc��j��,�n��Z$7J���Y������
ꪐ�*�J�۱��߅&�(J�X���p ʧ6�1A�l�D�QI�_����o�>�ۚw�yvWD���C�ʵ�xq��A5�u�Y.���)�If�`���]�9�ty6m­}�������yxIKgE�U{P��_��<�q%���bt�k�ʘ#{�Pr��ۄ����-v��崿����s�m|#�
�.Ȭ�3	V��X5�0��o�~\�.�G�T��
�U��D�z2O244�������4�lY��Y��`�=<)�.�%���zW�>Ѣ:(���zW�UT��ɴ6����d�,sӊ~�5mo���7��	Oyf����^F��>�ܜy[l��:\��QeT�
6����0��7���E��Sk��[�{)z�"��L�n)�=W�'a=���cef�m(�]�)Y=�P�\D*f���w��v(>^k�`PdD��}�,�.i��y_�#�@��݄�Y�|�}
E��{3�֏H�jQGU_�Ǟ�m���F�2z� �I�|�U�/3��z%��E$ʱzo�Hd�d��O[��Uo�oي�Zr�X�,$�xO1�ۮ��Y�hR���8��m��^��G�_u� �ȭ�n?L3�w>�<ͷ����sn���W�؎h�����l8�6�#ݜ�+���ǹ�E��B��%s�
\qT'zMo���eX.���BU�bR_)��?������<V4嵆�Gm2����ٹ�Fқ���?�b;��҇��үD���{0 ��wD.��!b ��$�jlu ��tN$)�?*��Xr�W{CF�&���> ����ep�ʑ�[4��II�{�I,T�Jd�D���8&��⸡���PMS[��j�����:����ylѭ,|.e=��`)al���dw�UxiN����Ƿ	ɛ����L��>��}V��)��5-��$f@�[����������"�@�o���nWlWĘ�.#�L�e��1���i�,� H�ތ�E�B$�Kw!��'Eo��� �}�7Y��/I���a.Z6x8�ՒC���q$ӱ��6 ��Y)(�0r�f��aq�A��9�?�/f/��V�!�x��cI�Q�L�E�z͟�k"�J����w������B��ng�d�i���z�(����Ez�#�+ǐ��so�$���^i�tJ@�DM-`<x������o$/+A�ָ��$�u?�%F����t����}`��iE_�8��:�6���cyay�Ĉz��ϙ�l̂��=p�r��U�y�̹.�{����~�?)���Ɵ�]3��Ǹ�?t��x޻oNH,��/��+�E$z��A:8�Ɖ�-��\MKH���R���O��)*�'�G��*��iq~�F���!t�#Y�V�o	,#֚c멛�}�U��C ��&ÚVV�� �.�tQ-.����-����zXr�Ah0�w����谑c�h�]N�q�*`�|�lۈ�@�ӗ��2���ȣj
�qI}乫,�\�Ƶ�]���Ny����U�D��a�C��*@�y8\Do��3����Nd�Ԧd��F��<|4��1��֚�^.�*�%1r�e����`�=�է����F�Ҫ@��^g[���흕d���:�=�����rN�����*�½�H��i�rC���)0�A���ouh	�|:�=��#(�������S|�	@h�o�E�9���:���<��R|[az�K��j��ɱ�ܱ�=���kW>�Tз�A)=ӊ.Y�^a��n����wН�� �6�ߖs�B@jO7��M��zx����3v��wnڕv��L=Vht�M��U��h���qH�sL:^M�6s��zs#�<��:^rE1�M��K"�{��C��[Ŧ�� /Fwd�~�R�#?���\���˸S�r���;fM�7P�r�.�����6�j�{O9lY^�ƽ�/��V�n�Sk c3�����HcOY:F ������}��x�;��<�G^ﮜ� `�ۼ�H��'o�<���H�}:��qV�ڿ�%�����'���?Fv���e@* b�|�K��91��~'�cd��C�>i�Q�`8y]] 6#�,q��L�˚c9\u��Բi�����8��A��yi�!t�B�{:H��
6�|��5ĸ/�<����g�H�EA�(׊Q}MM�+Dd.������ �Q�Pi�6��H*����Y�%&��9�5+*���3�͘w<��=�b���9�M�h����^J5>6|��n��jԻ7��fc,2�r�aΆ��,(9X�o����*�6�Jqȿ3<*�f���(�=�s��iGr��""4v�o�lk�4ʠ�,���H.�������~~�P���`<t;�f���h�`�8M@[�3��?)#ƃ��;#R(���+���}eG�6h��PRAۡ�b��z<�Y��-��&A���xd�;��ub{T����xeN�B�^�v��i���i��_�ta0:����eb3E��M\���� [Sq�ݮ�߾�$EXV�YA�`]R�aNF�S�B��-�O�b\��_�����X(ط��y��W�����E$�N{1&s��OڒF%�b�A�ܾ��{e�z��
�J똖���~o��ȏ��:� 0D	�V����t���Iا���/N�{Qr�hI�QW.b|�T�۬�){XX7eg��[�^
nonze柂��z^0�BH+l��>=��D��iu��Oi�ֲG� pWZ��U��Ai*�����"���\KhQH����h�����pۘ'Ł��˖��U�8����.~PQ���*~q��A�2j��1􏤠T��b�C��~%Ķ�eyctlx�������R��Ѿ?0$�?	gb�Z9��P�+��und`3��<�)����y;���v�0��k�!���!�/vT_K�J���6P|}�jH�֓|n�@��71׌x�'�W��Q�Ov�I�~���ѡ0�+�Wn�_�襩o��%l���]
���%�>�ֳ:<m�v�=U�v!�9�٘�<���a$�jo�Jqpϳ�S�<��-�'�TW��P�U�_v�~�zT��f�:(��u�|z��ހPZ���9\ �C� y�x�,�*1�<R�_)��1�-��7�_6kz� ����r9VI��Ɂ�A�A,�E*�(Ɣ��}TKh�͏��D%ޜ�Tj�Y���e~���%�w���'�%����s+� ��[�"�my4Jk���ぺ���i���dm(뇐+����#�8[�4ˋ127!;�� HW�L�IE3���Wft�5l=��#�Y���~�	�TIO�}n+Vo�ք��,�$�'��ITJ�$c����OY�D����"�=f����َ�s�]�O�P��^lPʘ�6y����L��`8#���ۖ2z�,oz�&ܨ���[��ȟ��I��2!��{ľ�4	�˺��IRg�4��c�F�Y�E[JQed�����Ή�p��	o���ؾ�C��\.4��S	���afX��1V��G������*�)1�C�gm�°x�aQ����`��@�ġ<1A�ȚB��HMYE�z�*��VY���NVW�� �Z{�(D�so�/*HkcHC필�F3X��:� P��Z��o�-6K����@n�d��<�]B���� �����A�n�)�3�� ^5>���s1�Vj# �}]gO�%�+�>�i�i�<X8K������퐇�hSRh=���&�%��ۑ,�[��8~�G#��8职�q\*��]�jp�^��`c�����nE�H��������q5dG_R�o�@%#���𽽝X;׫����I����D�t�ވ(�5b�Gp���Е7��f%(M�Ց�@�%Rr-�t�Ҥ�)��ݰ�d�U,����h�̳�\��;%�UZ��[6Ǭ�[��5�����{e�s�R⨶I�h=����6�o=%����pn[��*c^mB�,�F����M��2t��>AhHt˰�S�6á��?�O������bq�_�l�m�iT�9a�*P���9�z�r'����e����f��2놩�aRJ?f~�:۝��q�u �w�����抑�x��[8����io9�=~�դ�K��>{���������g�p/�k[��h/��x1i{�H0�Ⲽ?)g7YnYmW�\���N�r4�2�㝭�$G��rFv<���T�ujV. ���ޞ��:�����x&�!�Pb���褃+�K��ݲ��x�%����W���`
[6�	)���0�:��r�_���4H2{� ռ��Չ���^�r���L*����产���d�mA�h��݊��W����K�n|�|��>��n��w~]�3H���t�Ĭ9oE�vG.���4C�݂�,�1���Wь��jF�yu��ŀ�@h_H_���t�[�܎ڡ��3�E�Q\M2ȆfH,R:~���^�7�%/��n���&��r��P��m/^� <��Tl`�w�#�'��$�ι[��c��D��Xۅ���Bv�ً��m�0j��E����b�$
�`��E,�#G�PL����Q{����!TYNB�u�/ �Hn�����)���Ϟ�H9���a�H|��;�������f�3�W�P
_M�?�l�������|��>��^��pR��-m�/��pT��`�"�ҁ�jo�jx��vN��-e��%�$z���N:AJ�j}�n@���쌉����-�~�ߒ¤<�"F2�����0k�̞%ƌ@��"r����Q`'H�B���[��s���r/R&�Za�B�%�_�,+)E���b���B������9ԕX	RvR �}3��-!��o�`�Y��/oqn��l>=�h�:z�w1�H\�Z@/��I@x��<�[�Yǅ x�_K*!�H�7F�nS��w�J3���L]���6x��K�����J��l� w�XeoA�(?���u��p�N�`�i��熔&T�d���+-u�mo�bԈ�K�APFu��k�0�ʖ������Xu�P,�\�`�as�^�ό�t3��Pw~�����d	�AGA���4	�� ��[��a�U�<�<o�<6��O��Ixi�T��á�k,�d⨵�D�x!Rw�9]̵�S�e�9�Yh�6�6J2 ���Ι��V*`V�[���2���{�:y��v��P�fNB�ˁ���T�+�H$f^:���k�U)V��,Ǆ���>m��L{t�Ɋ�4?]'�OGto�<��] ���9s}6(U���]a?�C��j`&4-ҩ�3��m�U��L����rL�'��)��.�5�t Ch�����A޳S�' ��oVݱB$��	f�]�?���E����X�>���R_KZ	��O(�x�&��?�mpB׵Z�0.L�:���ObX�RW,�L��i{�)���Y�����'-�~jc2h�!SmL�
�)�T�3�F�E`,ꯒ�u�����=��Y-��%�c�1쪿���Z�<�A%�܆h����Z���m oI�+� �ԻU�d]��eس�i�Xˁ��a���9`Eߤ���q,Xe�2��Jɏ����[��=`<�'.l�]Ě{��e�`9^X���/�|�R�Z�##�M<�$�x��dz�E��Q��@Pue@;P���k1���ͺh�1v��{���s�!��r9$����'�f�(ns�\TzBY���׃��3�{Jb�����MF����e��\��R���c)f?؟���ʔ�[F��L���buGC$�Q&2hm4i�|&!?hu:��.�w���Qj�+�5�$�-@��A>�������|#=|��z�3�7|��-U˨����F�{U��\��>���M��ɡf�he�~��:��T��f���ͱg=�Jԭ9h�h7O/) �{��a�`�T,P�\^�Ht�r��������0K��Q���e<>C�ffR
cp{LӻK���ph�k8� K����e�+�Q�iv���ܣ��j2˿E�a]&�®�T�o(�m+A,������G���,�랾8�o��݀��j[ ����s�������C�Ds�%�ډs��55�h������_���-�oW6ͰX��7p�����{7��T � �=�7YAō$Ad��� M�{������0w�)V��{ ]���C&�k�ۉ QFY�v5���-�aF��W�Y?|��Gs��W�Q�^P[7Ձ�Xk}��.Qh�S>2Y�) .��G
>�J[8�X8���:%ClQDȄ�x���[2���~]�`L��T"�����ԟ��To�T:�[Sݦ���̠,��c��\?.]�O-1:�bIhmo�D��t�l�c�ty{����g��>���u����(R\z��U��w��0�!"�+=Ǳ�ε,���,���������+2�����t��2��?U����*�=���������*uԓȌ������ҡ方��P�	3t�q���U|"�[fl�\��[3@c�l�N_J��,���!sWyPuƀ=��[��&Պ�r��PG�	5�v��bo�Ҧ\k߯>��$��Yܪxq��nd��},����37f/�ܒ�XB�(t�;�_�g52��*DT��Lэ�-���Q'���NNH���р�'�Bĩ�&���׳i�%���z�<ȏ����k�������c�\�����Ca��ɮ_ ���tK!�U��)�)o��e�k���n���B��1BMmyz˄��,�BS��0�R���O���z s���;��m ��b}@��	�j�F�	"i��u��;X;����HmQ�-#J�0Ӄh5�i*: �aj�����v�y f9�\�=kW޹�6ʱ�o�]�E[&���)#c�5�j鍚�!p"��l��C؛��"�����I#��/9�Pl��y]2^�1�!��E��Ii��Fw����.eE/�D���\�+E�`ڲI=YS42R8K������^II�U��lR�oU�f�����ov�����;���uL%���h��>�͸j���|v#��;W�3�������M���c+\`wC 9����A������mE��(��L�\���F��e�t�mJ�����q���&����q�K�hYJ� ��O��w�Z��f����n��1Z���*���q�b�F����þ ��g� �N���D��x]�E9tu��8��2����E��R�Lr����r��@����x����g4��űƂ*!~��7U��N����+�B���r����F��*�2��I(�I�Y����7��
[[���i�M��E��ٜ>��-�*-�.��[p�'0c�j�-_����YB�K�O�%9��S�d8�9%'-�ÿ�э:DL�N}H�z�S��Ĳ�参���M'Q%$���@�� ͈)3�[�� �͡�I���9�HN��Z�b���>����'���Du�@v�!�+��x{d�5�R�n�)W�>s��B�9�5��
��xi�'go.���:"	Z����~�!<��%���/��P?r5q��"��;_"�t]���C��_ķ��������V�-K�{�!��˴ST��Qm��#�[sM%��q�"ѻ$lL�EFԴHL�S�>^Bͷ4P� X�e�au 5��}�l6�%�r�������WB��!��U:�!��"bj�N1���M��5�&�[\{�^_,�J�"%�l�ÔT����Q2�$1�=�M`C�ΧOMqԾ�����=��x��߿�d�&����Y�w ke�h�J�_��R��ɚ�c.-�d���+w�~"�#ؽ��̠/x��fcy&�n�P��,�[���Gn�z�*�lKl+.�1P)d]��sR8�1�>�b��1�L�z`x��-�m-���0l�({��03�KA�1ќ�`�,����Onw3O�����<�Y?�s�@se�ӍC�j��/�qz��;��A���_����:�q��,p���Z���h׃��+6��i�ydF�p@�8�?��Cݽ��-nNR�I�݃�ɡUE�e��=f��:���GҡV�M�{�l�&.V��Q'#����c�.c���\�ZZ�a���&��p8b��|���6�24c@Ʃ���Ё�h��d%�^���t�=�ن�]����m3uo6��i�ʮ�&��C[.�!�!_�@B��@E8d%���g�-�����P�\�5¾*+����=Z�l�sl:Q���+�.�tfY��Ǝp���|�7#@(*�X��g�s�n�g���l�v<FO9��˖C�
w�A�V��u������Sv����i{bA��}���Q廒��uC�"+R~�妒l��&���f�M�P��6Si�K��g��(�83�=�;�FP�o=��\�t���<�s�HD�!���_~,*~�ٴfS0�6�%���O�Y�۵l��K�<� ��ր+��9OX�����//"Ϩ$�&�1j*�,u�ӗH���T�{}�)����gNe炞)�ԃ�>jo�iz��w��� �:�!0�9����[bxӊ��}�?7���)�t�Z���/�:�O���m^մ�$�oV�cM�ܕ�/w�c��j����;9�x�U��bщ(��m'���ۥ��`]��8�K���	^�����O��>C�3�]�;��E8���
�X޴�ƞyR`JY��6�Xa���Dq>��"!�q\U�ե���3�v#������G&��?T%V~N�Mvg�WNi��J�*�QL�sD��Z69L���zF��h�>�U:�R"u <���}�rA�ko挃��7����#�;� N�����]��9���������B��#��v��ӎ�a��@���¥��޾"�j[�����s��q/������3+v�F'��~f�
��Z�OY���_՝���sc�T#�	��IF0��Sj���sf��N�!�G�]m��`%Lm^GOB����G]\�c���=K�N�۰�w �=P&^瀦7��*Ƚ�,i�~o�^��5�'�O����L��j~ *���G\����r��E�Q.��_)�K�iBB	W��K���ͧ��Ak'i���YuS����AS5�!�s?��tgJ!�P��˵y�d�gm����L�x�P����ő�Cbg��8�Ŀ
���T:�0s�Pq��p'�uʏ�f.1��Q�洘D�QV|xu�|vj�߉x�x�����l�x=�yP��9l+�d�Q�K�F轸��V'�{�ֺu����,N����Ʒ1.9� �ހ�v�)[E�^ 
�ATŲ�v�je������6���`50��J�X�Hl�OJ�k�A��X��τ�3�¿�[@�WvjO�YK����W��z�G��Ko�����iT���^@��b��w��.D@�ʱ��[r�h����`�ζU^;���(���*���ߗA�(�im�n.�*Qɾ@�,�����6y��z��[���D��B�l�x0�|%�ለuv��yJ����R6;�)Zzj�H5���(�"�o�B��}�`Y�Oڍ�BƜ��J�A�;�.+�!���f�Y?�Ș�~�R�w����C�B �D��E?��J��7�Gp�����:&��W�k0��į��O@���p��st	��S��o4P�HyWCV;��0�L&�8!;g��:1���$4�R1��'˓�#���n��>i�1��}vo��ٿ�с�fq`z�7����3w,!������w0���k�3�֠X� ����(}P�²�9�П̓�?�Jkt���S2:�ߤE6!� t���k���>&�|��e�9���52;�]��Y������>�H�ߜ��:��o͟�5�^��,Tw��q¥y���X�m&�%
�0}��u�*�������e2���f�E"TM�j� �0?��_�TǷ��~ � ���EX
�ta�nh����ǡ��y�$[e��Nz���1I�X��ɞ�X�0����if�3&R̞�k~���������*j1��$�apH� ��� �|��&/c.�L;m�5kA���ק��P�Tz���{�����#Ff��,��:_@q��I����=�8i< McMnR�J��TC��f���ސ��߲&�%T/�����Z�AE1;U��@R��
���m��pzg�݈��斆$w!��.zk�f�qw���&K L���A����Q��p�b�vUcǲs�u�E���eO|'��� yoM���?I����I���h7�y�(p�#J:�f��uS�]ͳ�ߐ�%�ʧ�;��FȜ2�h�q(��i�drH����;�3�n\���ٺ����SӮ�>V����C��-�S<z����À�ܴЬ~�Jh�׵~�L���rK+һ��şBUx\��lG��34W��q�B�oA�A�����ޕ�g�R�I��'��:!�_^�ƀf��$.xAh!2�$^�Qp�ѡ6=-�b��0�N�Rى��O�#���P�vq�P6yF�J%3����:k�G���I{����5���*���W�v C�E�!�?i��mK���,LQ���ek��ѓ��y�_��v&������-H.I��u9��2t0�QI���y��B�{��4�2�s`jxIW��â����0��I1r �!j)��3y@��Y�2m���:|���F���+l��'�ڛH=&)=T�!{�Qg�q���\�����6k+������z\śO/Q�62���L.~7���~l0��Q��J��f��������!�ӀZ^�,O1>�e��F�������F@	����yO64.�=Ir�p�7m�O���{����oO�C�����:$�+ۼ��F��� �E���F�uCp�� �Ԟ�*츱4�p4�&*-��?.�Ds�a�ڡyP�Fc"���ߚc�T�}l�g�!�Bcc�?M�`־5�n̊C삸>��	���w#�{� 4�6e����<�x��D��?��L3e
~�{<#A�Q��_ ����m�6K\ F������̼�Z ��.��w����Tˤ��~Re���>��}�&�e�2�	f`�&Ogr���w*:�H���74�f�>XH4���&���^h�$V9)�Q
!\�
5��I?�?���5w�5�����q�p�^���zҗ-���0�g���V�hrK ��Wv������ǉ{�1�q,b�Ց3M�)u����h#'�N�f����E��8yv2Z$����Faw�T,��B���n�`!������h�lT����x��ؔX�>͎]�Ou� H�H���9Y�{�2�;l�p_n
~H@��~����V�:�f"Dn��D&v��p���v��O`F"�{�w�x_D	�E?�a�Q1I"�0�=ӰU�m!�]Ct��g���b��މI�_��\T.U�Bh���+T�f�o�&��3�?Q�:�$�r��*���i��>���.O�D¡�»5 �N}C�E/p�� �(���%�sl{n� ���[' &��q��>BO��������pǷ]����&?.���N�`��'�Z�O�ɷ B\�c&]�Г�8a2$�`�ԾczҢ�@��c$TN_mL�G����1Ya��V���ş`��5֫�ζ��r
�X�} �<c3$u��{&���fd)�ϫU��`Z�O��*VR��ph���e�:3�"��ze��ۘ�x���N%��7xx5u+~���@;{��P������e��Wǝ�N��u-��6<S��檍`vz�X�����i��ٴ�ʆ�u�v��
�rc?aN���;��B ����ؑͪ��C|?C�.�"�<W`��Š��bd���
�σ�*���㯈���#7O��A��%g��{���m��s�`�ݥ]�7��QJ��6i����:�n�_��%������n��y�tRR�x[Xb�"�]���k2�N�v	���uci����
>;	��6���~�:5���*�r6c�x:�!2=O�����	�,̢"���6����$�����f��"� 
}v�	J��W,���T�v�����)ܿv�L0��fHZ���JJ���7l��X��v�s����ZR]<�H9!�iU[�&z��ܙ�Q%z�\���RV�A�Q�ǚ�����n�ZA8�E�\=~?��0��)V�/��f���k?��+Oq��~V�M5�L�I��o5�3��j�����ꇬ��
,4���?c�T��G��S4�S$���:45����s�⸣����O4�4:~�iA�P��[�0��	�	J�`��1��5.Қ��3ɽ�`)Hy�ʤ�ރj��R�i0��Ժ.5J�t���Z�"� _�#')�te���қ�$���I���C�~�a��c���J#���y�[��M�����7ݘE��(>��T.�'��� �_���4��lٍ.P� Wh7�(��b��l�����.�,z���ýѽm�s����؊7�p��Z��8V/_O
��o�  �puWD��QT>Y��ZlU�Z8�O_[{.�oݗ*�(��߸��[t�L`�D�x��gc��̍;b�j��b鄃� �JӢ��e��<�.��g���v_��Ald\=�V{�2S��� �^M����]Q<g��&0:~�`̰��B}~�nm�>tICy<�8���1�c"��T��î_�Ђu$�þ"�'�Xvc��G�6�\e�KTk��گ��.�������*�h����W�o`��=8��6f���3��j�?讅MU=P't�t
o� UU�vx��l�����Z�U~{�c'!�i|�/vj��9B�{yet�~���w�E,������j��m9��!�g�}ֆisFP�i�q��M�~�Ҭ���m�g��o�����t���q�������<˅�=�P�n������ٚ�3��M*����mb����vI���J7�P"�)�Zح�^|f�<	fEA�/�T�֏�ڧt/嵀����!�\h���7xS�k����J��N�_S�C�3�%�%0n8s^��n�D�Xo�DL�>���JM�-�!Q�Y�&ː.ڳ���c���oÍe	5�7m|����d�\�f-��2b~d��Nȍ?*�D��ډڊ��k�c6�B']�|
�ӴkKBRP�~�O�B˯��g�y����EW�0\@�LZK!ٵ�P��o����+%���)��X��B�ձ'N��,�u����Hq%�*�G�@�~(��jf��C�,����8D�+ic�E���t��:��=�ElE�����
�Rv�-8FFT������-Z����0=��Qmy���9�	�6[㨊�� +E��)�^�Gt�R�j�܆@^�;P��e;�r󂝈W�d�?vӮ�37�=m���%���9����dVJm�ZM���� ��_p�6z|P{����?K(ش	�~|�"�A?<��������Tu�8�^�O� M�!�R���DC�F Y���_��]��~Bd�"�Wʩ�3�@�H`-���� *���1|SB����uN�Y�.���e�
����_9G^&l$�* ��PV����( ��N}���y�Y�q�s�C��-�z+P����J�#Z���<|�Eղ��������x1|�k��F�X3������$M���>��ᓭ�^1[�Xu��!�����x}k	��֡㗾#�����uD��-����W���7Q��,�T|s�%ǯ���;x���$G�,�s��>��o1_��d�IJg���R^k1� ]Q�����g�x�����>0�>��96r��ԙi�"ő��l��9��DPs�C%ЅW��sdR	r��}�����\�(��͟;��_^����`>]F1<�D�<�2�ԭi�)S�"�e#a�ؙ/�/g=�]�?*��I(�J�T/r��i�r����LTa�E)	����٨-a��;�To߰�@s�7�eA�R#�v5/�8�>V���+�Izg7Uk|u��A���e}�D|�n��rפ����eV��̳�k�NA2yUe_^�'���Vd�~P@O�g��1�5�Y@�~��(~!d���)ծ_��~���h$KBe~�~9��q+��;���5{1R֘gB���4=QNؕy/���}Ι]pc*u���3���:���C�TM��̴5؏d38���z�5��E�_��8��XwuR[4���6�:r[�l̬�q_��2Ө��Y�E�>�8<�������z*�&�u�#���˾y�N��OSg&r��\V�J���3����+��ї�������up�����(|
'K'�n��w'�7���=kQ��ӯ�+#����t�j�Σ�5�����*�A2zB�k����c� �������к�v����u�`�tK98:�l���r'Ѭ�Rhm��Cs���Ϥ��l�Ylﲭ��I$t��� \s�G�w��d�c�N�����z�x�z��,�A8.^{[ݷ��\'�3�y�	����0��a�U?��.Ӛ~�u��&�6�~�cvǞX�Y�xX���'d��~��%��-I�L�B��$�9���i���"i�]�E�;��)pz��"9�@�U��V�u"�r�S����^�7�I>��L�M�1ݳ�����IAޞ��,Z|��r#G�=�a%���s :���Di1c�"�|����<!��J=�Ю�V������b����^K4+3�Z��\�a
�x����8��u
7�8\�Zd��}ס8��R��Y`�Kd�Y�p����KC (IGU� UP]ް��
S"q��6�m?�w϶�2nM�3�znzϕb'`����X�ј;���ޅ�2t-2���_����m��Z�U�BBy��Ћ�K0��0����"��c#�:�?�;}��;h�Fa"n�}-s,^2���T�,V��T�I�]B#$��4\ }��U�U�/Γ!$t�� f���GA��]T��.�P��5R�'Դ)� 3�[k���Ǐ�F.���d_���K!�Α#�r�d�I�v���X�����t*�-r*ƈ=bC;v��A!��,�8�,���=)�B|����[χ� ğG�啇�W2��Ǵ��V7�]�"��Kb�o5�_<LTS9}���<�{�� ��!�3��?Y�@���zl8�͍`��2�_B�/���Jo^r3��BS�;+�j'k=�`u�[���i��ԩ�i�4�خ�g�"@�F��VW·�bAA���'���:��U�;կ�,�<�$���V��@s�SIK���9�{�#z%a�͜����>�P߀�v�8���im~g�A3�*�E5�B��!5(c�.�A�WRJBIL>ܡ��s�H�i�	��`xƔe"x��-փc9�lDf�{뻩@ �7P������*��y���p���1p��6�J4��v^k��.�ִ��&��wt����,i����C�û#�3�$��������1�$�w	����v'�O����!��$H�J�S�u䗶��zѰ��Q]���UN��zaL�Y�}�J �Lb��kk�én��}Ӏ�TH��2�-vl�~�G?ZK�a��������* ���m=H������Y��`T�5�+k���S�޼>XK�q��r
�Q8\��.1�ϯ�R /������Z�e�	s�:Q�[��f������:P./e�D��/rwb�3.����H<>h�'W� �
��O2��?=�>��%�����o����q�@���N�ܣ\(���eݒu����/�֣�%��e�(�)Z��!_�Gi��(_�D�;���:�^SحK�/��ٚ�.�Z�'����9[�X����0�R���#�`u��n�{s��r�`��.^���d+ķ�^�a�[5�FF�yZJ~�v��kvȳYf��o�؃�+=<'}oN��bZ��V�2'��{邱B������q`�袝
�a�A̖Kd���?���>�/ڿq66�?�*�~Ռ ��+u��r�N��:Q�����l�v��6)�B�$�'`	>�����-t���:�9h ma�3T�2*ҍ�b���I��!�D(��.�#i���u�0��R�/@���:mO�ho��&��s�5���������+iV2��|7��T(#a6�(��M[�VuAǤ�d�a\ݟs���Y�+G�������.�,�F��[�@����[3se�IO�]���d��΂���<"�Q��޴����@�K��� )�E�P%e����֛O0l�����4�b��o�	�>.��ku�mW����e��I}؏}�˫q�ˢZ����������$��0��^�H���"xl�⤧��aAs3��c�����R��5��f J���pٱ�U��E�y�cz�_�\�*Ů�P޺Pܨ�?�\�Q����%��i��x\�L�4�B#ifa�+b���K�S����n��]Z1������4d��K���r:�����ԓ0��x�<��9N�@�pܧ��e��Q�n��6児l�^,�H�����~�Sog�xF�$q��qPU����i0��:i^���x�i�4܇� ,���[Z�eHg���?94��t�%�yfפ�ѝ�K����X���Q����fQgB*1:kK=}����W+[C��pS�4H�tT�]3���57[x8lOcӆ�3�z�J�����'j���8u-�K&J���j��i�/H\�(l}0��^��趶P��T��{�7��W���_���<<�֚sru�M����%��Ο�|S�
9����l�q-A��=@��op�C�#���[Qɧ��`R�uА��Ή�?Z�Z
�-
�	J��"{�uP�Φ�ztI�p<�U��i"�����[ֳ�$�8Pq��)x=�gi��1���zzQ���ۅJ(�j�¨Kïi��HE�|�/�$�A
 �ؚ3�"��w����G<4������D�܇��G�V]k��������1�8�iؗ�@Z?c~�n��t<��>��1{_>,��U}R���i%�wi�H�ԋ�`���[������W�ߔ�X��{8��H��|q����O?),b�'|�����xi�d��c>f�[��|q��k4�%�e�LLb������ٓ��E�rq8��M��bi�T�թ	Q~���3��}xy��Vn�r=�W�ۨS&� ?'������z/̄c�u�3�^�\+N&��=:t��,9����PvdO���<[�����=ι�{��1"�Ve�!�YI�v�'xB�#2&J�cD�Z�J~+��L�e�
��������Ob0���_5�Š7�@3���̣��g��3���N���i7�B	G�}�>���lQ"q��ru��o�� �+�L���BW�-�o��d����3�7ܽu&QWn�[%�"�"[���D�vY�����"�Df�3���V���-I�j�5��t�ţ�܃Hu_�$ �s9	BL�H��h�r}�z1�튣"T�_�wS��P��]��)�%��ril��皍.좝/�+���YEyٯp��� o&UV�V�������Ha[�"Z/�j8�/Ϸ�<�T�����.�@��	��SQ���F��XId���|��g�T���i�c��S�Ԙ�?�<�����\Unh�6ˠŷ��yJ�.���-!����CGL�����9�隣��R�0E��&��2[RT�~�+)�YL�����w��Y�	)7�h�?��WGz���hO�14!�<�a�Syxı��@�,(c��4�o�~����;�����M8��|�EGc��1�4+x�\k��N>I�%��h�u|7m�"�yt���!D�9�=y���ʘ!��ےLp��]>_9(����*�5d�Q�����X�� ��m�9��V�,kC�L�8�(�`_`sv2��̡(����SP�;d���ǲGb,��5�Ϋ�����������?��l�0��utN��g�>��"{P���}���oX����M�wUg���A��Y�	J���O�4v�z�R`;�N��iaHb�P K!��y�]#���eNڌ�ͳ�厎cg$e���p�n�$��r)�V��d����m�l�U�pۢħ��lL�;g�hQ�d���5�6��c@�@H&��T�4�esa��ϝ�}bTΎ�������#��$��4��RLm�͵*�O'M�okn�ߜ�~�Z�+�4	�Np�P�=1V���.A�N��m܎�	G�zd�}oS�#9�*����Z�eբJ�Q��{[$<�<��1ܑ*&��ԟ�4#�@Co���{�@��}FOw�0;����Rqy���A�={��ëdX>scе��{<�>���F��ȶ�� Կ�v�v_�?�UtV���4�,�!U���Z}�Vi+��ہ���=�;)��\:�'� A%�d���9��#ť�����࿳��?(��*�v�N�[��t8�(Ȑ���'̃Ϟp	l��R����N��Os�%��C5/�91_kr�z�
��h������P�5���X���
�Յ(�Be'�3a3 p�%�G�����t�ML�޼��=w�0�#L����\���t��Ho���>We$Йv���:_	�-��yNP�l/��.�QGk�B}���RXE\5�3k�u�k��8��� �:�[��ݓ��_%O���G��-��s�[Fy�bZ�Nƀq>Nc�t��~�M��ZY�ΤF�����!���u5;��T;%��fO�Bs{���9�h��i����S*R��s��T�y�VZ����o����]<�^|Ug�3��x���_�}���y�)�>�]���|�=Ό����U�n%��?%�Ǐ��$���L��Jj9TY,�7nR����)T���M���F����7�ou��Ha�'�MH��Rc�XٗVw-��J����h׉��9#I���z/��ܛ����X������l:)Yi?B1�Ndfm^Q��1�>�<>�7�M��:�����U��>���M�|7+����l�ꃮ�]��#<[�Y��?]*O�4t��,�S���e�٢�h��赺���1��y�vq�\�)`����@<Y�,�K
�J��v�;�eS֑ `n�v���GkFúQb���͹C���֔��Ļ���1�����i���a�^4�aד"�jT�J\Y-�G��Tih��N���w��(��:5ť`�d�������49��P^���~0�}i^	3�x���@�������	���4�ǋ�f�2
ث`�W:�F�����r ��D�7@���@������vX�ښՔ&�
��Ak5��3�,
(dH�K��V�(P$1�ڣT�/9��EM
����\�O��_C�,�C�_d��9����'R&�'j(�����~B���)�����*�F����c�n5��DzOY��|��)9�V�=����ԽDdF�Y�]u�E7a�%2��t׍p�����Zͫ��T��r'嬀!���뚖�Q��BM^]�v�qY$��%���zk3����h?|�
��_2z�r�</��@��̽XU�oBZN���k��uA���gp{���?j���\�<RzrR�O5��X�r�-q��W�cS�����PI�Y/�]��E`����3u�Q�;.�h�w�ba6E�g@��z�tX�nÃp��,�/�a���X�-بZе�-<���0{XBkƋ��Tz�6�=���Ϟ�nU�a���?���~�T|����8@�oE]�eXf=V-$��	��C��Q���Pia,6�%Y��d2=N�s=���i�}Ώ�!s�����St�0G�G1��?���sE�yJ�h����2�k_�����k�v��L<ˈ���)	��B�h�~�Pҽ�C&E砶#��Y;�m��G"\�5���Vŭ:�F
Ehj��m��:��1g��~ mKL��%��a���ޡ��a��9���:TD�������	�-!-�+�1c��d�b/�|\;9��t��<�I/2�c;��;i��3����?xn�&+��g!e� ：�Û�*JYe[��B#��M-8�x���e�(����ʍ2���h�͙���+h1�\K�/.�K#�U�;h3{����� ��j�n�&���2�ޒ9��֮C�}RvW��"m�l�@�R�v[$#8QU���BUMx_EZ��]�L��?��u���G#��j錣�:'
OiY?{�Г£�&&TMc�Z�*���x�i�8U[>��	~�Y\J~ s���R�f�l�iy��Kb����=�QrM�$�\�������F��� AV�y�E�A�`���z�a�
H JP�[Nx[���`�\�uu�`�E����V�B�,9��"���љ�������z�9���_�v ����X3+?єn��_��-�N?ҕ竈80�n�Α��җ��G��&�I�3�)��t��/�a��eYZ�ݶr��k�~�������:/�r�b?rgC֘��T�|��s:�S:��U����E�N�r�A�6l�=Z?�~��R���G���F��*�Q��)������T��"���_졥��j5{�O�����q�M�7r���D5�i�4quD���J��=_����t������"~H� ���Z`�%�}�Uķߒ���d�O	Μ�nL���S��UCI����	����F[O�%����j0�<�;��T���rp�H�����-_;h �ܐ<���
�[4��X`�m�bgj=��7���{���K)q��Ǐ1�=�q��T�
�~��86ұ�Ӹ�`��o���;����ض������$�Ha�"��39S���2H��5��Ivw�Tm���׮�̀�t�t��_�A�
H��]��W!��ޖK�XS�Xd{*HN����|f�W0(�>�x*4����j��,�Bc����3ѣo��;�<�!lq12��p��wy�
����.��4qA� ٕ�N^ҩ��;�/�G��a���w���O�H8]����	qI��� n�pv/�m�ЏN��蚌%d�۸z l��+�#���ݠ�����"ڦ����9;r�����+n�k�1�ɤud�ⱑCk@��M.C���dj��稥o���|"LAц6���9��S<r^�8O0 (��[���C���gzk��xӻ�5����T'-���;�JnJ'r�X���fQ��P�d �����W�����䅿c4�$Y6)�'e��vR1�_/��pO�m�<��"�[�/T��b �,π9_�%�3Y��>��X����J��Q�,AVTg_���o.p{��;�Op#�Ҏ%���na]=��j�_޸b�7��	=���Y7�����J&4Kl�@k�	��;�C$[2��ʹQ����Q0�֡8kv-9����?~g����j�a�Q�y��]h�X����M8��Z=�i2�@�����CgA�˄d��9U���B[}�1+l�p�.�lӻa=��o���o����U��l��V�Q9����D��A��,��B|�̩�������W��p���Yv3�rn�-N+Z
�Q�����gmLBJR7l�G*��la��H�X�8��7ϖK<w�T�䉌ޘ�3b[X���Z^v���J-�'�t�O�O��7�N	�D�T(�ߥ4f���W��%+Դ<�w}��/Oz� S��4�^�����d!�:&3�p2��+��*~�Cu	��ܯ"�9�w�ka@]���vIG��������;N���)�2��+Or�e�	�="��f�'��q��E�Q�
e��ҬD��M��rSs+w�"��x"*��15a�P����e��D�8Σ��u|�����T(ŭ������� +�6�0�	A*��֎���׵I���&LMY�, �3"@�Tݓ�][��k��x��(jK$�RmG�s��]� @ZZ����"��.1t����[�>�8ŔA�y�	1F����?�ÿ�g@��]�բ��SO	o����5^�D�$�r�X�R�!K�\�l����k��'�A� �_��9�	K��C ߋ�(�m)=��g3f:��%�������� 1�_^(I>���#lգD�\�;���������N��&=֚���B��x7*?i*�0Є�Ct�M௚T���Sa��������O�/�ϩ ��Q_
$W}��h��T$w�g��Z^���Kϱ*��x��L,�?�bg��3jve$1_�CB%�:�}�.��bC�z�D�<*��1�thnUЯ�R� L���6�?;�S�>~���Th�E�{%r�r�e������rV��F��P�OD&8��d,���8���M"���.��+�He�qɄ kr�W��Sw�4����{�ħ�1��>$�{uuu�[�������������~���M.9Xj��dKqDj�^�;Pr�<H*w��h� ȸ�s����Wظ���"�6�����-*Ie,��l�����6'g����47Y��=��SѤ��Ѧ<�S#�ۂ����L)"+U�	�� �>���6����C��P�%!S?qh�
�P�
�a{�	E�8��K�Z�C��.�V:����K����H�0zH�Ί=�:�+���T�ަ:���ve�jOv��t�r��0��P
P\�`�[ރȋ+� �ُ��TP�l:����s�Fw�����t����+��(��Q�G�#÷pDL�#�-h"!#'��6a�l�{�y �>F5!!����(��f�Z���C�j�(m�k��	��3�Vc>���eVLfő�S�����5�q�n�i�M�/6�RL��`L��m��ܞ܉!6���I����/Ӗ9�����j�o�x�z��D�s�S�I؝D�'En@�m�zl�����\0+m�H�X��zRV��w`��2y~Y� ���fD)�O����=!��Z���uk���c}@���ivB�.����=�MIZ�&|�G�9�m��'{�.���g�o7�j�ᥟo�x�+x��
��&R٘*u���*��u�ۙ7b瑷��r�`){#��j�/�O�^��l�z�o�r�K �)�|�F�͖��W �ۓ�C�� ����
r��V�~�����J�D�]\�=�pF�j����IJr�D�㹳�����J@-���?�A�������RtV�z�M����F���˜�:C:��	iDZt9TJ���Q��@{Ͳ�+̀����ӣ��;����5�����'�teP���+2��1���t_��d�T�qr�+x��i�P�{{+>�l@�0����g�
�$�
J%h\;�@|��5�.��x��������
vz�O�j�����i�r�ѫ�i�R1�hY��_�^�ć}�o���{�TlD[�!��y�~2�iڶ*�c��d���h�@0ij�yw-np�Cw?l�Й����ю�a�~�U�eH�h�t�"���Qs4�'��� ��֬nEh"�� @�'1}�w+n�
Tb�Jk�wU0��f5Y���� ��za �
�2��Q^�޺�L\�-d�C�09�X�-F@��%��� ��Ny��ڶz�v���w��cН��n{�����QSmG�	��I��ђa�Q�*!���S~m�eB���/�K!O�(�G}�F� P����ϝ��H)ff:T"���b��l2���ۑ�X��t�n�V�+~.�7�q���);.�u̳������b��BK��^b+َ ��Vz�]t���X��5