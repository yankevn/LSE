��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���!���	���V3�n*nL�\}]��0!4�#h�o�
5��R�U㏖y�~Rj{���'�$46JJ_�!F�����(������2w&k������3]��tүJ��$���z�Q�P䳨L*��=	��{�h��Sm��w ���Ef~���;��qCі��|z�+�t���z��m�\�_�\�����|� �_I
hG^�9�X�� ��(R|}������Gh�J�M��m��D�i���RP?�h�`[xW��O7� ���	�#J����O#Cז'n7$�}�"B-�FO�Ƀ/�j| 3� �ݪź��B����L�r*��P6	��O-j�|Z�p����2��gm���ؐ�ly�ӌ{+Gj���g��ޔ_pH�,����f���ׂ��̅2-n)+vȾN�,�zϽCa8����^�l}�tY���:�ֱs�L����tN���igC�h���#r�������-�,/bs;1[89����_y:A
Xe*5te��S4w��5���@��M[Ț��(���>5�0�ω�O���:~��}��[aŴ��)��ٹ����l]��5nA�s\3�Ĥ:�9χ@W��f�pp�m���xw{��h��Ũ3)
��*\�=���u����%2�_:J�l�B�m�������4��_�����[�=�Q~�g/ QbU�rS�}Ki��A����S�צ�0|$(V����A���`��4�az�o{���0�;���k��7��������8���W=���o�i��l��d�S���!mXlDю��Hh�Y�$�|ϐ�@��������xR�}+�tz�,i��8X�&����6�a���r_ʃ= �&�[�Ru����y��H������6�'SFPQ���ZY�7��2>�g�_+�3�@����ɧ��IJ�rx�&���|��ޤ�c>Y���6�9�PA�)�hh�c�ed�$z�����C�nЁ���ea�n'd��`�4{FHҼς=}����׸*d"�B�+m����y��V$�KH	 �}�|c��|k�KHOBpg���1�1P,�h�|}�	���e[�?(��UdQ��,&��w} L�l3��Y�Ѧ퐷WYʲ��1va7>c��%(.�@&T�fCn���c������$&j�E1K�/=����vx)6�qZ�+is�	.&3g�@�{�5��ѣQK�mH�b":n�G�G���b�|��L�X��P\�LO[LA�i��N;	CT��)�� m���p�6�QP�z�j��6��+�i�r���{�
yP%�+���H��e�:8��54���1�X���DPnT��T�na�'4�Ҡ�KX�����YM�a2���VvIa�
�f��)�ŨU��J�*�� ��O�2����x��^n����Q Jv���\4�?$�-h�(v��<7ŉ�BT=o�t�%�P���=�z[��"rͪ(]{�O���>�Ɔմ~���T�Ъ��X5������������S9Vo3�Ε�}��zq�H��?4��|IXΧ�i�����d�����H X�{)NkUslP{p'��<��K.��8�Wiɣ#������_)N1�z���#i�/@�>^`�����y[^�/N#�r�-	���>��˧,%��t��˔'+�fNF#�Ǥ���6���t�	C/���+r�)-sJ�-@9W�M��/Yg4�>�Aװ�@ڈ�!���"�:|���q:���������Ε~��Ql{9 ��e<����z�0���j����=#}�����$T��a\Ч7�3�K��q��V��k۱hmk��y�-c���CI�ptr�W9���[�+���u[N[&U����)��ofE�-��#t��n���`!�5�Q^�X�0�T�