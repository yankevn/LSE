��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���!���[��c�L��Y�w����s���\�<�p������%�6h�(���=�+U�v0�Y���Z�~����@��⌖k2����<:x:��U�L,Z�{1.X<G���c��*'6�ʄv�=�N�n�D�K��.$Lhߙ�D��u��z� WX�[���/N�2(x8d��� B��!�jWj�I�~����߲���)�5Q!�'�<��_�tbmt�ˣei����k�fXlE��d'7-�3�F6��xtz\�u~��}F?��m6vख़�>����g���q��°�~��M����{m��{3���Ú�0G���� ��^˼����FC"ci�³q��xˉ�_ +-�X�W�D��L�J� �r�A.���k���R�^΍��l����Ïb��$jB�@�5��	1?����'1E�?'-�V�#��5sye��&^}�RR��&�ջ�����Dx�}L�>�z��)�������
��R�*
v��3��3��8��ߔE�����oWQ���_�K$q��v��)�3�^>,��Ԗ3����9%�⥶�}T��t8�S��C{��*yh�#���>�ϊ���$�~�V/�T�G�
�Mx�g�`-5�|߁���F�W��RIM�Sb���)���s.A4�|�fFkG�o��mL��ZZ�*�AIq����u�J�jOFcK����s4� ο�)��8���(MCI���5mFL�=ƾ#(�GnW z�*�w'��u��\^���s�rm���0D(���J��9Q��+7Vr��[#�&[���!���'�\;��qM���s֜��[�O�\�K�,���6ѹ{��؏\a���E"r�n�L��p;ŇPu�f����uD��ٗ��,Ka�)�J��W���W�ʮ$.��q��O���?C����m-B*bk$,
�+�q��c@��3��^��6�F�z±Bg-,(f�{�#���&A�C�dU�,kj�{��g>�h��C�J�DL<��CC����0���S�Ѭa���7Y �}���a,��z4
4
o �"��!�](l���
�䍠���( ��[����
�S���^m
[!k!�!�g,�D�����UQL��хv��J�x��MGA��b�L�@j���k�D���,m�Љ `'4S���{x�)C�ܤ�"�U��6K�s�6� �?��%����8���>O��2c���Y��K���ϮG����fCq\�3��@��>b�����.I 
~�����{PlL/�f�
�@��A謴���X�\�]M��Uf"��Z��9|��75�y�|���������e}S����"#M6R�*]�H��H��J��$��_"OM"��qJ�VM���/?�	;�����%h�տa���ؼ��ۿ���v�9�d2ʦ���s���1��8��M2��Γ�v����A(����?���[.d�R��j���A�����Z���Hfh���Ԧ���~�C���