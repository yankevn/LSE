��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S����)1�
��W;tI���n�R��I2�p�ݒO��ͭ��g+�۲h��*���]��L�5= 5?ޭ	�6*���N�lg"�a)
|��+%vքj
�'�'gެ������[txPf�n�����S׀W*�Ǐ@��e�������/�1�)�H*u��q���
�>���qf8�բ8��F��U��B��%�&Q{���IV%L��>�h�'��V��k�2Z���;��o���m�(����a/��϶�#\��O�%�i�E���l�P-�����6��l���  ϡQP��~ ��FԂQ�u��8�%�Uf�1A�p,:����]�a2
m� �	ף_���Ү�Մ)��	q �P�dP�����C������zk}�����W%�_;p��(^�r��K�����M>r%pM��j�����9!S�y�D����2�l����4�=\O�euU%¦E��̋ϒ�WKl��#����f?�3�@p%�	t����ƕ�^�YG@���C�
tҨ#��G����9iI�_�l�ɝ+�4z�MҩC�|&x"��j QD����=���y&ʻ�Sl�T�ĩE.��۝���!*Y�[c�T'���C��"�q���j-�ɴ�.F�O�M�XG,<ѩ��4KifN��0F xssS��&%�k..�����V�屩#b�JE�fS��
<0����i�Y�5�_�8Diޢps d�����
��< 
אv��QKmWL&�󥯑Т!H�m�J��z�}�j���R>d}��)�ؤs{�$p=�J�+8�^c��KYd�~W/�2��|i�+/\�`�2�c8>�^v��q&��]r��Ac���fOoq���`?�{j��B=5_WSE�#5������h��1�a�|T�	��#�̕!�}�D]g�T��j�t�]���O�aͿ�=��O򁇷����U��(R���Uif�Ԁ�Rl@�ߺo��`BůdZG+n�@��x(.k��=��f�5 d4�."�_st��Q���}�cՄS6{���-xQ^F��z��l[f�9�%�ݰ|oW��K���!�/�B�?�st��x� <1��CQ����/���1WV 	�|VҵA�꣜.����K�/�C~���m}�b,kӑB��°G��Uv���b�Z	}x���{]�(Is-���s�r�K�/ɫ�a��� �0�Y~xvQ����8�PT����%wf���yB��T|Ѵڰ�����}`r�ݠ����	������G�{�t���=W]LL�E<8[�Q�<��M+�%���W^����-\d�`�p���K�<Q�U:=F�H�P'v�˶S��Ed���p����2Q��}�K{  p�����Te�a�,�7���O+��R���%��F]H'kl�g��A�f�L\PB�m���Qؒ��1��*�M�N�*;D����
���'5sBk~p���r��-����]4����_�]�iJ�_�"OJ�����l)7Li2�apn� V�&��J<���^�NK�٥q!h���ւ#
�":�N����y�2��޴`خ���eV���yù�6���!��A�*���6�m%��� �dO?s���קv���`�����5_���Hf5����<���?+�RX[���|Ů}><@T��bN-[����)1�~�
R S����x{��e��+���ܒt񁂀f�2�M�y%_�!ț`�K�	����F�����4�TM�y�Ȇ�RWE(@����''���y)+S�ٕ\U��M(�^��yex�!+ wƄ�N�˸�Ǌ�y�����Հx o?�6+ �|؛�	�U�4��؅m6��7~f?��s�!��K��%j�r�i��&G�b� �����U$�6�:�˩�����?�R��?�G�a�� s�[F�k��?�4�SH*�x�Fov�H67���̫J�nz�IF<t/A$t����b�c�ʜr����p�j0�a�M�d��r�oE��w��ˇs?�6`\ݏ�e��b}FD�O�. �4k�ùP\F�}��J�Xz�YgUkK�� �m�E��7=fY�e��j��㳁�;h{}��j�Z�F��� �!q����L.~��_7���k��G�FՎ�ʼ�w�]�Y���v��r\�����r�6�MG�pI���?� w��Q�/�<�$��c���T�c�Օ�t��<'1Gͬ���Wx�Ý*�`�L�o1Q�
\Ќoy��P$�͇�"�$^#��[K�5�Y��f��H%�'~��+4�%
!�bw�Mr�%�$��'-�N4�o��� /W������K?��hZ��ς�'l7p�0ޏ��|�? S�g	\Zt;E[�?Pusߗ���ه��>��Fc����L�Ek�1���	u�\r#Õ�V,�_��L��
��,�>�,�v��_k��W~Ն#gs�_�[�D-�	4��3+�x�i�KF���� A��GdkT�<�_J;�,��C�n�c���
 ����ȀҡE;��CMp�M>�+�������T��"��6J#����:LD]ڛ�}髯M��yzC��v��#`���޻�	���aBK{)����ŒyLN6N%�1�\6��V��|݈
� �"�ʑ�AѦA�������}9(�˺�x(�w�b���VQ�~�H��`�+V3~Gܺ��,ؖ�Jw\u�Q�Ia��!��D펙�c���V��(K����_����9�鉌��`#�!{�|
�����纭s�s�.�rp_��LO�2��'�L�ێ����{���~Ð�ƒ�N��W�27�>m�� =�CU�)5�R�W��Z�)(�G���ʒ���˰�-�:I� �bN@AD�9��aK�.���9(<��ڊ]B��ֲ黩����T�h�6�� �ɔ��^��ߋz����-Q#|�є�n�(���*�}W�)�7����Y�2?s�����J`�k���ff����U{^�Λ�o�V���ڹ��.?%�����!d;��bt@��P���o�R#���ڊ�ڡQң&)��Hx
�$��}�%#�J�H��[F\��mg�]y�}g��w����?�}g��5��v챟�g"-(Y�d�,*��u���~/�/��i!��)=��	D��bY��Gڥ_�^SX�<�d�i����*�CV�Sz}<0�\�ٕ��.N^�oN#�goDO��MV�^��L�Rts�-/�8�ti<}��wq�E}�T�H�\�`LV���� ��VG�O��:�nh��ZI6�3��G�9!�!9�qI#B�0��t��}"��??5����'�A�9���_AE;�Ҭ��B�; |m��"���tT}�{��J�YL���!�g���QAӯ£�pp֙��Lm d'};H$s�O��3�rp�dO5 � k
�Ym���x={��0�.��Ƿ�Źaa�5�X��-w���-')���/�z���`�RE�H�bG|����9~p�8׵ĶQ{~�\~�SU��ߥ�GF�VDm����FK���}�3��h2W��>2ÊN�p����r��$���S^T��ȃ�B�^��������E:����w��[���U=,δj��Wj�zT�?��i�voE����2��w����K?�F[خ��jsd�?�=P�U��npR���[]oN�ʏ?k�n�_���7Qz��Y禳�k����Ќ�����,d�]��`;jd�#�
��s�j��w|TW?�f�����;f�;Bai������P>��^�^ "k�WBr��ŧ���M��ԧ$Q&����v�Nh�`[GCë���J���U�D��=ۘ~]a��5�	��;��/�����{�T�Үj�|�{a�ƽ^���0 v�[�}����Hp4d����|⢶�7e!f�o���)Q~a�{굍�uD�������"�h^:��<�^����`=[9��Z�(������w�wX2�����_�h7�=��������*���l�պ[�(�"�rjA���.TF!r| ��U{k_�!X�g��ԜpGbʶx�Ҁ���0��^Ǣ�> $�r��'�p�h�_�$4K6�*��H�d딛��3���n��]2M�"K�7k�A�ֲ^�N��w�{H��Y�I�g�8�����Tҽ|�ٴ��[/8Ca�şC&������V�3 �ղ�V~��Xm��_聨 �z��������1a��}N^�e�o�dYh��DżA�svnz�\���ֽK��E^�ֆn���5qND��������D��T�uX��_	ZE�c������fv��T~��yf^3�]o4���^���� Ȧ'��&f��>���������Zdb���*
*R�k>ГiW
�f��}g �{8����5ҷ���B��v$��2��XH��p�+���^H�4<W�J^��=/pm^�0��=���\ཌ(g�2����y�
k�]��'l�,f�6�sx~�
G9���fH�fl!T��P�g�n9E�ٺ�t?��O8�C��)i�!�\�U	���N���#��.��ܙM�dz��e�e�s��`s��u��������	ɝա��	R�%��o��K���$�[�=�:hp����;�ɚ�Dl����x`Z�D�XR�\Z'��a��jr�A��Z��	ΐ>�����y7T�Q�i�@J��b�,���Qf*��`�{�:Mgr����>�P��;�Y�$��Yʭ���P�[/����K���wp  K��T�@�9�}�f�B[ar�ß���'�l�:�?d���g��睫���Y�*V�Y���eIn�[8��E��S��r�ÑG��PL�2��kP�S�qa7i�%��?�8��`#%P�[o�{�sD|f5TG��ҥ�,�mT6�Ѳ�O�<�@
�}Gꊋ@�Q߶ւo���Q�B�����y�����D�{���O��r;r��
�DF7���X�ބ_W'o����+M������5�~`>��ʃ�V�~W�;[R����n=C�(��p�G�Z�5��5�|)q����h��'���dndbo� Y߻��?��.��F�W_��=��������?�>��Q�/0�y^S�����`H�ip���DC�U0�����|l���s���B��"�?Xڐ)�lȥq����./����[S���"���xE���A�b��$����U&��)IF5H�.`��A.��,o���XI����
wFC�Ѣ���O�/L�Jqugn�[��ߞ�2=3-h����9��]��W��I��|�{ΕgF$Am��E��'�"s]����F�����`�[�����S>C� {���tђ(�B��o`ݳ��o������A��9|����]��;E;��g鲕���5�o�N���Q��ζ���;s%.u�ql �"	.�x�4-w[Ҭӿ��7�D1�䓏����E=	�����T>YFC|?})hzH7ٖJ4��ZDEit�[��]7�))�<���@�W��HU�eœ���=E\�;�S��!�:��G�R�>V��|8n���}�n^�:C�«4���������tJY4].�KE/�ް?�M0κ�(�ƙR�޹x����]#��%_D�u[��٪��&Ez߷W0MZM�U˛�`z�8_�l˪��>J��Ȓ�܃��M�Zf�1�C'�n�h��aɂ��ͫ	x�n�6l�����m���ZiV<&\P�vD�)���p�yP�\�f頲����}�����=E�Vh��;<'�����J-V�㫳�GT�Q�gB�z�&�d��VV ��*�[����gT�s��s�{"��ڲc�\)�f�^�,�8�����S:�C�\%���" �.#�Β�ݰ��3fu�.W��ڧ�L���3��`���oG�j�}���R��&G	V;Ȫ��w0���(�y��]ՙ�?Ng��1A�H�l�-�Q��w��huW��k6��g��(ߖ�z�;��Ki_&��9V}�����SV~��3-����O/r�@���8���na�2|:-1�P���<���L��T�5q�M��r��;7�
½�9������SD���W��`
d&�W���&SZ,�����g�D1�����`6hٰ��x�=@i�|���VQ��(vB�j;,�.�6�r>Oϛ�kE.e��qnͧ⮁�d:P�L��!/os�ڔU�;�[����|��C�l�`֣����D���;��c�f�	��f��`qg�'���_5Tor��.Tb�,;�1���vb��jSHl0�]�; n;iCY�{�Xsk�M�	�hNk�j���S ՕoKT�ɻ;�q���
[(�E/�����͝C����pν�Ln���$n�l�3P���ԩ2���-��Qp�%�~`�Y $���nI��\�f�G��d��nj�Ό�2�@�ذj�Mtk0�N�/|P����=Z�p�U=��:O��a�a��&�������&�y��P�������v��{����h�/�p��߸����,�IY�B"Vq��J|���%	��e��*M��mj�~G��R�MѲ*}s�&ͦ{�`a��^x�m_&]�QҪ��?M��Y~��)#$9�b'r��Aᾼ�����A���Ø� �j����>�F�� X)�������S���>�W��k�˱��b9������W����9��!Lם�����MK��`v��+�6WW�o9p��rQƄ�1
�Tk�ٺ쁿#�a��5�h��yz�> ����%�QXTU��<���	�~�,���R�P*��?=��ȃ�n���(�=2ur��h& x�0���@광3}%,� �>O�gzի7�L�J+�C��$zoC �+Ǖ�
�Si� j���k9Y�d���vv,���56���en,;P�Ӕ=���a��C7���N]�xo�VS�����˥Q!Yo�������u���	/�,	a兘v$����]�c�����ZY�y{��4�ֈ�V�\'V�o��S՝cE����ͥT�&�;�ިs�j[����3b�+�+�Еd]4痯�Ϊ7B?`�XAh��ۈ=���7!>����u���2�W}��b���jv��0c�4�(�<����Kw�"·>%9=p��n��h�F ��D{z�|G
��T���ra�l��~|��OPa���9-��Nn�3��F���J���ս%S#F1���A�?+�T�]�N�Kb����+HEF2�k��|l���թܘ�M�s�����F*�<l���k�f/m�ئV+�#Ur��.�A�}/ �K[ⷎD��0.1h]�r�A�,�w������̲G3�9ar#�<P�1�x��5r.-����ڸ��5p�Z���.ʹ��w�Uڞ~ϭk!�)!�z�B���-L���u	�l/T{O���Wl�5c�y�aG�v��1�s����~���t7��t��ɔ��-$�@��ez*G�^��E�J���ؾ5��{�*'f�%_��2B��S�,v�p�j1�;�%`5���$fAU31.�j�*ޮ��<?��Sa���.�2m���Z&��t�
��X����)3vD�x>���]��H��b�BrޫN��":@� �e�r�L<�Z��!	��{Y+q�H�Op=�����+��7W�a�,��1�Qln�����ҁ��՞�����@��+#8�ai��Z/�K���0�T�L[�doB���+�t����V�"�	���<��$G>JZר�<{�x9c��p�<�H��Wψ|�����/ ����a��ą7���T��7v[涺�h�t(d��*��������*/��Ip����cO,�<Lvǥ��>^.l�����r��������N��`I�F��Q��sَ[��{&�����^�8Af����y$���"XC���#���f���kq�`�T�0�*2�m����;�o<��3ەOȻp4�p�`I���V��Y��{K��s<��9Sqퟋ���˞Q#z�Վy؏�������M���,]]n��i>5�B�ay�GU7�{d������b69�hOo+^8$+�c��@��#��&���9:;:�Lv�P�a�D��XX%�ӤRTP���׮����srf?��1�H �Q�j�8�5¼��n�zI,[-�ٲ��C�C���"?u.����bK;�v�8W�ُL���ӗ��i�$�#�3��m��!Tz��k�u��&3�o���C�� ���1�ï�ө����X	j�{�"%�z�^�WcՐ���+��,س_Z	��M���	����G�[���pF*��|d�K6�<�	s�Z���H�خ1��V�s[z�j]8��u��0o�ßJ����t�6#T�/�w�/ȓY�V6�AzQk���x1����>��F�X���c�?��,<Ы���ޫg;\�D�^�T�#D�L^�i,r�@�,1��6���4����V���hkp�ů���H�喚!��R�}�|�<7���d���o8ӷiW�s��=�t-������+z�~�$I�;C��k�M�x	l)��,�^�:n��.�'�g�i���j�1��`�ZĲj;�����I�4���X��S��*�7"��9�����AN��"A	 ��?K��/{G���@�DA���Os�v̎"�;Q@�кD*���f="P2��X��j��Ћ���\Z�g�8Dv�ld�)14����R�5Z*���2�;����%�GA;�V01ݱ�t���3Q����!�uU�$��bO���ziw
g��oU��)Ǫf�#��m�vV������"��L��Y��Ƕj'����F폭	��m �֬�ͬ>��w���S�b������v��?��^`�	d��i$���_��WŃ��WNC�w