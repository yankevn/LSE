��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� �����
I˧:�-�Gǔ�=���atSƊ�|aui!?���c�?�/���ڈD����_���Hs��L9���)�_q��)���8B(V4c	�2A��u4m�����zH*&8�Y��\Y�ej�9��mmf�r�$j]wC ��� ʅ_Kz��{�����ۻy(b,������BW�X�e����c���pu\�����5(�"��C-����4���;�aL���������-?���&Z|�87(S���v�h�O��x2�S<~zX��K�p�������yB�V���Jt��{��CΡR�7?r�%-i½$RͶ��(�Da#����2����XB�k}�YO����Y�X��C+V�u��B{�w�e���:3L�\MF��0�.@q�ztM����A��%bruo!����.��4�4>%#@�O�u3�h�u��|i�W���.2`,��Xߜ эm��&��l)K�υj	Q����&�ϕ�[�
x%<���(
f��7ġ\>QPi])��Iq5��D� /*D��%���.�(q�Zj����XR@�7�=Y�� �0���se�n���R�Q{|�q/�X����V�H�����d����� fR�ԁ�}c�U;ݫ�b$#�-����D�!� M&�����ڰkHWն���<�>t�)i��H���I�ֆwp��{��� L/���@��3o@L���p$W��2���J�&�l�H�^�r��;U#��B.�o��A%_�n�q�Q��#���s��⽣J�:� N�S�_�,���&�f��w;b%[>|hW�k)�x�U�[�B$/Ž�(S���^d魶
m^Y���8CF���{�jYPqE�L��u�Ao�E� 3�R=��7|���:�aeu �Y��6V�ha 6�U�ue�a��wŤ�&���Nq|��P;�2�t5Ò��{�1�<čr��.��8RX+xn\x<<[U�iW�F��V��`�rE��N�}9����P��8�<g>��m�� <�sऻ�z�j5�)��C��LXd��+�M�g�VE�Y>a�b�I��Ϫ�(G��6���|�5����1B �O���)å�]2DҰ�@����bTD�@���}.�Bw_�Yu+0�b�d��p�dZ�B�~�|tg���ʴ��#�ZSj[�b�(�#�=���RN�8@"vh���D�c��5�|լ�B�	�R�ƿ�C�/=)}���e\� gu��Ϟ��w��b��./�_Kʝ����}ܜ�yU�� 쭺�Lvl�]F=�A�fs�<ehe�ɘ3!�l�j�5������������bF��º$�'�u�����ƴe�Gn8��?�5i�9;*���ab�66�&K	�\��{0�������yg�
xj{��h��y���,o$��9�2͑�������
o	w.��*���M�f�il���Noڂ���ԙ��&\��y��nӤ��Be|Z�n�S	 q����=1��H����	�s�����y�H!�:��D�'�|����#��ZeA�K�3���ʾ&�/d�t�W9��W�?����r�[�Y��Q3�ޔ��a(���]�
�G2%���aõ/�Ë��K�2�E�����B���i��x ��ƻI7�y��+=�E����7����yQCN�����.DTe�i�Zʉ�j�sdT�Z� #�T����U7\���4g/���w'ј/����w�ö��A�69��1�h����(ȑA"���13S���̐��%N��"O�,{�/�~[چS��O+r;�$��Q�7���HA%j%sU���F�W��t��C9e����E�C7L R���|�
�;?^�AԂbJ�ؑ$QS(7j���^
��O?��0��Z���_zB�T���1�c��F�Hk�<�����u��/�[%������=��g�	Q����C�x>���I���ִ���^{���
!��������T�n۩�B`T���-����\���챬C5�<�*��+�m��?��BJ��lm��r�載�8�	�u�@3��ֳ��qH�A��Q|ux|�197�І��ϐ��/��������S�� /ސ����=���>߰���a�fa�v�_��>�5�z����#k���E�)S_q���(�2'[���DUq	�S�sa{b��?��/Q��H�
T�m�_n�=E?����p#���~d�V�,/uO���v�5�Y�-�6��	�W��"m�^۹�Tg���='H �p�.��s�q)ʲԠ�V���m��&��G�{��b�� >��� ��4��D��dչ����7]s�6Mu��ͣ������G�gA��#*�Q�����w���w"ܰ{�����	�}�ӫ�J�,��E;��*�8�[g��K�F�96_d"��ê��Yk<uV�{���Q�1��L,`9C�u�'����a�2T2�'��o�v0\��QJ�����kU�L����X֍��,���`q �����C�0ml�<o�ֆ�MF���qa���}R��w��K�34����_����S@�nL�M�X��
����*�s�ab��:�#4$�G��DWr��C�xM������l�u�o��5�"��u9of|��ς�\���ؖ��9���wk��l���L�b�	F�c𦆈�'Ȉf�w+��IFj�:Ųje*WwWaKY�)i�$F���%^P���]IR�*�t=� ��l]K�TqD����T_��XUQ:]q�IOX����W�D@S����sV�0k)P�V�i9�Sܫ�������u�[�*+�>R�C{G,��C�=)�s���,J�w��O�y�?�[�@��� HR��;�vf��hH�1t���V��%���[��&̟`ĺ:��B�o�}��%ۇw��t��C�<4$�g4�v@r���z�<J��\�5PZvyf�j|`,B1E�̈ў>����e����+͟��F�J�D�M!��Phy�Β���q.�����v�zs.<�5[�C���|�]CPD4�H�nWr�A�k
+'����\b�(Y@[xNc5�&c֞�Fwk@�z����+�m�O�W4��4�Q��%$㡱�T���Mi�T�@c_�O��XE��Ac���!��OZѨu;�&ײ�m%C_�)]�9��u��P��67�W}2���.j��ҵj�,#����&�-ֺX�֫1����Z@.��`Q�o.�����������'ϧZ1]�Vﱎ�
I ��1Z7�����������v��4���� L��C��������O.��L𕥢X|����x�$U�e�^�"���ƹ�Z��6����XWM(��;m�X=x2�����T()��ԁ�pb@�rtL��u���%@_�����0��B��/��d��ܶ������.k�e+����~Yu{���2�md<^f֞^܂Z�@7�0b=�F�������h���VH�"%EB�/_LϹ��~yp��>W��6�ض�����v�1z>��puW �lGqщ�Ǟ_{K��ڻ��d~R$"2~�o���n��9�96o)�[`a3��25�Wl c��h�_f"�us�J%y�F�
qn|���a��Լ�O �H�d#(Z��cEq�[��r��d�У,j�Z޼��Μ�����R7���x1i�k���Qq���c��U=w���G��岼
6q l�0~pUG�lI���Y�\��T�}ٻ�"Nh�k�7�i®�۽�y�^lS��HTE-9�U{	�M ߉ܴe�{��� 1>nOz�tob1��l(l�A�E�]�=��,�݅��C�1��Wa�ȑ��+`c	����3aW�u�cSR�c%�M��x�������6}ｦ���~�� �Lݨ(nn|%�y��V�Ưoz$$Vd}/�ї�+c;��1���5]��띋�C�m;;>T�1p>	-���v��