��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�Pkk�ZK�P�18w^�9�u��0�3��i�?m�a�5�+���4���_����K�����x�}���0�$!�*WV��|xϮ�y�n��A��&�T�*�qY�q��w/������u!��$o36�7Q{"f;Or�̞��{�4�v�^��h$	��Ki4�,\��M��>Z:�BAǕ�d�׷e����Q۶C�#_i=���-�da9	��u�������  ���*�T]^��f:I�!W�������a��ʌ�v�"�?���c!��3��9=�nz�G���D�����/3փ�kv���H6���J3�KRY[|ε
H��&Mk61��`��I
��l�9�T��$d<Չ�C��č)��b�o��5��u�^���r�)�u�a7�"�e_{�\�����:��"_b9��8a����
��k[z�t�ᄉR�KU5�Fb��ϟx�c4����w�n�S��|M�yI�A��f7ҧr�2} �6͇"�MCF��C����/n*�a��f�j{�9.<���k����D��%:��Z4�.����L$�,���޶o}	!��i=��Փ��8����vt��?�ߛ��'B�PL�/wK�v���&�׏�d��z͟��4J�G��7����#U*`�
qN|sI=R�j�?��s&��sm(�����N���zj�6�St�.��O����ۯ\�7}�z�����n6Lj��/�Rlf��)�n�@���f��->��+��ų*�&���e�)�W�x�c�a$��T' �����И:����6��/�S�R� ����qUmN��׺��k��\d�nq�"�򿟷e:�E�"�Tr���1�~��7�b}�.r��I(04����^<S��Z���R�����M�idχW�7�|���Ѭ�)�ŕ��@C����gnZβ�{���<������H�y���M�c���m��qG�c��a�7N"s��%b3��g�䒯�LrO*	3�F�n�X����!p.�Bd����I"$p��Jo�D�rp��p�h�����-������Bn�[��i�Z�W��׿�j�f$�|-�*w���;����b@�����$��_��>���sD�mZO^�����K�xDկ{�O��t�����,D�ɟU�}a�JiN �X�/����f��f��^��ݤ�z ����O�i�]~xL���,i�Oi8V���<��t�F-g���W�g��/����!F�ҷ�Թ��#W;�D�nU����U@�	R~���)�2��<dYа!q�A_�׏.i���gv)R��Ga�V�n�&�RZq�F���EF�𲻝���Y�W� �.q�7:���u̓f2�H�Hؠ��Fz�)�����Ϥɩ�m]k�~��bB,;0�%����+��$��X�Z��R��Ԃ�b��Q�&hv����Q�O��c�km��%%o��~X8�|���^4�9��7�pckOY�`����8zpt�'˂l4���N��֥��w9!�D����=bTB0h�h��=^�&VA����=?�*v����r�����$���ŠzI&�iB�����V�r�9��A!�<�x彙C������pk/*T�ü[�qv�����R�-�H�$ר$�*Wd�7|+�+�|�el/A�LM"?S��gO��B���R�ݮ��X��� ��(al���ټ�V�Y�DJ�륄�M_'�9�X�*H��0�",.P^[��2��¾"���v/)fj#�+����2�$�K-�SK�����VC�R~���\�����f礱I]�!ܴ��F5˻h��"v���p�]E�,��Y�|�����+؃Sq<�R�l��e�9�Y����;���4L�;�#��M��ɨ�*�4e�vD�IЍ֡�"+(�h;w�Πd"bOO��:bs�z���� ������Ǐ��F��ٳ�J��/�&HDt��	n�xܬvK�t�IX
=,�c�lj붞��<��A7��N1�j �R��x�m;�wo�2�r�Sn_���}�� ������gy�UDgf�@��b��}a(��q�~h�f�}�0W�����d�Zg�z!,9�-�3��Y� �Z��~�]�ĩ-A�����YֽLu��S���ZȔY!�������@�z�m/o�wi����C�Fʼ@j(�8��qT�7y3+!���~�H��l��g�z� ��91
�>:ǣV�UI��\lͻz�0kØ�Їu�o�N�n�lÄ���!F|J�|��e+<t��K��&�-*��ә�ک��R��5t�Q�D<x���d4��0��v]�c���#��� 7�r�C�na��=������u�C@�x�8�5�DA���D!�V�U"h�����l �h��G�;,v�r* ��l�f�͎��Òj�Qn���7��N�#w"9�i��J;�*����N\��Q[��t��s��WI����{G�e٘�������WI�~��M�2n����>S.��_��w���r��{8�Ա������	L?Cͤ��]ـ��u�W�U ��b���￿'����2r���i�ٌRw��-V3�/���t������%~�Q�Q5A��~���L�q��sl蘅8a�G
Q��~�����]��YJ�`�/���;hGa���-W�	]�tJW��u��VQ�zҗ����ʭ���ړ��|W�	r��@���3:�N����9��j,̂F�5_�����c;����nc3I�-�jZ����o���WUZ��2@��������[��(�	m��>��0㍔�p	G���[������}+�~�쓝�����H�\��ֹ���8&���>��H�7�3����t��))S�a�1����dn,mX�2竀]P��N#ҨQ�fc�ZQ�W�1���Q���ߡrM����U{�x���<���J��d�2t�
N/Ż28�Pc���N��cQ]�@��o��a���*�]�O4�B����w�0�ǧ���ϚL�N���^Vq~�3���oii�Ez�]4'�	�F�-��Ժ���Jt�"T�f5�D�m�$�Qy�����hKl$���%���Geo�	�F�6W�MI��6���=C2LX�'	p�|W��@�8��2�7�A�����ϗ�k��Y��.}
��5֠����ֳHd�CǬ�@f����(̦���&����-�	���H\	��ga��0�!6�\j��9�������H�r^�V%�<\b,<q)�Y���W���,W�$ �NjWws��6��}*���C<?rR�zz������a�R�t��s�Av���-�,���G��(�C���@Fk�|+�N�Þ�/q���Z��ѳ�NUZ_oy�Ew'K-K�����vk�2��L1ؤ�4o�h�
�rH���V�f�����<�.���3��B�fa�����n��3�<�/$<�*���ޖsJ���%{����Q��i
s���Z��/QQ����h&�>����V��j�qU�ڀ͌`������h�XD��ѡ���@hB,�+��x!��}�Y�UN������Cm-3��A7���׳�| ح*A�(dev�Tvǟ�u��u���	�F����n��I�渝,�L�^\�M������_�X��CKq��	�o_�]��o��D�k�YC�P'�w\m�u���k�u��ř�4������!3��f;Ɖbi{i��}'^̢���}�n����f�,�UBu�(��o�T0ډ�2�2eB�2�<� ��s�G+y.�%�����`�7we�	�Ȃ�%܄��RN� 辰�R��ѭ���~���W�T��C��Ka,�K�� �����&|�n�KW��[�����$��<宂��{�������|FY�B�?,R<����`�Mgi)��f!#�:qMl'���8��~U�L�NW��42{�a.���/��Π[ě��j���5�l ��k}�_;90��d
��ƙ�d7�x���uk�tz�UB���m�6VO�C�B@>����#ثK�z��"ߖY����[M� o�dV���/JGҹO[:C��e9�7Yy�>�.9�n��ܺ���!�4*-�)���nU��RA&U^�Xp
:�xƟ��4�k8 5��'���&���G���u]���l}Q�bU���p��	N�jT�ퟂ�簛� ݷ!>��mq����5���2 [����r���Ha-��WZr�������dw�m }�ӏ�-�br���QԷs���e;z��S:(T��:�����F�6���?�����al���Wq����B1'�=^���c��m�^, �}��V�ey-@5�Utt)*}i��6[ќ��q�TI���@�È95�Ὰ���dD�E;^<�u�������
��_�I�	M�&�<�Va���oh�ޝ�nds�` ӱ�6EN�H�CsL��t��U9SP���^����j$�_��>���(W�{�2��C�N�B�4Ð�㱦rFvT� ��حIS ���#��L^��vDx����rB4أ�Bo���Ӕ[���0�L��V�z�3JZ$y$��6��B���[Y�ۇ�P��&�m�ߤ͘6�rTY���x��g��b���
!��a�:;� R�Ōٛ�X_Ys�n��!B,څD�iM ��H ��^�Ë?��`��w�'�=;ѿ����ka�5���蜪�����Q �ş�%f��,�#[��'�#+3��G�o$�dܽ�d�H����[�=x�����c 7����m6�j,&F{ma���&2���pP��$�̳���9+���d_F�o<��Tf�J"[��S���#�Rl�5.� �I� n1z�����`�u�����?-S���J4#�k(�na=��|a�V7d��--�)��gT=o�4~��k�߯�R)�-��t����V�`w:+7��˒��
�W�[����乔_���ߎ&���]�V���yiv}�pX+��XB^H�������s}����V�E�<��Z�,�*3]j߀�#�0��z��^U���'a���+�O�ȭ!���flEb�h8� �� f"�>M#.�l�JN���+~��Ô�G��mv�� ^{�.(�3@����B2������n��L`¥���V?�vґ�����,�0r3��e���\IbOY�l�	��E��,�S���(��Y��[|
�|��4�3�&�Oe�j�@-�_��v#�|�0���D��I=� �����n�Pm���z&<��IΎc�I��F�N������0��#��;G��v�E��o����2(C��e_��vk����Ψ�|N�Ͱz���MY����+H��B7vO'��&8Y���i��חt^��coՄ�q%n��9�
��a@�Ջ0+F�/��]B߯Pz��m��r,?K�#��2b���Մ��8�|V��\܂�X��r�$�yw�DN�JEl+'���| 	)]�Zu�[�8��.��yyg�[}�@���c�(�7��ܣ)�y��=N]f��5>����ZSȮ��z��(�8���޷%�y�l��o�����&�����3bbT(?d�*ps=�_S��S���ɞ���eC����R�G� �x�����q��5�&�wn���o���ϭ�;�p !�� ^?� �A��]��=|�ؚϱ ]�����H@����Ʃ��r��*��V�#��I�q��-�^;���h%�|ǳ��n�C�ҳ+��3P���j;I��R(���i��{�y�ۇ�����y�������#2�������Z"J���dp�Q�:��8/���%�KD�\�$p�UX�(��L%��Hx��>5_���LX�J������I�;�U���U�Y��*b>�Mg*9v$Q��(uAE�m����@�w�T#s��ŭ�����6�K1Cu'�t��~uy<"��cC��i�w�DN<����d�7�M��b�D����&��P6⥙K�:q��k�a�\6�����!C�Nxq5�PC��a/eyI1f����c}� ����I�?I�y��&17��D7!���Vj��~��h1z��I�b������V�"���)���I�}��*%�P�7L�6�	�m�k{`��ڿ*�0�����ٖ��&"�_vP��I�n�?;��=Q�o�[�¨��Z�[�,�/�A���A�N0 �� ^�.��UE2H����}W�N�9��)�g���0��vj�ႁJ8�.E�3{L�Fu����1,���r�������#Sz5^$��UM�`v�3�qF �q,^�`$�_9�L�	��ԃ�Y�7|��qn#�{Ɔ�V�YF�nw9x@��T �������cX��X�KR�>n/:&_d�6h�(�|���Ա�*���3R��(%�Æ�۲