��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,���D&ů�ަ$6n��o��x˱��� �*�q�\�e}#цr�cd.�_�٠&���M��xI_`	Jjڣ*��+����.$E=���1����j"���E̘��w\��jʽ�V��^sG`+p�O]��Deq���QQ��_ �=kƂ�Nd��i��[���)m�#4{��Qu�G�;���D�i�BY�j5Г�uvY���S�����7{��G�l=���BY�$PFӍ[x0V<g
k5��i��D���m|eC�T��,gm��e�8殾����M��!n�	�'��he/_�0�8T���(��~ЩQCM�0�B9�Oe@8�ux�\���į�����ͳb����_nR�:��YY�	�%��W�����62v�@��]���z��t��w�0f��j���甥r�f�7#6Ӭ%�{i�L�r�gv�x@�^�sd�LI(��ˢ�?_���jd^,��\3H�>��y�⭊�=�A����V�K1�?y���{s�:�'c�BSV��ʹ2A�H[F6��v��J�*f�ء��Qt��k!)ѧ%E�D� yA\�f�>ǆi�kAO��#�E-�"�z�<D �jz���$}p-5�;���U�>k�t�L�Q����o�q=�&{�g�
���A�]������N_��rt�.s��vN��ڷ�8���o�aK-�S�3�����:Y�d���!�{YG����4�a����q�ȣ�̣��"Z���|:Da�����3�R��N*L�r��Vv't��[�J�t��?wfn�
;��蹭F��$b=#i����[z�o�GOr�r"��~�+��=�
���3�}�V��:��TR!��x�*=ϰ43.�*I��g�1�����Ů��[֢)��db�i��EE)�w���z<z�@SX�k&�.�Q���c�Kmyf���W���'�*%s�n�ZX�q�o����wo�����l���9A��L8"�{���3?o�g��+*��������{^R�
J�2(?
�<��\��]%
�H]+�Q~lw)�`�<[���m���}z�9b���h`β��[Y�G�W�LoAq �N�o�$XP�.2�q);~WA��+�������/�oY��9hyX/ƚ%���e����c�H�F�0�yeR��b���!,�P`'TW,F
���s�Ap��լ�莹3A�A���W���fqT��}T`��z5�bx5�gHU0(P�����?� ���� �����������L2T��ҳ+N�����4�a�vޕ� w�|ʈn�o�Q�WQ�78h������h��6���b�,�#�\�%�?�2
c e���L�Pb��Q�U������������3X05�h��IIQ1n�h'L6F*>Ku��B����	��F8�ps�D�q�V�ە�Xh��҃j�qé�Y��X�A��bk��4K(c�2]������=W&��bR�/�2�~��