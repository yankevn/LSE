��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��z�B4j�$+�x�G� �H��$?R��7���tD)$\2��T�!������#h�_��F�����.K!7$��Z	ֈd�/{J����f'�*<�ԕ�Vu�-��&��66"�G�1���f��A�`���f%����F!2>;�gT�'�z�o�ϓ3���2����kE@���!�V��$l������
�k����{�˘��-�K�Uv�l��j��Ì�+�	,�M�#S0[ƫ��C�/,zLH�v��d �IeR�v��Ι޼��ۑ��6)��i������o���x)|-~U�0��J���p�Q�`�	� {�5p�\7
2#B�bh���8'��d��͋x`6.z{�u$�o��|,q��~)���*a���6z�.Etф@a��ɏ�M�����9���uk��	�_(���W�"��,uS�'�p�t�1��B=�e�LS�5�!��$2��Q�]��ȐA�8�aJg����f�+!��#F��gu;���!M8N����#\v�C���<:6��Vc��{��\9���	���:�>��8�>9.��X��ѿ�*�G�ӑs�=u?�����(
�
e:���N��.m���L�R�Ȳ�t�\��E@��B�D�U�Y���&i� �����7�#x�xz��:��zA�+-�s�q�aĬ�!˩?<*f�{���%���t𑘒RQ_sV�Kbjs�?�#��4�j��)ِ����.����]�׾q/su-��i�+6���Q5�y�k�B�)���Xp+P,%���������QZ��r��0�͖�-��f0��)/���4�*#�IM��64�h eJNM�?�����y�`�/�G/4����r����?���1Ψ�']{L��$3#���q2{���cJ׫������)G�8s��n]��A��{'��#u���/=�J�EP����%�@"���ݴ5�S�heX��'z�<3+���PcAf}�r�Y��;� Q(����Y��}��E�vb�h��, S��z����<c�"KT�I7��Q�	j�l��u�>�қ�pX�ԓ�ER�̐I�4�>?�F�.�G�X>�$\y��T��O�@��^�Fs=��+1$^��H^Ы�$4�3#0���O��Y;x.��z�nj�g";6�-0uS*c)�U�kt�?Z��U���+����I/�$/�0q���X5��u�ᶄ|h`c2���퇿cE[Iع���4ݨ�O�3'2s�'���aG������,q���Y]l+�J2�R2���&��m�ٺ/�:�,��<~i�tx�<��Nu�HE	���#��b}�uP�"F���Yw��U8	(x�t�(���I%��GwVqQ��ZZ�~2q��.o��l�*:����d���y
V{b�3t	f��f�9ݟ��?3Wxd�e��tGm�����Y�0�#��!�O[d+��`z(&�V���+"�L�����5�Ѽ���ړ����v� ~Fcώ���W�W@�oȿ����@�	��~sȤK 2O	L�9.�lEhaxWM�4�+��V�.�ž��S$��W*�~9�.?%!�̔�0;��L�6�T����t���a�Asl8+^��?<�P�]VL�?G-��7ߚV��`��i��������v�r_̵b�$�Yw[��x5�����	?�R௨�����s�mi��H�ĨL/���(;<�愋y7�v�����c�+G�����PO��������+�,es��|��5/���]P�,k�:��aK��� �M������}o5��ccF,�\��h�;.���N�)�+�	[���D?��8]�N�g�ᦡ4dd.[��
�u!�&���fxd��"��~Чy�?&�����I���ū:�T�|R&�e�$	߬$���Չ)��m���!Lv���\p�W��:�W�Q���ƀڵ�J~���E�FW�G�d�����a��4T��U}u9��J�ܧl��u|a���#3��pu�U��V�T^i����_`��l�@O�J�����ķD��C�6�:�Y�3�pͨ��z��A�����o_M����#�P�"2�99�j�!��uzg�ر�� #�C����>^�xH���9�������[F�
1�o��A�j���h�4���.tx��VX�h��Q�P���|,TҨ���g�����$wNy��t������P&%EL>�|6��+p��l��N9}�X��=�p&�����V��S,�>�6R3W|٭�-S[�d(�B��~�B��iE �n�`�/W42C���
��VXzT[�����a'�Ca�����*��sã2��pYP�58v9�w9Z-0N>���/�Ul����C(�zVb����%�����aciiG�N�ᯔ��d-UdΪ1�܊����Q���_�yKL�8���#�vfz�s�Ư��;qR-(��Ճ���
���Ձ�f���R%��[J�v��I�o��cƸ<�A��n���}45gt��q({<^���[6����UE|��eK�s��L��	,�������k�7�������Ls]�J���Y1�E��޼��X��k̛�}��C���ޔve�z�ʫ�K:eخ$R0=C�V'����9m�a,�i6=v�P��4�#>I�&�ʐh-�1����D?�)��յ �p�����_�vf8�mn pdH�"u�mC�f`6�r�g����I^[����Z�8��¥*�e�p�5k	��@芥��*���h�$�e�*�=P�e�N�|\�z�Z&B���ɗc "3�F�tp��Ü���K��&����Iq�!O0&&]��<8�`x�l&����G�.3�֠�4��C�<��O����'W�7��d�Q�؋�owt �u,J�<zW�:H���F��;�� �B��}Я!e���Ȳ���n�!-Se2�45��r5lIV�����[������������"��Y�+��?.n�3@��J��Հ/s��%�eS�q��K.��9����5zHu�,�����R�7�%(�V�[�{(>��y!�w�ԗW4�F�`�u�l}>�0e@�U�V�9vI�[��t��+��4��|�Ҧ�k��u��y)�r?lX�N���2�ڂ�kc�Â�� � ���,�q1������*א�Hv5m5���pO�k�R��T1���*y���~��t	�ƣ&.�'p��;�N�`K�ͦ�<���D�%�[�?.�?7��%�1� ko 95">JkЬ\��B����4Z�4�u� t�IA��Y��oAo|��W�e�?��ճs�>v)�'�����Ӷ3+j6֨���P�:�¸>�ACI2�H[vum%n��S�q������n�{]�vt�����6o)��0*{s���zh���Q�Y��f���'�gߥ���w���3�x����yq�}B���Y��-�g� Ȗi g�d]�V$���L��y2�x�<&�����;Y���K͕�����ݕ�|+��I���a�B=�Aa�C���!i
�� n���	(B�dW�t���FJXV�i��=�V�{��!,O��2�� ��{����,N)��ċ��#J�bN˒��	g����(Y�n�n�;z,?|��p�w��ө���yrl@�L	s}�a�
�����"�߃I��A=������]l� �|t�a8�h�3��)�t�@n�K���$(��r��#���Ṟ ���CG m�%zo��B��	�$�(ߍ��O���|r�HF4�t���e�}��Zz��zm�D�A�c�����H�o�n ������8���Q(��5!�e���[rrU�K\6��u�D��= v'���d�Ce1�1D�ć�qam�o�����o���̄�G��z
a�4V�!�zz�9�..��Z��ެ�)&��I���f��͚�Fp#��ͳ\���j(oM=�{A��u��1���&f�F���P���g�Eͧ�Z���Qg�K�'ʤI�ۇ&{��v�}AL�;v偛���kJH���Ⱦ9������iET�VLȧx�lFk���v>�l�7f_r��Y�~C7�kO���m�+��t)?���d>���\�Ȯ����V&��M}K��¤k��pJ}����"d*Ԙ�2�^cr�NMO�D��E�W� ��#;wb/�j,��a	FrP)F�X�8�J�S��H��m�?�=
��?!���o5�'1z��	>����8�0޼{堉a�]�MF�L �aXޘc	��u����xT2�.�NJ�Yf�ڲ=�L�E�Ͷ��}���`�&N�\߅���E��Ĵ��d�{�.��TY˄Ty_C�e�U��"�)�/��YL\�[eeĹk�ָ~\�y��z���R, ��xZ�M��c�3r�,��)\ѩ�UFy2xGU1�Y��-;]�U�ӎR��3SN��h��=c2�G�>I0
f{��}���`���F>G�
�_��R'\٫T�&�mʩ��˛:\DYk� � ����4wu���b;��V]B��afӁ��g�y���?�<euBVD���n�tԤډRX����Q��6VKpPt����0�؏�� ����81�fP�'�8恽������(�ޑq��I<���M2'�B
���I�"����{��0�S��z� j����:�G�K��Z���1耱�9BH����ɜ�quq(�UJL��D��6O�s�{���/�a� r�bJY6ͬP���-�q6qcE�c�1ڦ��mӣ0ʻ$m|y�\'�1��57��i��|��!4�	W ���ߧvGw��C)�KR�t����AP1�E��+m-��/���F;����~A��_�7���?��]���i�uo0i!��.C�r����Ѭ�r��4 ?喲�g-�D�� ��	��9�3HjV��+�֭�&���'�+^[ݜnҧ�������r�*G��%MDmR�����Џe����ACMh^�`U���y���5�:��a�L�^ݓ�j��q��N�:��0�Q02�*±���"���64��{�4P�ֱ��o�~%%��鄇"��_�5!�E�G�$LI$�IF�b��cO"wve��������ub��a�)gj��Es��0�g]�EEL�h;j���8�!&��9f5%eΏ�g����#PI�����$���p�-�h��U
Ȋ!P�p��O�3���+�J�V�K���|f��:��q8&��=WCW'�u�^7��&��h��U+�m�a��2ud{�8 ̰�<��a�r5�-c��r��'	��RΖ�Ҷ���N��S>ۦ_;�٘V�S�OJWޕ~J�C�Wz���9����,OL;�Ė�G��~e����?�7�+�:$1�
�\�{m ��I�.�i>��z�?���:�m~�"̅;�k�����J���u�{SiÒ�.��>$��W�	��1z-4��q>�,���E�����d�P�si��I���#Ր�;Q���jcv;�H�n;�[�x�cG��V�p��v�.��#�9O�zeh�0 �ʝLkj=C���N�d2���6(�O���ք��V#����+
u�/�&��l��j�'wyV)�t�tT��{��-��T���sE2{E�-k���,�_���MF�]�ܝ) �c�O���L�������uіҌ;+Og:|�W�8&y�$C����b%9,j� 	W�(T������U�>�'g)�cg�b�%�5G�Kx�%��WD��S�i=���q�����8�K��ETj��*R�x1��E�&V16��!��|ޏ"�,���/w*�˩���EY8VIo��^ރ����k����t&��:K�װe���({Z5�Z+����9X�	����,�ם�U0ѵ��l|<�&0t�$f�3�Z�
�O �͟�'O8Yl]}ަF���v|d�֦��6}}y���y"u;J�V��gdb����MӼJ�����i1���y<b"�1	�e^%�L�r�B�Η�' ��o��|������k)}��p��}����~#
3 j� �,����,�Hㄶu&Đ����w�l��:x����x��M8���|�Ӄ�����h�4e�G�)U�zc<����5W��'2��W���\��2�!�4��.��{sR�Aw�vY�H�D����D� ��N���e+�V)P4+Zƹ`ΚC���^�p���7�����6YY*���?��V﯆n���h���l���g�񤑪NY�f ̛Ԉ�.ܲ
��jC���>�RG^V�c����DC�v�#.N.�iJ�{���~Fñ?�8������&jW�3ΠR���va��Y8e�N�z*�ca_�ڠ9(���7u���b<a	�7$�����9$T���m�c:>e�:a "����u�	VK�J���+��e�X��a�PXa�%r_��zY�c���AJ��g̨p�f�X���y�

�����Xbl��k��Ƿo�zЛ��ߘ��/�`���1�?�"�i8)ʸ�lO�($�䀔�IE�E�x-ʡ%�B�]���h�D9Z�yG���ՄV�����xi���=)��e���F�������gs	/m�i ��O�<>eIٌ����$�.�?t�{ښ�W9T=�`ʺ�z�r����V�׸oQ�%�^�];�<
y��M]�P=!ל���PP�fd6@Q��m���p���d�$�.�����;�q��T0���b^��27y7��_�b4������ ��W�Ϻ�T�ά@�v�~�a�A�4�u��fGs~Ub�O9~ڹ�ZS
h{��U�p�5~�(�ZŚ
���$O��(cU,	0�K���q��qTPg4A�R�>�8�O
)E������Z�����o�ի�?��rۯ���j���F�U��R��U�T� �(+�n�~7z�!Vm�fd���*Q�!l6*�oh$��%��7�X��W���b�3�[ ��^:�s�e{@�����ry�Z�fl��|�E�H�w�[��_��\����IjQxl�F��R�mua��(}���e�C�	��(�$�c�Ae4�aڏ�������).a<��F4��:�=x�3�BA��2��m��c�fޯ�|�!|�2���=��IGc[�Ok�K�_jM�y�#*d\�]��]�j�j5�{]'�3�V ���sVoZC��O�ĵ�~���$��>v�4t�Ag�˻�,��xQ!טw^Ol�1�-'���>�DO���X���K�c8�
�[v��e+{j�C2��c}Q�"Ѯ1DUx�c[��lD���:H�K���X���u��П��l��\���O�=�5��R�#V��VGK`��	������B3�$|��p6,y��x���㯍�t�ξ�&�j1FV��k���;.Z꛵�zp�38=v	֯��`C�.Wt�_Z�oL������-�|�
�Y޳���S���y���D=�D���1�j}�02D>�
'�4QiBu��f�QJ�S�s����|r�e$-ױƅa�l���Lq2����a�xw�����d�/˵��J�z��٘{�E���Kp5p+��r���C��Z�����iۿ�@�!bCn<��>�U7g|Y��7�I��ay�W��ح�=���f�z;��M��c�O�a�t���=J�&��W�']Z~Lo�w4� �r�\�+�}�(wC%�_'P[1��a����fՉ�&gQ1;��m��^�_��wOsǞ
k����Q@x��%�A!E�,����c�!�ʕ'��c������+sz��"��CK�K+8YY����P��4���,l��Sr~!��G�?��`a,o<���֙��8���t�LH���~���������nAB٬D�����z�6le���cg-NK��Ա����z;��QC pEk��Jr������K�	\)�"�:342���؏��NL�V+5� �*�ϩ��58k*�����V�����m �]t��Ŗ��	�j�@�L>���^�.��%2��v�H>������H�2b��l���쩩�`.�5�^,��a�3�v}�Flb�
���k�ɮ��
�
:��n���Op���Es�;6�{o�UN��D�9�E���s��ީ�_�EJqnrF�7��4#�d�Z���[��
�>�0���D%�����~;r���dce��B0_"���,�ӄA�8��h$���
�b���Ovv'���&�5aK���|m�i%��\��n���U��6u��	!��_�DK��:����I��E�[<��xy��#zoDP�W���t�n��(��7���n�Q��Rz���7d��y��/�Ywjq�t2A6�5��R��Wvp�zr�Pt�֔�r"���Ʒͨ'��dJ�O����f�'0atoD����B����)��O_��M�STɊΓ�=�s^FF����+���p9MM�*�AC���_��ȧ����\Bv��wO����8�@#X��h��K�Uj�5d7��j�0Ѡw����\v6��������#�4[���?��"������R�"dG~3U딻�X&H[�p{$\+�m @&�����Y�ŶM�A�\���eX�N���dd�0I�ri��I�B��A�?7�\vg)��+�u����>�t
�r���Z@����>�pG�pЄGM���s����2*M'��kh�o,�D�b|�N��?\I@�>a��|j���
Հ�v�E\�p����!R���yz�Y�R�'+�%)�]������#�����R��^�^@)̾c�B!:27j޵�#0~�v����"���R;������T��r���':�ઐ�O�faR���t����������
^��ڊM��}��_דS��6��.4�h �9 �^Um�ϥ"�v.�P��5�bϤ+J���b!{nzy��J.����]5!v]��t1XJ�U�ӄ?_���l����`f��lj�/��i1vdݽ��W��xzh�;�́[���a��S����?�c���'=�E�~�E�Ĕ3��d9r�����~׋"��!;Cb�/`�@8(��q���
�n�0������"�����ql�UV����%@�55KX@��?5�����ɻ�V�
����˓*�J���
1+����X$�ۉOIb�ހW�#�0d1��g?@��ာi�H$H �8�%�--\��j>#���������D����!�����`5ǈ���q�諅oY��T2!E�����Ó���±Jq��h���Ce!3�sS2��S�y�a �>9=�җ��Qe��cV_�����fHP֘�͜${Q,]�C�R��,�G�~"T���(K��M��`�}.���Ġ�����1.O8t�K1yhb�ԉ-b���|����8}>q���CRL����`�uI?^Z��/*Ť`S��S2���	(��-��.�+��2~q��f�ׄ�A/��a<E+�HR�3C&��1F��v3�t�����jV�:�JI�	�2���ݠ!�'�ݬ��|�1�r?n��S�,����S����m��Ң�m�I��
"l�4˱s&[���n<�*���e�Lk͌'u�hr4
�,CIH�Z-u>��'�;l�p�%ɷ��0L�Y�z�&����ι���ݨ��Z��p�g�Q�_�9��w�u_X��ÝT��\��c���y��>�jJ_�Mn�I~�W/)�Z�Q6l���J!La�->&:���D��������3��h�|�5��f���fX=\��4Q��c%�˙���0�O�35�ɷ�Ӕ�0��|�}�� �&J��ԭ>s��R�8�t���P�BZ��hG��o`e�9K)�����p�@�`�b��~߈9R��}�9�"]Db&���u���j�𳉂��缫�Ͱ��mc�k&�5P�	Ѩ��,�i��0�D�L�]��d�\'��{� t��h����[5'�n����07�t�~q� �)�y��.5k'�q��U�Di��g�pI����N���t]�����C�?p?��v��63��>c���{O��I���ق!��] �	�s�� �$�t�5�����5�mB��l�jQ�ێn�8SL�P��޷n�8^�@��x�᧟(��X�D�P��g��
��٨�ͷ�Z�&�*�ͯ;
xU�t�!2�K�R�=i@�ѨU$m�x�m�+۳mC:�;N���T�T��T �۩�fp��Z����[#s"�W�-0��A��2�P�k� ��M��-[��B+,f�,���`ئ���ŀ�M�Nvz8����M��tz�����p�Z��9�3��$��$j�g���"rQ]|G���Y��(/Q����X�1��d��^&�.�b���gJ���g�۹��ܗ�Й"��IK��ĥf�E��q��j�߁!sMZ��>0%��-.�@����5��g
'��#�a�~��U�Ŗ#�>��9,42�4!|��mJm ���?�J{oÏs�m�d�>=ņ��c�󅉲am�bDJ�����)z��O	��Rk%+;u)T�y'3c�m&�B��M<qO���� x�
��RMTƊ!'��oQ�p