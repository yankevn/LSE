��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~��[2�q׵B*OW ��@�8���uG��.^���`:D���������EmQ9���@�&w�&��e�Z���,] ����r0g�c�����̳�<�hK���=��3ksXH��>�
�uخf��)��y�	���PF3X�4���8���5J��v�{%s �L�7e��_��:��7����(�>
�te�f�d��N+N�ȏ��y<���h�*U�Z����ꠝ��2����P�_��7�*�\U����=�ٗ��/6`��G̧�7�0��?�H��16y@lf�j��W�{C�ͪ����@�^��w�o�ҷ+�KoR9�(���f�gzY\��m���<@"�]-ܐN���|�-<
����BRE�3'llbsQ?E�A�Y�{��i(�����)��qD��t�	A�b&j���|����`�C
_�GW��v���N��$�5ܰ�p��{	3�c�$�:�A��a` �׈�n|��h�3<���ٔQ��g*�l��dWz �b�?��ޕmp�>{n���gۍ�hc�J�\.dR9f�x�Wa�@�"��~\3�+���k5��մl��ra>���i'�����j3���%%��?`�e�ڃ5?3�t(i(WI�Ͳ���@�@�{�i"��4S��6��.YJ�m�v�:,#�Y}x<�(r�=f��m������UJ�ҔZ�grad�b�<Ĺ�:M
�����Cɇ�hW>���&�Fˬ��'ޒ��p&
Т��D2!]_׸���0��T[G��&��a����@u�a��X��gKM�#��cU��J{�#M�K��St8K���g�mn���u��ٽ���z�sT�v���Ua�[8���֦�yW<J�뢊�S}���e��\E{�y�QtU� ڂ��!z�V�2�rJ�Ru���0����?��6��mD��;��#b�'շ�8��@�S�Y�05qx5���?X�vn��`=���l��BJ�n�^��D�:W��i�Ƹ�UY^�>�h]{/M\'��3�⛸�_.�I����Aʷb�uF�&B�{�솿7�tD�x#�9V�+/�!}�m�N�=�
�hL`h\b�rј�9'3~:�&�>�t[��<W�4���M I��u��_��r�����d\a��G �!ḥ��αl�4��.�d�g5��U�!����,3]��S��k�ҡmk9�`��q�����4xFڬ��m���Uh�lbL]Q,��˘.����
�P߾�R��ㄖc��ԝ�m�K�ێZ-~��KjOIC�+>���G ��oC�ڕ�%����Aǖ��̮v�$J��;��s|��fZ�,��]��o�:!�t������1ԑ�Wҵ�n�-�T`&㋙!@��f��.)ǵG@�8��9���6*�8��ZȦ��3{�[�Bs�o��}�݊@1X����.q}dh�dJ#�n� #"eh�Shr�Z�2�:`���咖�+��7=��Z��>IH��@�J@��	����#~y��""��'5����<@���9��������Y������h��۳9O��s5c��N��YB�"������4��;����Q��*"���Kв�K���P�o�&�Y�ho�44��3s�T��Z!�Q��a:�⋊дB��]I��~��]�~7�gײ�^Q3K�:�0�����MjE���/���7�H�����Y��c1j,.��O��%���E7����7B+�$�w�(��ƶ���W\���uñK�o
�\�g������ą��D�:3��D����\��lg�+�^�_�"7u�V����S��GQ@`��Lѫʧ�hTݙ���MV�(�������S�.�LA|B�����d��^lT�^�+��rn 	�z��V��*���J�����l �`�e�],<��:<�vג̯wX���%2�s���b�I\9J��/�w�{D�Ros-pŇ���-�]k��d&�Bꩍ��=�����ҫ�2���-�����]W̾D���wG���@��e��������7H=.0�6t~q����¬9��L�G9�6�v�yS��]�>�9>���VG�$��2LF�Y�s��c����h�#"�F�SD����ԑF
�D�8�.
�Om)Ά/�$�l�s��A	60ڶ��~@�H� :ѧ�(���N�~.,a~kdω7+Vj���Ȯ0�<�f���(�����e!/u�i�FS0�mrd#Xn��i���ݱ�륮=�����Q�^�U�I�}:��B ��$	79oV'0-��J>�����Df5��$Y|rG2��ݓl��X�^��O��}�[^R�h���c�O����Nb~}��n��� iÏt���4�1����Ց��P'^��;���H���w�L(�� ��
��j���H��1�ĩ*���s����z�V�}XE8�!���%b� Ͱ�r/�]��9yHוJpx(3��T����1�,�oJ$�Y�����v�}�T���+Z#�l���T�C��<���b�v �z�ޗS��N2��гkyhPA|[�lx�YI���u,J�RAu�|� ���� ���}.�
��ԉ��]�w�#˵[�)@�H�a;���7�H�|3&��r�n���L4<��?�k)`��\E]��E�ߢ�8o~V
����%���	.P��LЇ巅"�/�WA�*8[��KM�'u�h��#&���z-��E�:_�M^��R�^I'<�".���,����ڥiIļ���9�u��mE�p6ג���˲��Oxr����m��64��|��"�&ɴ̦�3��#��{�"a���S;ubesϟÇP�@M���/T�;���S���X;G�mÊ84x�{��*��j���@�|�B'M��t��+��$��k('v-�����|��-����|֤)1�%i|�G*iG�l����1|N�Vu��?�Ⱦ`�8�xt�q����אAjQzQ��GJ��7�D��)Dp��4�*�|tʇ���*���iB�c�]� 	�yJ�����PE�W�rB"��ܨ���8S5I���S�����>
�Ym]����G��?�-f�1Ul��0@M���؈�E��|��Y����"�O�*@���Y�./_6ׂ�Iv���@��G[���@DKW����CџS�ǟ�z�It���l�+aN��<L�Y-4x�ZW,T��\Χ��Ҝ���n4R���?���ڣ��OC������F��>�"a3|p�9�q._9��)��lK!��lBV��ͅ9J�H�z�}�r,��L}���>�u�n�Y5Alr�U+j����4J��Mq�{vb�U�DQ��Ža���tj�s��N��Hv��ǿ�19���Ң0��H<�ryQ��Y�i$r%�h�{s)[g�=Br�4�����C���®���b�?^��;�-�\	��e��*�>tjw��?jw3#<�L'*8o�����c��x6Xa�T�����wz�Sf�&�ҡ�(WW�#M5;��H�+QR��I��s�zN=�g7��~����S�'%jY��1_ ��ɇ� ;4���U~>S,��m4u]�ĝFT.�(�y�bz=DlTc�]��I��-,��\�������D����&����%�r`��|13�c0z�A�RA�н�!�760�R�b4`W�BMZ!TE*�בW}C��|5eI� �N��Yl:_@
^I�/���v��L�[,�`!E�9�{FFa��&r��������#iܨ�D*t������"�w�Ox�r:k��i|m��/�T�n�>(5D��?Tm!q�aI�>4;;Q
%�;j4&�,@Dx��<���k�x�\|�g���YqER/%]E��_7l�N1vlo����Id-:NF���57������9w��@n��}b��6�����']V�ﲴx����9{�]�(��g��s�E��ńN��P�n�aܰ\�3���%��Yj�y��_�d���s�bŝ�t�>L��O_�^���F�t���jCb�}4@;���D�@C{�G
�E�Ȩ����k;:!��f��9du����=yJ^{]�6��54�b�7���g]����7m�с�G��� �~�@xWoWA���-�h�������*��0��(�5�t��g�o�sqk���g �˗�i�A�DI�6i� �S{�c�H���m�3�^ y�`U�����:-�j�T�m��+_8�	uyĪ_�ǘ� !2�iP��n��z����QvW���3=����F!];.@�O�z<�{3����@U�B�M<�>��#�G5w'���.�N����{e�<0t�+Yv��+�@!E�%�j�s����ݰ�\�d���s���.��6@`�|�L�!er%xt�Y��(��2�h��$��h��pn��y�h�J��%�^���48�o��7����UN�M����^�L��6)�|<�0^l��ɚ��o�B/���0�L����YKe�N��
���9��f�N�Lٱ(�ty<�3��#�P���( ��m@ն,��k�P��P� V��b���'�z}v¦����(�̽���3(��xp���׏)׺�=�.��̌=���&�=pt��!�߼��Kzo�-��lVc�q���ֽX��AjY���K`��\��0��D͂�6T��z�C�K��In+�ACk��%�w�+�FO�D�En�zob�����<=�$4�_�33�Jy��W ��}��^�K�����]e;��E�DV���+�.��~X�n���/��#���C��ip�RǍ�һ�4Cɖ8��Ƴ��F��߹�.��k]�x&w���\,�ac�����C~�H�3 ^��6ic*��[$5����$�@^'�9�$����=�()k��	�}���^a��0���Xl����'���ɴ�=.�C~\���1E~_�:�5�{��o���׌�@�lF�X��>z��ɢ�h�6^��:_E�pI߽m9�m��[<��T���$2WSz
m�����u���1�a�w,�
�>�~��_H^[�Ƭ�g�sb�J!&ER���<�Bw*ґ�ꗚ�G�Ŗ,��nCXãr�N���DD#Z/П)�#��;(ԟ�^���'��j*L��H�l��������o�{�7����4��s�S}BE�OhC}9�6�u�̔l)��z�������nP�ԝ��@���i�2=�G��`M5�V2��2�Og���]�pBc�ؽ����ě��0� ~ Δo����������Y��Ki��'��-�qn0�ɟ��|�{~��	�-S�9���6%[LX�OV+Ϛr.���Go5*;��za�68� �S�j���H"ݙ{[.B�B�t�����!N��Θ~b��KVd0��3ޥ���l`>k���J�"��+��<Ou��L��d�<~�1�t�-���,-��@��Knq�s����-;^���O�l���7D�tݺ�?4Y�{�O��/w�ҹ���b�Z6d�T���0&��	�!��-
?h��(����3݉E���<�/ձ/�Q���(���{�$��b3(�]����,J���Sz�HƓa]½E9��S��a�R�O�����)�r�T�
�K91���&E���ſ�9�E`u"#�G�3����_�qz�%��Yq�
�2�]��P���X��X�4*%6��������.��u�֍���#��ff�_�(38�,��+����$�h�{qw\�5������8�:��b��3��!Ev�$��"3XJ�r *����\<JN�|"CW9�S���D���x��b�c$	#/uBE�2Fk��S��bҲX�@Z��Y��Q=f� d>{�e+��/9���iNyn���$ݜ~Oqd�u�`�A��a���ěD�+�CK��"������4����L�]�_���Pɶ�HZ����P��wY���Ɖ`���"��)\�o�|�����f �޹��k������9�ڡ��n?Af��� _���a1#j�\�h-�_��m�5�,�( 9��sB�$�u��P�-s:oH�N�߽4�`��كI؏$ߟ�Vꅚ�Lw�Ϙ
��d*�лB�u�bYa�xp ���ԻC�%�҂���Ζ���0ţ7`t�Ɔ�3��B��L��܄A�49���