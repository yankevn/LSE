��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S����)1�
��>���yOd9��_
�h�a6�y[q��lm���;�	�f|�	>U�ۗ�#��1�d���"")�˚��MmҠ���n�֙�a�b��<K<J����j�����.��/F�%Ix��7�#-�gG#��a�OP����zO^�1U��{�i�V�U�$�V��uʇ�~Ţ�%ehA;v�����=&V�Ə���c!��5�g��y�]o�)��ؒ�<C_ߊ���ZWP*�cC�i�Z#�_��/?�b	HS�{t�^��&ʽ��ne��a��7�s����Yި�-W(ϔ�OK�j��4���N�do_]n�H�?��x�@C�Y�(��.v�Eq��ryG��D��Z�f�,��R��zu!}��l@�Ɓ�-�;	�6��xN��#)�����k������b=��H,A��X�3�*M$u�"�ڎ�?[����$g��Z݉��v����f}�����5qh㑬�D�Y;��cNqU���k]݂uq�@��*��[p`�b`׌]�������\����}޵�I$:�0���#xޛ�i���#پ��Ǳ�-.�8�
e �f�(����^&'8�un��FF�1� ��U�,Jn��9?��n$�d$Y�}� ��� ��'����ElU���P�:��ux�6�U��*ݎlz:�[
�G7_nE�+�r�H�\ҍY7��~���}����"���z$�t� W5��T8��&����p,���FXݿ�#O�s����H}�]��!K||��(Z~��F�jPm�d��W>�:��P��=�o�;����<ǔ��+�~B(��z�4�=y!�'�-�2���wm1�����פ��?(�|K�����)�����R���|˨r1�џX)��W�!�+��߼�K{I$C��q���ZEq�����` 3�9y�Íǧ�LR�o���D��n
���l���Z2���ܪT}	��@�Z�e��*s�i� T�rkN�7g�W #�ӯ�`qR��1K;���5},!Sz̋^`�}�&p�VqA��;����Ü�KYh��Q�8��$�|�ٓoj��,��&�>`/�yc�	��n�3�>�p�K0����[�~�
#"��Lȱ"ie]<�����QJ���Ě&��s�� �G�~�>C�}x�K�:◒opY�Gr�&'3�z>������I�N.k_}\�����1-��t�M�;0�V�e�����d�f��GYԍ^\�WT�[(�Ni��)��M,n;$˓�Ip���� #��ʖ�$>����mp�oF�n�Ѵ���y�Ӳώᡁ��Іڢ�ؚ��<1e��脞KZ?���~(��\<ȼs�$,�ٙ�1�_�l!��B6��=v���M���YJ"������&�5�_R�u>_R��k]���b<�u�g���G�؟����~G�܇�T�,?
Aetb��l䕆d9�-��H[uK�d��8/�Sܠ�c+�L�#��>��E_�����?Ҥ��nSgMϼ�(�-�Su���gk'OP��@7M�[�I�����j�{��H٢�
1��v������cPp��7�ko6^��	��E��k>��dh�#��?5�]AjU����5	_J�d�N 乪�YW�2���Gǉ�? ��Divj,1��h��(���U��<��ҍ�u6��B�"�h�AV�� �x��=�)�e�2m�%�MZ� �'����?)J��s�)��Ωy[yYKv���*>pCc�Mgp�hw}"W��Aʴzok�f�p�Zጥ�pU@�F����s�\�ta���,|�<�w�/�79^�>G�X����w�^U�g&Yc�]��u�$Z�
a7yj!]�M��n�y��k��\�j����^k�ɵ���*��[ύh�1�k3��J�^��\���Xއڮ��G�0{�p�9f$0���$Ei9����e����Zj�k�Ҫ5>��$L#V�>Ņ^��q�X����M��&tE��LY���rx���PV���7�E�_��*�6�(4�S��-F��&��j�V�3��it��k��iPZ��S�'���B���#�a�d�d��wX.�[��`��H�%��3��!<���|���2��6O���NAh� xҍ!q��`�#&�yuQTԉvT'��������un�т}a�`i?&eu	�]A�������|�����L��A����=[mS�QwX����������=^�(2׹�V�ޑ��9&$��3Fg��5�����K-�c��Ϗ��{m�}Z&9ߘ���~p8�<OK��d�Z�ae����,I@l�Fc�A����Д�ts@!V(]����S(��w������Q�Z+��":[���|�� u��f>']��ͤ��hp����5�S�\�O��=Z��n�S�"-����ªR8P��!�z��_j���k��J]
ˊɯ|}� s4�+[�e��5楗c������Iq`p����{P�a���3����M�����+*���-���\������T��;�(��Q��-�'�)4LL��*�0� M1���T>|�u��,-(������	��PCb�dT�3ȓi'�(h�����)ޤ%EnMSs�Oqɗ�YF��bzy:��y�i�f�co�\�L�&9A�J ܫ�ǓL[��U�e�7/Q�^r����VG�ڍ��*iE�wF�:��쌺ٌ�^�Ǒ����3:P�� ��Չ\Ϣ�>]X��ל���0�k
(�U���%�{:nA3��h\�uM�1�R�;s��8��-n�gc��3������b�$"i�Fw�WX�C�{�v��o9(��NU�9YVx4����9=�%L 4j��v�pBC|KR%���Z9kH�Xk������Q�x-��|\�G�L��=�u��a�Vc�*��9l��#DQ�E�8�T�M���*� ٰs�|dN&&���������cxT�&_sNnM�xI$ ��C,��v�#S�/U~�� 8꯲���c#��^���|y��R"ށ�#��Q����D���b�ո���M��ʧ0D+�ȥ��A�j��;^#��0H� .T�iiE��ߟ,))u�=��s�qL	�:�A;�T�?׆��u�^��Ol^��qa2�"<c](.*�z�L��.������E�b?hZR�y�&��R�����%j�ꁈlm6T
؂�{�Ag�)�C�x�j�b�?�R^����}�[3�==΅��^ �늠��)	�)G�l��P]�6eO%n̒!�GR����>�X�;5����Q�?���l�p�d��D�z�̃s|:�7/6��d+��=�}�AI9so����\�����OcӨ"�_1�/-}��K��H̲
�TY�O�:�(p~���H�o�������~��"d�ϡ�]A Ѯ r������[jD����!Lǻ)���(����͈yEt6~F	_� �K�	Q}R&ڛOKB	Ћ�A�*2�]+�XA�#�|�43y�����w\�`���]Ƌ4�s��㪬���V��Q.�TZ*�װ�s�>������"�PR������F�}O��|��ɯ��I`a?^<zGX��Uƥ01�f���	��:J]p�k�J�	����Ѵ(�|Z��d�N��7ƣ���;�V�x��a����=#m�a�����gF�8��|�nnяT �K}��_��D��@w���k��#9�)�꤯�5J�{�,tm���A����﹡��l�������l�<�	b#t�ik�H�@��'��֛�DJT�M��(Ü�`�t
�v�Χ��T��<�[A�k����ȅV�9��%ĽY��,�V!2>g�\���+/���_�g�Q�&��`�vt�<�qO��s+��C����)�mQ��̬��<���x�w����4r��v2S��+=��;�*U��I
�op9�ڶ术ɄG=%�^��1o�S�N�3�Ӌ���U�t�"N���*�J����?
�!.��8e�/6n�|�4��S���0���?9�}�َؘ�N4��,�^��ǭ쇤r��l�o-l��5h��iۣd�Q�E�n���!�	���@��I�+s�F�nL����˔s�8yKĢ��9����
d	���0�,��'P�[���-�v����)a.� ��]h����@��'кE�k/a݊/���K�4�wS9��� �ſ�6�j��e[<�[�w�h��	�L�0_ ����u<��ө�e�S���Tiė��%��)�������ɪ<HY�m�����A:�����2^�cyeD_���.E����ܓ��ڕo2>:��+��O~�^G�<=���b��3��X��E�E�K�m��ǥV(ia�*<\.7ڙ�x�,n�B���7�!{����`2b������4�"J�h:���Hj��~�4�1���i	�r=�(�&y�6_�\�&�!��Chi{�I��Ȩ����w�5E�e_I�z%�c⨴�I=R���M�{�P+���k�'���KI���W�X
�jF�=,�J{Ny_F���J�~	�9]����i+_������q�r��c��
n�S�����x^Ƅ˥���,�>P�����	Ȅ�pʶ.�0�3}���u*��'������_a`����	Ϛ�^Ij!�����&�R���ҫk�p�k~�@ԌEl��� co���~z�5OUȰ�F^Ή�C��mm��ɧ�R\Ėg�Hu�qM��b�{v���R�h͉d��Om���ێ����E�Y�DG�J*�^���Ft���O�/e�8�S�|�P�S�d�ѿ�6Q7��y`).8���:��=��[d�l��jZ
��)�L�kt3�,�|�}!	ן̍���h�m�q��ǯ�����=T�cL��8�#��m��#�}^�)��̴�����(|�1܆��M���H��0��hHį�if�A�Ce�n�|�#�'5>w��]���|-�a�<�GQ������>)��J���.�AzBe����4�2�5h4?��Th'��&]X�v��E��y�̩}g�8�Bq�8�իm8S�Tf7���نI�%wis1��}���c>�'�h�j㮳P��>v�g�,U#c�QB�b@d�.�hq�x����)��@V���J��̿s�L� 8�o0W����O�z|���)&/m�����X�煿hi�]{U�� F�q�����/9�Di�9Bj����S1 �m��