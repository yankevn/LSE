��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*�G�	3�`�{��G�W��;�
ֳC�?h��_���=�o��n�(�
b}?'Ǯjք�_Z�ϵu0f���Y�q[�m1�pp����&%�a��|:ꃸ���)�5�N��4k�, ���o�p��Z�c>���H��]At�$YX}�+��lj��^�E/��7c�1�Z~�$�ף�P�7���Lg]g"�θ��>`A�$v�.)�0(l�q\���i�es����,����e�� ��c�Dk5��̩�t��z%���"bD��p��Yރ�Ҧ���B���۾�?�У>Т��x_·|����մ���V),8F�g���otp�,��V]�d���J���6�`Lk�n���,q/z":��!Ь]������u��ف����R<p�3�[�my��o"F���/�Ӡ�+�G��]w�\_�+Јw�Y��DCn�4��&tO6C�2D���`8��r��tEH�#�??4��#S�S��w0N�B[Ht�N�0��V`���(�yV$?V^�r��ܖ-��Ս��&�X!�]����^^��B-}����^�؀�2	_�9��6@u�W�;112��6Mɻ�\��>w�B�i|�꣩���g���E���7	î)�Vb��l�t��
z�1R�N�P)C���T�G�D�u7Ŗuic�	A���Sޘ�Z�j�v���T�pc,H����A[%x��.K0��1��/hfCبb��>�5��"]�����������`��w��9��W�����,�ތ������`��Z��"3*d��n:�"uѷR��+��������BP���xl�&Єϼ�G�I(���X�X@�b�c�;$y�O�""Mˀ��'%���G��;`�ʦJ���!`@�d�e�.�:�ڗt�Rx�mvL7|'��d����Q�ЯTΊ&�lf����/�;C�Oߋ��0M�G�f}Ms���%W8�TJ��qG�7�yp�x�m}����Ʃ)�#��2��g��)����L{W�˩���z�����Gu/t�L=�����7%��qQ)ڈˢҕ4l!�M<�^�m&ǵm�۵��<-�.�&Q�[ϛ�O2���DF\��X�&���⌙� �,�@��}�ڥ�����&Q`���R�c'��u
L[�A���W8����S�>J���,b1!6V��V��]?U0	k���	l�D5A%Oj�拼V�5~5��s��ƺ�_�,Av��U��2�3�CC��I��J��~{�:+�QK��xM�|��,����D�1��*��Y����2�^r-�p��!*���A0�d`��n�i:J���{�������X��[�P�M��cW�$ñj.�#�Ir[�����2�Y4��*e�E�{�Y]S����Re�L�>w�
�0#n���Ky>��*�M�\wN��擴M!�͓�j��g�o�ǯLc�-�'��d&�E�]e�_ ��pJ���䯴yw��~�?�CY#���,�tݗ����l�b	΍�l����%��S����7�[m%���xZH�Q�����vmU;��kύ�g��D�'���a�-O`%_ʬ�N7�
���F�[)Y~쏥�pP���ܷ�nX�z�
����}E�I�X8�C,��Q�(t�Ѥ�95�"f����4$F�.
�܎~"��>>\Dޒ�EM5Zs`�k͓��v 2$���ڒM0�SZ��o�Y��u@������o #?uz�N�a2�O��QJ���F�lo��~9_mC�%>Y��,�����x�S$��I�B��"p����7�X��^dJp{�<:!-�Fy�wo!�����(��I=����:�W�y=
�g�h�����H��Z�a��
��L�ݓ��L�?(��x�Wm����A~�4����l�Z׻�DS���밠*�#c ������ps�y���T}���"�4�b���=��Ӛh����S*@��@?Qz�x�m�	=V�ڛ~q�,�31Pj�������l!]��h�o.^�	�E[)�d���^p���c�U��� �V�I�1��/��o�C�B:d�^9� ���-n���Shě���f^Rg�P��F4UМ����d��$��3sQ��{o�M�|L��/QN�]׉���Z�tܦ�[(��u�@V/Ҿ��ޑ e\KJ/u��69>�ͧ=�Uu�ME��ds��?]�D�o@�L�E�����J�d��
̘�hPSlz�`�lcoة��cr�� �AG��(��� g��/�ש��2�W���o���;#�^r9H�[��B�0N�li��+�ߢD:?P�dwiӖ�4�"�T7�f�Uңb��^:�i�=c���#�E�T�*<`�C�}g��8	�L�#��)�����<Yߵ�!������M+G�5u���¿�)��{ַ�Фq�ʡq1������^�v�|Ch'�؈i�H8e��O�@�2�����W#��?�r�"�h�W^��C;�l羃L�ޒ90U�,i.:���{���&���7�%A͞�'��i���v�����e�e�R]<7i� �r�Z _;�Q-�����^w�1���ț��&!��+Hc����O"o�1�^>A*<�b@m��y90B�r�-�#�@���g����w\����Cx�f�8�F�S�Yݸ7� ���e�;!&���M�P��da��E�Q��1F^P7<�^%���G\�9pAn������R�T������>1�-Q%��z9���]X���e�E���]�Nk�� *[�(�;�&�����-��7�$��6o����O|d�>�
mt�:���_V�!)2���x���&�D�˿���+��Β��/�ل9�^X�Gce�}.��c�R���L6bf����r�N��l�Wu�`L��5d-:7)�mG�����ψ��n�r���!gP5#��&<_H���������y�#&��*H��k�.����jI!|iD>���q�㒳����C�n���nR�8 �����5吝�~�[-93�]��$���^���(jY�xE�4Qq�ƥzxQ�?ڰD�e�|�EK^Ob�l%��Y�7��-��w�T��I��&����p`��7�dШ��Hh2�.�����i�+:u%J��db��P��oO��lN�g��V�;�a���>^��6�.4B"��{����w~l^p�K�4]���۷7u�KZ4@�j���n#�Mi;��Q�߮���%��Lz�������_ã�d��k�-��)��1Z%�����RA�<W��|T߱@Z��p�W���º���kBGs!9'�i�����"�N���&w�4�I��@"�\�g*r���ǽw��!MD,Q�����IV���"�\(,�������zz��I���ώ&0&�a^�h/�A��x_��D^�G�������:�}; �R�{��G���
��6��l%JC3� ��c�H����7���?w�ܖ�(<ʲ�t��M���S�d	*ZD;��'�/k�����ٺKc� �2�����hָ�&�7�������ik�n7�Iѝ��F���N�T�`��&LZL�ı���$`Frg��Lʃb1E��o�?r]!�`>:㐅=��q��~'6�-�s�T�զ��:�P��Q�T�F� bz��O��9k���Z�����S�o��`��G��a8B��X�b��[���)�2�i�tWV��(F�ɹIm⺫c&�|A5��٫LE�p)!�����f0sD�O+/m@�R���=E�Qp�5�Ԟ��P�8"�^�o�~��d㜾�<�T�L�B���5+���p��C�6{�J�$�.���-��,~�3��53#�ld!�l9��ޔ�3�F�Ƣ-i=�"�Qp�9��I��{Q���$�.�/q�[>���/*U p;�4�!L�3må�S+�o\#p%a��)g�c[�0C�K���7�j$�7�vF �^�j^]�Z���4���ۮ�XU
�@�D�\�5��o#�W���L�NZ�=U䦓oP�U��c�㗋���R��W���62� *��	��O�1�T��������� t�u�Q��sE>~w�Q���źAn&9�������#�%&i2���٭�����͟�"��みQ?l���,�R��U�O�x��+s�S�݈�4�+&8鎫���*qV��ה<�5���im@t�U����}f �a|J	��D}���x��{��~�iM�u�CK����'~i5�"��0YWT����`inĵ��R��I����2�܈��a���'��Y� �?��^��e;��T�ݢd䛺���I6���h�('e���sT�;t���=�3�_+l�*7z��#�7_O�>���W�������$��9�}ҕ�$q1���. 1��>tg��27ņ�<f�����31�:�q�2 �?����[�ՅQ���І��@jP�N�Ӎ�u	����ѡ^���E��O�T��O�nv���+���6�FmFS�t1xv'EՍJ8���ѫr����[S�m�\�i�W=A��2���]&��l7ȿ��/i���I��h��^}�JbfU��'	����]�_���F@B��Lic��t�$��e�f�
�o��2T�J?�� ������X~��}m��^��]��M�}���U�����C��rl)�V-?!���`�[����	��O�����0���n����,V������bώ3xǯ��
TbF��pov�)"���ٻz�T�+�|���̷��b���ZL�5i����aذ?l��#����1t{"�(uݧ�A=�(�D�2	;�,�� ���Z?�k�|�/D v�TRi�rT��29�yN���%��9I�[�l2S��d�+:1�rU�%8�mk
0�fY����ʑ�%��Y�̣u=�N�E����
o�P�k�YQWl�1����ȴt�H���X��B t3�%=�y%, (�i6 ,u�Ē�S���"��"gsS/��m���ߋ�G��O�~�N pGJYpBrw�=�ȪT���˧�°���E�s�g&���F�ү�7��jzHk2���!�&HmYOF.�I	�x����/�!C�I�K���� �D����U=5U�"8�mud�]=f���@b0�K+q){�,ԉ�c�
�^����C T���������)�^��F�}�q.����SK��5�X 
����҄����Ɯ����/���E(��1���i-`���	a+�U<�o�<;�/`�$Τ@Q?v���5l�%� Z=^�%i����r���ye��"��&��8@]2X+կ��t�A����ARddo��W*pth5�x�������!��� {CN7Ck/�b��h�ң�
�:p|�"�,x{�6��� �aN�w/��s���.��� .F���v�{*�Y�B��+}l��t|���΋*��j��8��Y�����8�&�~��+����t�2Y��@Yq�E>�z&~�ʅ,2���=5���(X/ȁ��N���=X�E�m���י''��מj6E'{�]=ԝ��>�CP��Ss�Ly�^�x;~�r����Cv��u�v5p>3-�UZ�Ҧ���m��Kȵ������n��kr#ǒZl̊n�F(�^~�����G˾{P�����f�UG��4'sˮQ��9+=ds<L�?�Y_��8G%G ���bMpIr��|��2B��DZ~�� ���E�ä��X�q�x�XGA�{wM�)����-*��8$Q��P��0����Q�*������h������
�]�`�T���5�T�b����7�g���K`��4�Ķݼ,s��N7T������F+�HI#�@&�a�u�H�S+��{Y۔�Kgѵ�S���`�&��	Z���/����+��!Cu�����\�ixP�B��.|�g�I��I��x9u�����ښ�M���>��8�[�4&��yYK���#q�)pj?h-LJ�!��.�Ep�!��>hщ�c	�4N�Ln��ǅ�:�d8@ΔZq��5��/��J���1r_�ʓG<O��N��_qs���Aw߹�oT�晧르̆�Q���\>Ң��r�]��3�K9������چ-�f��kC+0%�����QF�PR��'6!E�-?�0�&!� 8C{� V�&|�~�mh�Gc�3$���p�	L/����*:���Z�|�j�4�,���=�G,I�k��*�A��O��D~�ڽ����9Le\�{`w�;��V�Ӗ.䟒�8�����R~:b�Nw3��Bm�We��Aȕ��g+P��������L�Y�~���,{53q����93h�䷱�#i#B`�W�]bYqX�ur��}��9.e��%��D�4$���h �?%x�z���"�z�vϦ�BRM����h���JP���<���	0�qA��Q3e���C�_c`-Z�eC�K$0�-�A\���Y�!R��~F��>b��8�D�O�M��]}�Y��ٰ[�d'H3����m�΄�&�d�0��_땨W-��i�x�=�!�&;�p��=�Vq��3�S��6�I:��%.�g���g-Kb��|ж8dǧ�H>rh��.�ͨ]���$"e�8��z�0�'��pE��;C�>J�AP@c��<��f]�s"C�wR�bd�ᅷ���?rsg�-�=r�v��5�u��ͤ�T�� �*�pZ܉������>㨗����&*�1च&���1���o�1�ϝ>�7/��%���5�Y�<��%cѵ6/�o�43:.Y�ǥQkV�zζ��-���3ִCBo-��f��r0\�H�_-4D{���ˣ�P�
H
���� ���i8���S�d�5����=�Y�kk���tƝ�k�d��<l���݅^V_���o�b�X���|a�vꕸC��u�2�T@�= ��*p�wt�\�,\�������%�O��ǖз������_���@,.�/��qL|��"�MrX�J�C��YiU�I�4�=�X@^L�%y�T�4Qa�$sLp�Y����2p�-/��S��8(9'��2N�|(��G�n\ٸSKb��E:ٕ�"��D���	�Þ"���hC���Ӟ�+)�Y�H�@1�k��1��	y�������N%^Bf�gƭ���W��f�
�RN�/^���-���Żn�UqY,F��'&�!�n䵧q�|Ɗ��K�����a��4��j�t��7�_�9PCe~;�l�=����A��>�8�Ƽ���,���C̦t6K�/�k\6�)+��eae�j�&�VH\Þ��+G*�먞d��t5�5 ����x�{�S��j��7b�/�`e8'3�J�I��
;����������W4�+�r�������%٤��lY�w,��Cq-Eױ�Kp�Wc1��c�c��7�Յ��3��G�=s�HQ�Gc_�����H�[a�<i�.,���gnZYa��̜��|źr�,�����1��Xs�/�T߅yI���fS��b;�H.�������!�xE�5U2&U�͟�r�u�^��sQ`h�Ő4I%�?����Ygjg��C�;�5�Z�S�U��Q^%�R����.���10a��P"YgAm0�@�ޏ� [}��g��X �]4�)������K�3(r<��fy�g�þ>��zc0�Q�2k���x��H�8���r�_W����k5��1a/ 3p���geo��n�����Ʃ�ܢ蓪x-��o�ڬ>���+�</wş��e�<�0=m���\+���������S�Fn8�}��C$Ei jɷ?7{�N�1F{�l���#�['Yh�F�7���ީ^ 6 �ww-v����D��2�#:(�o���R ^o��FRR�6�Z���v�#� otv���"N`������H&����f	�^1���1'����Vy�E���N(%Ke6�:3gM���:�}PyY��ɴ�c*����{�H���\�τ�m���	y�M��.b�E;�Y�4#wY�]fB\5����R���vW�m$�o���
�)r�N۟��r[���M��R��wls���
˲������¸��PH�Í&�c�sr��E����"P��=ϲɰ	���1	��߳���Pb�2K�@� /���d�L��r��3%ɑ�( �|����#X�"c�%u�tB_��8zd��R:.\�u�o�5.�a���GR_�/��*��Y���@=�u"GDPM�E9K�ð����Qx���aX��	A~ɚ�i�Ɯ���ru]�X�ѩ8�*��Ec'�L�r�C��e6��qc�s���Z��l��Vۇ�/�3�b�k�13X~	��+# |(d}E� ����%�QE����
�H�ڌԇR��T�
�wN���r�h QK��"��W⬹̀�r���}��'�/�K{��s.�Xc���q�0�ϽO~�븂������y��i��lŵR�	��C�}zW��~ĉƞ��
D=V!|Q䯦��m���r%Y��i�Y�%��s�I�����3a�Yx������"kM��L`�}R�8>�W^��N���)8�@pq8�@��/�2��`���vT4�}�K���ן�lb7���·���AHV#�WUyY�&�g�����������ɭi�}���������[�d�}d���n!Uy�b-��d��+�(_���l�����������z�r	6rS�Fw���<�.��,1�L�s�@��ͱK���%�[�hL��/x����cG����-<8��Z��+�U�9x.�͑���--I��}����	h��8e���X'�bH��r�Q��	���nj�<�����N#@��7����� ���x�t<zj_
��p���
�./�P e��{�@|(��'��.��c�x���Yz�Jh�� |qEDy�H���o"%��q�o��Dlc���m<�X:�S�)��M���L��c䧔k����u ��'ք�V�94��ߩQh��XĹ�=ee�/0�b�a}��3��i�:'�s$O����(�%��7�e�2/�#Gڱ�%���c�8�|j�4^Ͽ�+.����a[�~��C�[j46l.	�K��
>�CZ�俖h]���	8�|,#"x���>�lUx��fǄ�69n����^����c�ߪ�2�s^�J�S]���>9�%h
�Q�U?Ny��bQk��S���*1�3��,S�p����IG�ba�[Ci\R(A�!���_	�;�r:���B�d��ɟ��A�}J��t>	+�l@�r������N����S:��#u�M���\z��K��ā�d�S���tvr��W�ϙ�����2�\>e;�� �5�t�N����\�DD�:C��?��0�*$�����T�>�5�\sM<����#����(�A��Q!�*�{3�]&}�ɍf��>!kO�ԯ�d���� � �3��gf�M�ҬoIS�p,�ڵ$FV���$I��D�M%�CI��ǀ}kD-��qۣ:\io�9��vJ�����-�*x䑙[ �����00�t�TFR[�$��P_*�K����W�9�T@g��P�v���e������T�i�-S!�8")�"�or�!P#k������)�o�Quf+����t0��e	I�X\W!p$�M� (����K�N�覺 .�A��g}�����f1�:���M:����N�e�@�"���S��۬W�<��h�d�\�%Y=���bqO�*����*Y��$!�5�Q�=@�f5�)�����Gl��QP�b.c�k���^�G@��G��[<��0�5|+g�M�$�D���˯���u\�#�r|oO���	�X���	��s�Ck��8jd�-m?vK��jO����}1q%umj�r ���\s��>��5��e���t8�@)��-D��*�LL{j���y,����o�Vo!���3�NBt�zV��g����+��ce��4U�߹��X҄A�{����a]R�9y�aTK�˛Y�ƘP�:�H4�޿#��2v{��`klh9z~>�����=	
�U�mڢ)R�T�}6&n
:f)$�!lR��o++�6`��B�����r����ZIݺ��C�%�Э��5��Ǯ���z��4留V�ٴ���[�0͛��Ld8�=q_	�C���[T�������6�����,V��鍿���J�B���&i�h/6`�6���D��y@^Yo*&�T�w��*�)�E��g�ao��|�#n��ִ8��(�e��v~ѱ̏y���K��J�i\H�&����=�$�*����$)Z�J�*�9x�\�p2�R�&���Tx�G�#�J�j�~��=��^K�9�u@J
�n�4�ܾ&��"�PJ�va�?�-y��/E��e�g'�@�$T(}O ����^�F���H�X�^�R�n�,�'z�/y��_n�-μbLI�p��D�G���?ځS��TRS����دV'0��n�0'=���d�	!W���9�4𮈧-3����Ji��3�\�R�B��Dg2jp'�bJ�`�,!ww�ki�]@��3���x�[{���t�S��Mr�y^�~0���%�,j@�0U
̤ϓ&����)�n+��M `��F�2�ƞ�p�����q�α���/u��V�l6V�"d�zw(SO��C��p�6�]"/W��0�,�����n���S\��d��c�_}�w�04j���ԇ3�^��L�O���O�}��&���_�F� �v��(驓ܲ�]��S��cf��Ģ6JW&����T-�]�8Ƅ��� �=�^�.���1�&��	b��s�quY�
�2���o.���!O#Ǳ\�$�k/��#��{\��~�%Y��@��OBf9��NJ���T�	��������h��z��Nx�x"�s[�Ѻl0�v��qF�YU	����=�KK��ѥZd���4���3
���ώ4���ǂ��m�x�e�H��"b��I�.�/�S\�?�fB���]�ûl�Su��fG�fK����}h��Т}<����F$�Z�V���t�J�r�bA(��^c���&ߙ�t���5}����T"YV���r)q��sj��4�ʢ�yT���r)4��#mR��-����;�YR����Y�b#��'�ߡ�����7��!�^e�{T��VĽؐ��;M�X/�6=��;������W藧�ݷr��W�vK���tًq q�[qR\�&�?���\�{�c;M�[���\�kmd>R�k��b�9l-ǸtQ�M��c�@z:_T~�ES�
�`N��X/�Ǹʇ��5�e�:�P�Wm������S��dE}�7$X�$�h�K��g�(�m�ޭ�s*�%O�'�ϥ+A�߰^�K�u} ��YX�K~S���7��� ��z;�Ha7m&��<CR�����.n���e����y�e�Jj�!�����ms`RF�a~����ו'����ӯ��@ �bPFx��{���n��;a�1W��@�O1��'�0'Z�!�;��zl%:�ew��_��c	}6�Q��~�̻N8[����j�sʹj퉂ѫҊ�r,�ޟ�S����p����<�;�����O�}2y��t����HK��9�Eh�����i`gd.��1�*e��uH^R~���ȘŚI�<qdE�gz�5+��8��ʞ�Xf��ޢn;Qb�	������Ir�,x��ݢ�zv�8�(|���osYHQ���M�W_\���~�<SΒ� O�]���"�E=)�e�ku�ՙ���]����o���ZX��ᨔ�@��Q�?@�ٹu�dR��l�'
\��pS�3 �@e0��9 ��VNu�%����q;���x{���[I�2��|��>��k7�Y\�� :��Z~�����%!b'Q d���S�q�A:��
'�LeJ��!O�%���e��&�� 4y� ��G54h䊢B���<�U�!���]ld�-�@���e�i�G���v�L�=�E�V��Vw�oQ�&17%���ť������!�D�^N ���gf7��({^?J��>��s'��d~6�������Ե�l/�i��P)��8@��^ie�������{�[{�`Y1 G�Xt��oI�Y92�ɥ���9�� 9�^ �MQJ�$L07l��@�T�i��X��-"q.�)�t*-Jđ�8m9@y����ń�C"+�zQ?0�|m�Z�	��0�����X6P��:�܂� �[p�;��:[K{�8���D9n?��{=d�X�>���������Z���4Q��g8�O#�����B�Х�O*�]d'q�F���a[A��M34zZS	1�xq��m�_��`��Zݽ�׸�B>f�&�{�O�1u��W�@�-Z����W 6&3�&_6�Ε�5������;�P�{\y�������ѽ�3�!ґ�w��CE5�����kf�ʵ��#xt�
�P�v����>��퉃6���s=C�YO�l��f(�y2�d�k�L芕�Bv�ËZ�a��a���g�����Q� 擂gm�Ua5ټRe�T�Y���.����.͙�h���:�3zG�_�b�%k�����`��S,��:�K񙄜�(�?�@��N=amMen!��_����1(�u(UsZ
�W&�h4�'��F��;��0y��/1E�> ���T菵KE(�
�����[��]��9˞B�*P(3E���&���<��n�I-�,��<+^�JUʭm�D_�����!4�r�ߍ��K�á
n/�Bњ��!8;X�������x����{\��& �r���
��/A[�50��K��+�gS����������k��Qbл�T8�0�����ȂǓX>%���,�e��)��a�l���f���{����N���<�3x٦].ɲ�RWc���}�3���0�&^�LT��{���L�G��[�#��m���]F(\(.E<	.!��\y=�G5�x��������.*��=u0p
�����g�n��L=!�{Ua�O/���h]�����`���D�^_H&E��j��z`|v[U$@�xG×:�Y�+�̣XK�}��FUr]��d�L��
#���x����~��N �7��ڮt��:4������ͷ�Nʴ��M��Rԗ^�n���0�bp�i�9H)fӘ�머���tè�����@�v�ƅ֢tF�~ژkb�[B?�9��w�8�b� ��/6��������\�*E���p��#�f,,� ��Up
���%���j�q�W���<��9�e��"�\�&k ,�_	%-��A�zӭ,ۺsR{�8?jV�F���%d@7?�(�����EZ[k��7�hn�%�5K����o��Ƹ�OB��"M��B��/�A��ߔMىMRu�LU��"������\���x\��P����<���9�+{?��
�`�$�kRĚ]�N.r�o�:�7�������'>�_�C�g�͊�xAi>�*d��:�!�����d^�f7��~�ë�'A�V��wB'�tՒ���HK)l�����C�V�ʵ�Y���p �Iڬ����5�Qv���6�fx�����,z���ā��{1��8*�\�fb�|2��G4����D0��������X�e-��H�C���v �O��3��i�H:*���Zy�;K!��d7�+v�/U8����<	|�g���J(�'��?���Pֹ��iN`m�l���c�b�� �����*�4�M��*���0����-�P�h ��|� �ʫ��&�[����4� ��C��V�HO}����,C�ّ���iu�~D��7�w�Z��
\���'>"��0�O�Dq=C*�}%�i�QG3>w3A�G39*['�K�q�B�K����X�t7����d������毻{8��CS��̜w��r|7� 'x�ki�T�9M��@��y+1~:f�ɀ�%�H�I[�V��^�K�F�	�~_9؈��P)=o-�!U���zb���ocՈ�m�,*գ$]5E#z/E��|�;]|��:Yn�"�4
㭾�����n�N@f��y�����}:b.�au-s�� �5�C�f&�^�`��ٮ*lR��9�-����L�qg�'��xMd
"�:����I�S��������Q�D���|
�O/ƀ��,���F|	���e�)~Do�=x���xaġ�e\񴯫Nm�V'W���A�XSQ�-�����:VC5hF�Ym����J��o�͝��!0;�A��"w��nK�6��j{�a�q�Eҫ�gZY\~+��A�SWC�>R���=&B�܇*����h�Z��6NZ#vҗ����"ۅ#jJY_҅3�������e˓�p��
���c.�1;�R*"Cǚ}j������%����HQ��	}p�]�NG˕g�U�Z)�]�N�*�b@�U���$�֑�	`AX������#�|J4MB�] w�!.�o�X��TiNyK��+�9��٩�@7��3�VG��'����rX��)�ㄊ0�U����{ȵ!�h�0���?%ٮ�z�9-f
T%+1�4�L{�C�j������)�+�V�^�gTS?;3�{W���9ck\=��Ӆ믿�����P�<��� FF�Ӕ xǲ]cP�DK��/�+�	�+?�ZA�����@��$�@}�U�g � xy�Y�5`�i*�ǩ��}�-�UZ
�s{�N�&67G�#���a5B�P]Y�y1�����oP�d-2l�?j#�&�wV��[�{���a�R�Dn�y���n	;���1�*I����B/�g��>� fi5���9J�V��؞&��=�`�ׅ~�&T��T,�P��s%pRN�9�m��!d�|n�;�X��-���Z�6v�{�p���/�����Q؂�|����.\g�@c��܅�4%!�Q�V	�	�@��1'��W�m�&>}����<S�����-y�5sL��b��]�;����D��C7$Y���B�,�Q�M�B�\�Ȯ��ؾE[�tSDF�.����P��M�&�O�	�RC�4D���x�O���e��D�������_>��ɬr0��k��C�y�2z���Q�71�q��Ȣ��e*��h���w�e����o��C�t>~�=�Ū��12؆G��Y�r��4<��fz�K�ڰ��Hŋ����M�-���fIX���XwqTY-�Aoy�$E^A��	V�L�=��K�����<�;k����Q�*�=8Mթ��H����o$��l^)��k3�M����0�?Z�.�K��C1M�i�e�+�8؍�[�����~���#M��u�G��خ|i�d!j�0�j�@�h���-�K�	������.WQޡYghS������:Q�
��PX����9��E�ҁ,�\d��p�Ú�1����ify�ޕ+�l�&tw���d��2RzU0uʊ��R3gn��J?��&�ҕ-z�u�,�	��ZF��%E�G[i�HS�[/&x� S4*(��B�V|A�`c��q��*��Oȯ���L���.�	��?�^�DI�8����&��O��}%ڭ��t$�gl�k���j�e����(�!"����J��FQ1��p�&�X�$/�$�4�?_7��Ga�Ѣ��7�M�:J<��{g�� �p|�\�Y'��0Q?�JZ���0ĝz@8�e筱��)�'x
����w�!�4Z����`h`H�#��3~����i�������E���ː����[��,1̊�Ƌ?aYL��oXhP'�_
�IY�S���ᱤ�)��'��|b\�f�/����,��r�P�q�F�~m���b��Jwt�"Ԏ��RH�/� QiS}!X��x����1��\�YH3���Gӻ��k��8���[��R2�
Ě۔�}j����jK�˰���U�����^���<�"�v�s��!
�ګ����G���R<�v�f�a��j:�ص+���U��_?���V��qr*=�$�VWA���ԑ����"(xq&t<�/4����8tY�V�X��m�;���-G�9�Բfc�����h	��e>mms�}�>���Ct��H�����u��B;��׏n��7V��|.�����B�4�2��#?�

��|V�uf�4��>ȉ��Q��Ы���<�](M�m�6��2�u������t <GN� ��/�f�.]\#�ϗL5�n���'���`U£\�nI<�c�$ҟ��S��`΋���P��U�%��	v�徂��3u�y�F��z�/l`4��jJİ�1~�����P[G�kE!���7��
�X��)*n}�m�M'�s���|pm~vԩqlN�Twf�8��.��V��OKÃ���M�7r^swO��/�o	z��o�(|�ss�J�����e�/t�Lˈ��Ev��F���u.�hH����R��b൸�9�K�_�r`�LېN��?�K�v��+�`K�%��->������B�x�c0��R���"i[R��[c�bY��	�Ř��Yp�@�/���`_nr�9�ݏ��E��G��'�i� ��&�E�w��:�HYf��	��4��W�-  V^�=3�
a�E�*�hzj�BZɦ����F)�!ARW�`"s��5�`[S<�Pa
ut����C\���9(�����)��(8A��J��֮܀��.�UpG�vB��O.��z����VچrdeS�^g��"��>G"��I�H�	�2 A�J�w����K��^���1j���10��/��f��BKB;F������ȑ����F��8��ܞ�`0��T���
]Q��j�+���B;�Z!��B�ف#R�T�:������n�m��4ޅr�=�1zԳ	���Ji6��"<�
�Me�A�;Ŧ���7[�z4�Di�"��=?�)p��ż1��b��六e���0c&�N�n9�Ȣ��j��ݟ������ ��\K�JP�G�D�W��l�:L���	�;�-��r��db�������wH�.���K:���I��y��@z�n�L[�ujM���^���8"�z���e��+�|q�Ē�ў�RӵP�?������^m#�	n��sg.� �Y�A��3�I>Ď��E�*zݮ�a�'�$�����R�O:�A��)�?��
�P�F��r��D�߶�;)�_f��|tz��{�;O� �ˬ�Z���~�<kǂ�w3��0T\s×-	���O��5T܈�~S�OprQ4�n�2[���v�~$B|��t�s4�K��,>�D#�`�\����9)���4&�����_8��=gNPȳ5)�na:P�r�T�p�5�z���������r��=���6�p �g���yoN_�
-�F��t���w�E9rZ�nS,������b�J����I1[)��?M�I�U�C�W��$O�6�5��9m, g�,$�3����b�s�b>'9��n��F��)�W���Sx|/�oXo��q�C���^V.
L�U}�Չ�j�:�^tk��'��f�0G��on�X�
�y�H��"aP;�g��~��I�QͤCwxI�u�}�\�([	P;�7��bJ�X�w"�A�W[5�׏l{��Ȧ?gn{"��z�A���;�w�
�ۃ�E;+�:���gn�O����&sH�Ƈ��j�ɦ��/>!Jꋹ��Աf׋g�Z����W�M�M��ڳ>�9������o��6&�T�,�%A7�!=0�`@`�`�(�u�Ϙ����P�R=Y&@�N��I��<��~!�aEB�V��X�1y@�Y�O���q�~'���Z��̝v��ϛL���$Z��.�턭/"엄̪UUt0������WpW,*
Gbi�Z�|�`��ӻ��bU�En�ˡͱ8��eL=4���w=�T��<�r9�T�64�HQ�[��N
�^�2��λ,{����.�$eJ/��C��:���w� ��a/c�na~0/>�P��>��Ҥ�@�P�#��X.���!>�A�����4�%/�8-�FQ^�d�q�PG�f/�M;��V;Z��
�R���6�!Rm<&G���3�|f�y��^hp�ê�I�@�tPV��[iݯY�h?!����E��{��\�]cs�5��a��("����R��	��v����ؚ���c��w��@ߡv��� :�0B�(X�����%�T��ߖhm~�䩒�9��6����!քH��"Oc��'i<�l�b�{�U��6wI�rng#30��T����L#ڣ����G���A��'TQ�Q�v9���,J���C)�(����y4vV��#=q�A����8�ř�K��*�4��ղ�y����Wi6�
���X�N�2��b���P壠��U�	6/0���k�;�%V�7���c���GװoIK�ܦj�O'b_IMu�V��_�]}�"�Ś�2�4`�^g�_�U�:�$���l;������e4�t?;�"~���I?1����*��Z��UBȍ$>X�`���Nff����MueXhQ��xҵ�����b�-�﹇�Ɣh�e�wE\gt�< �Y|(��b��Q�.zt����^�b��Ԡ��,�fEq;=��]����_���䩿7i0ܓ�Y���'�GP�v���K@n�kᇤc*:x�ÇS7���;�Byp���u���	Ʈ�|M�<΅�w~͘��ҫ����s�nH]��g�&�<�ٖ�]�V���Yޢ/�4�@�K�a{J5< ���A��$wa��v@[G3E�������c'���ZQϑ-)-,Ig8(b�o��La�"e(��eX8�\G��wk�&���Y_��Ĝz�����7u4Z��w�V���	�
�{�e��/�8F� ��[�3�����2=�AJ}�����:9�5sTL�p�Q%�$��+���xLu������v�����O8�7�q6���B�o#Z�E�B����g��e����o�ܓ�L�����D<�_�
�I P�������3½T��l|OY>Y��R��_�B��ܼ����i
|yd��"������g�(��+܋?��v�l�C2�;�h�<|u�e�u�/f�/�AO���/��p��m֙�|r�?~�P�#TT[�m��������-t���3`����!1p��*�QfM:�cp]�B�:ȩ	�v��y�%֘���.�������;Q���~~����������3J�^�e�}GL]��u�^�u^^p$z@9ye���g�TR>�����ߵ�TFL��mDJ�}������O���&��CrȪ��z��2���x��g|z��Q{,X/��Fy�<.cP?��"�JR6���8-��)рu	��Ϝ-��!Tt��ݚB}�A�->l�;[u�'�$��%�-C�"������u��wl��]'_a��ҝ��V��vУ���?���/žnIŋ����mo��ԟ@�Ԟ0n�=��L���f?G��ò�@�*O�)҆�4Sz��E���6e���I'`6ڱ�\�@o~o�
j?�4�Ov��23<^w��*�5�c���s*��)]�8�U�,�Y�1'�����{S���A����}j�����U�{�*B�_z��~��W�:�|F��\p:�')�$q��(��\�֩C̸a]	}L�d���]q{��(ܮ����?	l�8őI���Y��[��f�<� �&��K�1NI2��b>�e��e�p`��"�R_t��%�[�����(s(eA�& ��zA��X���`f��wJD����E�8r��E�1V�B�4�A�P"�!=}6"k��{g�!\yV��E`>���4��)��Յ أ��2`P]D;��M��_�J����_�E��k�Y��)/��-Xi����d�']�x��/U��<8�J���1��F
�Wx|��Ag �e>���б� �38��cʵĬ���?�)wu!\�)T�$d;s�,-�{�I���
7 �м��۞!���j�Im
�k>�*�-HѾ^�$��:�wd�{�F�U�������n��Q�I^��lI�����9q�M�y48*1��W/B�wT��u�6�'�[2���� y
̗3��|v.��3ey[EH
�MA�fS�>���Y�p��N�X�zk>A����\���&�1]�ʦ�ȑ�Q�� l��rS/��?@D�"�?ڸB�\3��C�ڂG�3���!�/����=R�m&�5���F8�U{���А�
j�F�N%�XI'�7"�����k���<�vu]��`$��i:!S���چ?�Lo�1GM��%N,q`R�ۇp�.^x
�|
���(���O�V�͌�0&]�j����o�Sth���ߩA?��y�F�*5Tx�u��G�E�ZN��,���,�5�y|��hF>~���,nS�~;���+j�������lV� =B+��� Z񽋲��9�$}sZ���v�u0Շ�K��L{b~�S�2/7�Jƀ�920`�����	\�<�D�o�C��NŘ� ;�\���./�,��E�|2Φ%�d6AO��pi��@RZ�䗗\*ct�Q\F�m��Y��U8�a���9�ϸ;Y�x�S�
���296�T�=m�6zi����X����MދE���̜È��������d
�s�nr۴�ٸ�������c`_�bƼ7~���K��Іm{��QM9xg[>.�c�0� F�V�N-�1����L?r��x�[��-�a��/?ᖞh
�r�Yf�>_'#u��+�H�Z���~U���dޮ�Kج���́_jʳ`	��sl"l
��;6�Q�hP2��Sg���NxE�0��n�f�� x��PK�1J'�:UI�a������$*��8
t5�� "��u��0 ��o�tx2�w��4�E�I��F!P5���z\�*I�;è��S3�8+�R�0K�מb�r��!�F.��������7.��:<���I^�����O����m���-)Q%�:��%�j�~�=��x'��"h)�պ^ųK�B�8�rЄ��S�IQ�O�T���E�wD��e����As��gc}_�=T.k��!;-Dߢ�:����bE��?YB6{5A���?av��$\���,��@�3-/?�UD0�����M��h2)Q%��@��S|O�ն���6��	¡��j�	4�W{�;NP��U�,��S0i:\�z��T�z���G<W�Y�zW4���,�i�'������OM�H�,ݨ��u��Z���ⵦ����#&�^�8G���Qw��e�/0X�_qTNj��	�@�6q��=A�X! �"��Ks��%�F]�i���t�K7/��e��|�Z h�'c��E!�:�m� �/2�q���"��}�M��^�l�����L��5�L��c��El���#��=������JV�Z/w�Pa-gq޸��'_��ciD�i� �������\VD�~�zw�2,��^Ӈ�,^�S27��W�\M����v��iͺn01Zt{;��0�=d����m�������.��]����B/��p��н���p�g~vBQdʠaڷO��80�*l�q�퇂)gUi|�Q[y�څ��oU�4z* �Qy31�ʢi�9r]�$n�����^\�)p���O�pf���7-����4g��o�.�H�W
���ԥ�A��{���U��X/Nryj��x�j̶*��������%��<m�p�Elv��o��V<:���"� ��k����C��L&��睧�֕h��h�<����<�eaa$O�#�J �>�,�?��gt��9O��ۭ��DYu`jRYw�8�����[��[�,A_iv)����添f/���!ɑ r~��tl�R�(��O�VO���n�*�f���i�<)6��� �޲��K���kM���x�Ǎf��J�m�9�/�����$cp��v0ѽ���ߵ�_��Q/�t�1:P~�^�/b��Z|�)n���#�����#>8~�O2;���T�!d𸄫�f�Έ��8q[!�7#�D�$W��,����Xn���pڱ�^z�[Q�F�t��!-���(Na߲��x�h�^�Ylۖ���������I����k�4�X^`�j	���y���F{����nӁlD���X���Y�4�9�=��z��ӣ��%���'����]��i���om��t�>�R�?*��5	�]�	]?��x��x)�*�7�����*B����]���������k�G�����G�{a��l�1U���Ƨ���jr�T7Ŏ��-ݻ�~z�EJE��OmC��cwϭZ}������������g���[��lK��wŊ�@mv���̈́o�#��!74��D6��Em�Ɔ���m�°3�H��Y8�e�:<��?� -���#�	S&OO��d�%=�d<:�Ӡ��s�f�N���D�fh��YzfDv��?�Fep��4�G5���ճ�F%�T'8�1;e�!>#B���ax��xq�)��^�o����;���h�*>�ѸJ�
s�fy��M�*%I�;��ۛ�n�g�,!���ۄ��d��l,�J��
�{��`#ԃ/������0���9-@ء����a���1�:��6 L����(�]���"z�F�'�	�֗'
 ʛ��fM�޹@e�w����o�������ES��j*��k�6X�Jސ��P��!��4���!bWԵ
3l>�0N���f�ώ��_Īb�Y�W��9����-EΏx^;Z�5�_�{&lqi��},	48��Ғ���鲭���Xrՙ���[�"�@he{������t�WA�㿙�cb�h���Hӵ|z�\a�\�z���ޕ�>�
�)I0���k���b>�&m�B��[�#!E!T�D��_�����4ɞ�ݽw�v ��f�d��U��Y�KiL��o�*��
e�@k�wC�����G��c��GI�Q�Zn�'y�~5܁�ޠRa�C?vb�E$D�]	�Tj'b���FM�W�m��H�0����tfƛI��/�H^ �7���	�����PA��K��n���]�ׂ�0}(���g�7�3I;8g'�z�u��ŗW�h��a����]��y��?0Љ�:�������bD;��/&-����#Woi��(1nji(1/D!�ްS��b��gK�*�}孴B���JP�$a�`��:��ml=."��1?���.���35B�� ��䵵�]������"S'zPڭ�iXi+	%�0��^�Y��ϔ��������8<���/���щdz>7@��~�]�R����n״|J�4c}u��9]�y�rܒK�����Ǯ�e[���װ?���
��x\pK�*j&���ѷ�If$"hpE�&���ۗ36DV$��@�e	�J�� ] �zcbZ�T� �;>�n�[* ��]�o�Nq� K�X,����k�- ��_r"c�v�ʦo�Ɠ1s�����G��ጐj�5cZ��ybc����F6��eѿ� ���^���_�S�"��(K)*'q��BM��2�O�
G_~�R����1��,�3�znu;��Ύ����p�6U�A�Lgq��'��qEţ9=k�ъ�d&#0�wJc�;	���*��lWr��4蜘U"}5�e�o"�t�>B**�~�!�z*����uh4�^��i�,�:Ę�nN�L���1�=�Z���t:��4��cW�w��"7��X5O�H�@�Un/zv����6D&�yC���ɼ&�:�g��{�H���E��a.ބpة�,��s��|����Q�ݴ��,IsW�C:�$�GNq0b7�����R�U��!=rW+����<cȩ<��1�#�l�P�Y7���?>�/5��%O�����]�f�Y�~����,�6������J��퓾A蟤�M�:U�qc�L}V��m7���U_�fCh�̖0:ꥼO�_������u���y�Pl˥���ͩ�Tᡆ,�˴�~*.�0�U�T ��VD���;��r��#ix��>ꗲ�n��_�˰��&JE�Zv3�p�o<kK�7���b��C0˓������72�6�<5fS�^�� W��~�Q.�E��iIm���x)H<��^o�6���cP������a� �>!a��ܷ#�L{5��9G��=t��e���gP�Đf-��IK1Z�ob��E
1?�-s��C��qt]ԇ�_�f���]n���V���6ov�m�u;"_ێ��vx>���0�JR�����������+�Al`��6�y�w����:;�m���K��<]�F�-�
��?O#�Ќ�7��:���b�=���n�ى�H�;>��J�'�i�P֧� c�f5T�H�^H����'�a����EW�ym���(��I�`Ŏ@�F�J� 7����jo���\.Ԛr��2�� �Arw��q�&�Rn��]����b�r;��m����]�>����T���89Ji�)ś9%)�x�_:����U�"k;�(��#ʋ>4���͕q�n!�u�)��^ ���{��6A�J��)�7yf��	���Fy�w��?�+�O��s/��T�OWQ��lp��o����I��cd��+'� (������ui�w[cB���HɱV�՛�.��|	!�2��L>�!���&I|*t*���Gɖl��
�n�-���}�>J�x���_Ψ�,���t)`iW�Z��y��/�����ue̬�v���ͬ�	�L޳.��3�I�Ÿ�q�����1��M٬��R�a'5#d�#AVѬ� 4��Ƈ�3�yJ�i�r[ګ��v��)����h=��0��mh2��g���-*I���m�,����d�>ق�����R�g_'K�Z�{&�Wۨcqb��@���M����&X�i�A�r��H������e��
ny:��톽� �,�ι8� G_m���3S��)��ǆ��D
�3�:���<�h��6��(�����[4L��7��t��Hy��GlQ�HXՑ�"�S�½�\����`��5��R�bǂ=R�`�y!��/띹FÎ�hD��8|~�Ō:�[�6JZg��pl��|;;\.������m	�inwP��d+�#k��蹬��>�]RP	�t	A�qj��D��Ɔ	�i�͟�5#����$�-�j�6�������?&�j,q)l�.Z8���aaŹ��)�w�]��t"H����d����T9�� YEy���"ۀc�A2�h8��+������8��B��(ɕml%5�#oݍ�6�����l�܉FNuU,-�n�8h�J$�)��G�5�X�}�&�57�檡&�P�V������o��!�KD󀏜�����|����;b��?�w��{�? ��
��/5��|��x۪�exD�*
�VL<�o*$C���m�kܳ�Bv�>T�t�S��*D�^n�.ԭ��D������!�� #�*ˢ2b��|?�u}��K�ˍ&��+��.���I��t%�4U.�Ә��ǥG}%�.W�ą��*�Z5
�m���ن���Y6���������ǭ�:��Bkm�Ty����i�D��||$j�|)F�8���3'B� ��teO�:j/{~szd�5h{<�V�������?�~f�Cu�z��Y����~!��y����Ǔ�/���{���&X����M�i�{_>f�
�?d���kr��g�m�;��D�fK}U��H�#b+k�I��J����wen<L�+���5O���d�@��S��,	�2�E�k
��!��I��2h���K��@��Pq��OO��R�?��+��tQ7ؽ�D�@V���ĭ�����n{��e'ǧ�t!d��b&F�
��R�!ݮ&p|8�AɊ��� <��_Xxe�^�O�e�ظXc��E	���/䁺2�p�0�,-�z��O"v=yq g�|62�q��ȴ�J�1vH��/��g�`�Vlk֘�hB�<��w��C���7&���;��U��V��K1V��'�U�Q��w������t6�7���q����}��}0����"W,E
���ey�-
�|F�Y���Vhw���Ȃ�=���k�A*!�๓��n��)DR�5�)��.�l����p�Ĉ�I蜗}w�#}�6�ZlQ���s��Me�&j{5l�t�j_av�xRO�Qn���<ĆAn����P�*�z^�8��M�/����G���QI��\i��v�tԩ�?��A ���P��"����Jy3V�2�0$͍7pIRt �j�i�~:��J��U5��f�����+�S*��K��n�wj�0&�ܒ5��q|a�1n~�28uU�P�`O�9�L��7`d���mM.�eN�L����F���?}5��Y�����/5!�ɼ!C��j���3\�.����� z����<%D��|C���tf%/���>%0Q\ug�����1���5I��p��0��vZ5<2��;׺�uP��f��������J��%C�J(tJB��X'Ǯ/��KN^�Z��v7��gD�m����3xR�1��MI��ev'����J�<!͎�(~��%F����v������{f)��x�t2zn��X�C#���O��LTq���h�_f��!p��#M�u���g��B��ˤ����S@����[	��$osv�9�R����qGsT���p��d���P0�ܢy��E]\ī�-֫>�&�?=�P$,�Q'��۽�n�OX9�p6>��&�RTw��o�0���4I{����SK�ś��z�#��n���H	�6ԟ��̤�����g�w��Y".{�讱�?�������y��Z�]*>[��e�}�����n&�������8ކ�vV��(�=Jr��<��=��Wdtɥj��B���dţ"��̎&�t4���������;e�:�vU�]�U����y��8��= ��b�!��D�������>C��o�!W��U���4Z��V�k�4c"h�0�S�a��L���:H!��2�<����D�Hv��F����_�A�����oGY�?{�ͦ$��a�-Mv�=JIs��י4S{;�aJb��2��R�Ԉ��ڋ1�{�{ruv�%��=��u�5�-����j�ݪc���
	[�����c�Ve��������4�ip/X�R5�WWV6�^�+�%jL�6,Eԣ���!��*!��7�of�'"�//:��������Ty=G?��q�*�п���~�:�G�R��0 �Xz��Iê���8�������(��'�4*����{��w­�J�|P���N�3D\�{�Ǹ>_�%� n��,�R]Ɯ��G�F-�X��%|��� <����;7з�����t:P�5K�(#%����ʅ�VMc�@2eFa:�7��?��搄Dœ��Y���gE�5��Q�<����u�+��.�(��G�*Hd�)`B�ħ�偖�S6�?U{�Xw��u�	f�-�4JO�