��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���ڿ���͟곅	մaן�Nfsl�(�~�(A[��K�+6�K���>��iǔ��e�L���F.�iG�7�y骰�3�a5��$���:׀�0d�)�A��Ǳ&<þuiku�+�l<7��ˈ��Cwl�ϯ�8��;�����?ה�͸"X4gv s�D���	��C϶�O}V?V$VK�L��	���<��$�2#g��s�jo�3Kx�����؜�}���x�
j�}���V�OV=C�w)2��	��W�*tgPeKC��*���\�4)��Q>�D��z+��;��O�Bn�ʯ7�'��`da1�����T���W��Q�ë��0��$%룴/���� �F6�IZ��2c�>��ŋD�4Eh,Ww��*�i�|�U~$uA%ɲ�A�F�Lދiq@VQu�)<�q��p�����U�I�*/&HJ����z8����N����cʎ�A�q��_�3᜼�e�T�vy�	��يo>���юa�[�3^&XJ��]a��=���m���|��U�t��`��Bl��<�?mc�*(���d�Bߐ�������X����9sWY_�l�;��QD��v��)ؕ�8�F������{�ۄ}Ck+����V����ɥ%���!��`I�d�s�03�2H0.�Y�w�DHs�f�u-4��yږ.|�M�S2n��ui�m�C։�=���V "��xE�':�>Mn�B���S��rG����K�J��]K�sN�i��_=O0E;��t�i�Da�l�i�E-�������2��;[*�
&s��X�̤Cb{����s�F\�8rv�qY����yŪ%1�r�r�|&��?ى�4�����Gh�.7��l�/�E�s�8B�|��o��ts���m� XB��L��f{���}��D��71��v���c�"���d�=thE�,W�z��n�&ט���,,#g�,��ht(>��>�L�co�@ݿ����7c�A��B^��ian��8"�&�x�YǗm_	7.��j­�߫B<��)y�(N��LVt�A����1�FMOߡ��1�4_o����٭���v��1��A��pֈ�X�:.�301J�hB;�#�5R>꥘!���zF���pQ:���C (�	ʏ��h��M��c�]n�+n�mFR�}�y2W�s��M�T�q�o����Ŗ� k錒��T᭫� ��#Íż@o����?��;fs׺|�ǂ��=����j�!'���R�7�Q�T����Y.�E�vaz<���,�M���8�����(��9���e��/p�rh�e	*�r���p�W�M��Xs�r�[����g&���Bxk�Q��G����x-VRƹj_"�+-وf+����%���LC�'�����EC�%ק�.�Y�?}��c���������t*��[�]K�t:QKMӖ��Glܼ��{dxݫ�KZ7�Ć�>���Tk��������#�pNb:�>�vg�y/-@�C�t��	�{h�Hok������q�u�%�~�i�������W�/�[�������i"��Q��2So��7&�]�d��{��s=���yFw���R�k`L%Y���?��E>�\��^�9�̻~kr�_��3c��i"/j�s@��G�G<j�����G��V��}��*Pƨ&B׎-k��L��Zv+l�౤���Ep�_@^8��L��h���10�����ZQ)�k��o�?[=Z��$^AE[
��{䞚x�1�kۿTԯy9u�DI � ]A�"( a�͉�5JMb�!��"-�� �O�����׵��~���ⲣ��*q?��2��5��6�o:fS嵦1���w��ǉA�s��M�ۛ�X��ȧ\�.�_��#Xua1���Ri�;�d��3<�vy�vF��Zf�jLW�Ԃ>�bw�3fƥ�R\}F)L~���{K�x:���k��Yd�F��w$r��W̪U��(�E F=��I��qO;�wyL=�d��8C��7��������$����+�h�v^�����|�3���E��ڈ�UC�ymrd���5�1B�\��HS�-�Vw*��%4��V��5~�P��)r���Y��J�v~s4]qY���^���W$�P_jt=��ůV��Cܓ_馇�΄g�?��_��Q�tD���kYdT&پ\�G��.='�T�e��F�`[� ��3���ҍd���^K � ��*�V��K�3p�5�r���%]�+��s�|�;1ޤ������b�d��2���㍝j�>�!��|���eǱ\�:� T:@�~a���sv������8�|*
�خ�)�=��Jh�Ll5F�t���Ca,i����	�6�g�C�((q��$���œ+��ܒ4njLIk�|�.vL-��M��Pߘm�۵�^�"�Ƈ��^)ml�*��,�K�U��J���[T�ҡ3�ݑ�'���ᨆ������3P_f!."8�ul�X��'������S�M�V��t�{�t��<ґ�����?��
a�W�s��P�K��Q�Ab���r,�F��|�_,�q�" ,o�Ԟ����k2��~�k>7�p��r�#Qn���74��OJ���^#P�co/,.��S�U3�*-xM|^%@�Mϥ�s~�����؊3��%��/��i4���KA�7��y��mÞϦ^��N]�v�����w���c2J�y�}6%Q�=Ma%��]���D4�Y��_�V8�.f��쀴"r��pWŞ�m_�7ԡ��d��=��%)�]���I����e��ki��vg�B�\u�V/�Q^y��~7��4�ĕ�6�D��Z
<��|%�z8�i���D�W�)�ԃm���@���6v��~C�� �!�w��w�H�o��a�/�O2�i���oF�oE~�� �^&a�j3�Y����5q�
D�`?ƹ�,;5�*� O�f�:�9e����w-�@O�;���J�5L���9F!X�����߳�K�s��f͊
�d���q+X*vn��,���ǲ oo��+7��|�x=qI�${=[�:W�V4�(�}���_��JqW���.�{GH*E��2�������"#^��׏L5��05˺���S9�=��5���`�wL76�L>	E���#L�WEU��P�r?x��}.�O+s(���Y�7�_Q
�n�}�s̭�k�<��B�Bn��Sѻ_!�0I�O 0>��؍#z�=����S�ad�3*��,G���o����5
t(�xS�ƢS��Nj�'F���� \ŀ�� �
ɳE�[SFlR��@%��<ȻE����v럝�~"�h�h>&�W�\���UBT�sX������OyP�����6�����Ζy���t�6:xS��qҍ���1��<�N 8�hy�i/�b�����dFm���@���"0f��JVY�9�ɒ&�5O�7lƭ73��u�t}
v5�B�-âg0�ӧj�p���`�2:muo�x�.�oZ�dʲ�����8�f��7�\a�}J���!:�Ec��m�O`O��å)��e\p��QK�p�����/�;�l�u�˶$;�#��{�q�k͂-J�`��E������p+�9��(SF��S���+�%��U�b�\�����NN���]S1"eu�X5J�}/�Y�PZ�i��>ќ=&�~�L(��B4L׊a�����HI��8K��5싞xŦ"&�*g��z$�+i�Tv����M	?f,��E
z�����(��� ٍC�ް���nFY1'8�w����e�[�����
Y8G~��A�vÍ��[^z�x�T�X@:$�h����Yk.�����ڍ�@�����׏�m�$��	�tљ\�^,O�QH�bJ�ERS���n��"�ܭnY|ygB�"�h��,��V�#���5JjEj���$�_�3U�/�۩������IW�����[�i�I�l�bFC����2Q&�c�{�5�[�|z��dO��V���$9��$�k�^E�
�F����>;�2�L�[xs����%T-��F!c9��B��(q2q'��CD
��jr ��t
�c�̓�S7��D\�#4"pA��O�K^b�-6"]Jܩ=���)�OV���W�JNԛ�Sj�?�܅���A����k�)NA�&i�w0ON��+�3����=NB4��o��e&���Xy�e��=[W�a����e�f�x_5ޝ>���Z��^�Oaɶ���2b���08L���Hj]㠕�-���66^eH�
��?�?��*�j�
&_h��"Z�ao��1��S���5Z�+$?�0�S����ڦ�B�ԍ��2�l\7���`r	P�qFS�D���b|J-=���sن�Vz�Bk��#h �R"s�0U�h �i�4��0��x�JT�Y�ǲ)z5t�0����\��8�+��@��5Ig?���8H&�j�ʖO�� �H��o�)���J�5�h��-|x��'��NURTs%�]�z��TXK;����4�uޯ3��oM����͑[��:�(�,|�&_H᠔��X��(�E^�����p���t�R%6�!Q#�2)�>N{��0��f�%�yg@�P�|(��.���62g�^�r�_�4�n������4�`{+��ʒ��i�ʆ���k�r�]>��Ƭ��~7�d���w帓�]��ߊ�*��k�|������s�`�*sJ��{��}�kPwd�pna�!d�fOC�5����'3.�3�Q��HCp���7+�*P��ki�ݯ�A�U�)��)�:�輏袽���f�Vd���t�����3��Y�s(u	�@���b��Y�r��G���4����^1N�f�SV�\K�f���Sr�"A
�/�Vݿs^G]�����3Mtw'> ���a�|�07I�y9p� �_����������n��q�.������J;J/�<�[z`bbN��9Ş��z����!m�(�_R���^�*{l�DX���� �l��Q�}�?���iVU�^��I�,}�RWr���u�k0�YQ^$�5s��K+���s%�=Q�(��0��	l`������ �	�s����J��%r`�[j�$p>�Џ�8��v1�c�h�5+V���	Ωr�CW3S>Q�s�n߳1����v>>�Fl�0I���B�gxn��o�$��by�ZB�<�>U���r|8�9����$!��D����	Fx��T���IF xy�x���@�i8�4D�PB ͳ�Z�Q��yՇ�s=R���
��B�N�����y!h�)������Z�?+#0sڱ�Wؓl����~�%�+k���q��e���欼hDI�,� D���5�qҡۀ�u1�#����=���
�PcM�_�3��N���g��I�L��NE��*<f�TQgs�o̌�"U@k'��6�<b�^����{d҄> '����]&9���~kv�Z�w���>B�٩�8����s���FQ!=�C/'�Qޱ��^� sYfz�n���}u����Q�n��#�pS񶪬�B����*�\+�����w��6���I=5�����e�L�b:kX�X&z���d9��_}�	���7�N�g�v���:>6�`�`�_Z��ӡ��,��2#r�<�ha�#�z,W|-mw ��[t���ܸ5�1��ݸ����6I��)S#Ǯ����$���&�h;]�?pP�Qv1��ؘ��!F�:�9 ���"��-e�2s�x��s��*�T5���sf�NA�{7�(TO�^�xt{��Ӻ}B��
���Q#J��f,�� ��ͦ"\{�5����$C��Il�<�k��b����h���u�\ڕ͸�ZU.!9\*�D��-��D�[�!8 }@ˑ0�l��Q���/&� >�!�n�G�+������:�1�yy��o8���3B�!S��$1+�A�$E�#\w�Z�Q u�j9+���@JS���5����[z��I���ʿ*�����ů4�2��=៕Ǻњ%) ��<�>�V�t�&�S����I�� �"��@=�A���X'��S-��t��V���ZdX�;�X͍7LK6�0�U����v!ڞ/)<�]D:�\j�6����~Cd�����!~Q���m@��s�m��S޾�|�!��J���׫d+�n��̦k���F�q��k�p����m�ob \F4 �@��6�7!�7>�.��3N�~����(��k��������cx[��c�Y镹��9ez!7��-@RT��Z>>kb(�bT�~���7"�G���{M��Ó�����c�7��#83�P�oj��q�k��9�S���$#���剶��L�[�;��)�z��IY{��"Z@c��/���|����h@�ͷP4Vоh�3>ѹ&�Jv@r�Y��L��y8&P�`:y� ��(����E� [�~�%�9�H�� �^�̎fc��AU%�Sy⭣����e:�B.sBa5"K���y�T�`~�D@z#c��q%�+\Ŷ4���a��F��o��Τ�p��0k`����.�N�Y����K�˧LJy�͢.hy^���Ej␣��e�[��G#1�^󚣤2���#��}��JE~M�R<�K�M��K^�cL����P{*\��l	QM��e�ehĘ����̗���:G�o)ڞ���Wa@�j!$=y���01�9A%iӈ���G�_�����n��u��FO�O�i������A�	h��͸�������X�@�n��PBS�r�r�Ē�e�a���e�J!a�
v�u�`���0xv`Y�Ĥ}f(�(�U��Ź]�����M˯��]�g�;+q3�J�qnhS24g�w;מ�O]mR�Rf�<�|5��z�A�{��{��3��Х{����,�
���_����� ��޷���'��a���"����<y�e]LA���n�nł���#B5�cz*�Qv�M�����S��;�/׻��:)����I�C����ig�����=]jw��Aޣdf6��	t���3y�;V���L!�t���tGtF�]B1֚v�Pl' ������+��s8i�����k��b���x��6�N���TtXT�	� 9`��f�p�9�����0�m����}�]�Bb0a$C��$s�`�z6�N�Ĺ��6�6Ey�ө���iJ���
��l���y2��׮�o�*�obE�'�u�Ml�x��Y����X�KI�?*�7|��(����KL��Y�Q A;�Z��ƴ:+�)4�1�<�E����s�i���@Q��i��x�7��:9��Pt�5Ʃ�y~��P�����B_xp��g��~7-sb(�0��X��C�oB�U/�u�N9�*ő9<$�9�=\�p��\#��I�i@�,��E�,L�{�~�Wv!zNį	G��d��1'�0��R|I}DО��3��TcA���dR)�^�$���q����!p1�X���M��T ]/M@e
~K8M<���L?f�/yo�:�A�G����J
"[�g��}�On�ބh�N*' kX�����
�BX� �^���V�(-z�j��E:��p��ED�4�	rY� ��9j&}��,}�AP�*�.�؅��̼TBː/��~�l��F����\�1�M >4����R�3������7���}��9p]L�/�Q�C�M��7�4t,Ɍ�v�5����g����0!
�����V6
z�[h��vyx��?�:oR����,��(�k�aZ%u��g���U��������uYW��H��L�J���#�h���M	C�|G�����ޯP+Qr��L�j�,S_
R$�ϭ��8F�O���̹HD�p}�q����.����͑l�'��d���;+o�l-�=�;��~
d�t��)�Cc��qQ,-_;��O��p�|��F,r��&�<�N6��M����pP�{Dz������I�,҃�Ձ�!�t���p8��<P��24;�p'e�u@�H��z��>J6�ox�I
�,5�&m��?#z5~K��rqg�$��2����c��Q�3�������A��P�r����w��w֔p꣸֏�;#�R��h�T��3����hV�q��2*��U��
�<r�*���|��m�QW|peS f�e4?�2Q���ʤ��?�ܶ::���j)���r8L��i��!��aa��U��}]ko�Վ4:$DkY���"��Q�ڮ����(�<�S���Z�VF�RD�o�e"P�CjI�s<h4���J'�j�|�#���/-�|D;��m����6���6w��h�?4e�}���~�x	!ׅ�����S�H0W���zG��S4o���ʆ��zֿXA-�t��a(������6���f�db�!}�@������c��`��;\�$��<ST��Ԙ�U;.�:V "��0�?�w?����x��X�˄��ܖ��S� ��^�u:V����S����lU��b^%��`$c<�g<&�K9����3핛P�_щ�����zH��~N�jF�KF����$X-�9C�e�J�Շ���gin�4Ϣ)&����L����k5�Mi���	U'����nr��{�G(%���|h����w�@�e^�o�>��|���U߷!���VW.>�T~��55�l��}��f�.���ID�+gY�do�/x>�Y�D��{��v;uo_�Z]�v�������B��4��߱�Z�*�Y>�ݫ���Y/�/W+�p�b1unZ
�'��pp��qY��C�L�E��=�rsǚ�4'���l����Tݲ0����	��R�}�����()�.(����g�L^�3U;q-�v@j�9��ZD�ַը/$��_S�@����;��~2L�NC$!�KN8�G�2d}�/T0�-�!���i�lwRP�lS�����h���Rd��x�8Q���PIU�~\�|w �^��[1l_�����������H,L;��G��8�&��;G����s߶l9��S�f;X]�΍w֘j[�gm0B!h�8m�f��)�v���jՏ��a3?8�DUOz���B��
u��z���@I�Ċ:i�` F��e��,��l�+�vMb��IN�Ks!Z��*l$��za-�O\[��>���j����`���١>b�N�:3���VM�y�M�e��Hw���`ت#���]�C�橦�̔9��9O@��,U�ct2F�u6'QK�'��ӹe���?��|d=�ZyĐ~g�
�w���`�n'�G�0D6<N/ds	d�N��s�A�Fc�cX��[jVN-�W�>d�R�Dp��%C�F.J��?����݉�|�x7�S+��A����v�6h��=�����kO���M�+�YГ$��
=rt)^��ݨ�r���w\6�	v�@9�M��T%�(#`��H`ᡦv��-�:|�!�L�	�]R/�nڌ�������@��UiY��w�����o~��[)�V5�Aӱ��oLg��� � NC^}�j�֑�5� ��~�R.~Ơ d�	������/h~�a�'��0#�l�,�a���?�l-�N瞪��!Krrt�I��/���J���3�+��~�3g�B�����椰�XL��B_\�1��3�7s���%]�@꣇�喼�**�T�m���I�V渽�&�誙p�r:ϐ�l��,ɸ�.~���K��gn,�B�8�Zퟍ6y���.ًa�f�8���1�ib?��]�í���(�[p���Vy_�0�7m���1XKfu���9���qN�(y� ���g��M��n����|���α�� 2H�Ev�7/��4�� ;�`c9�b��"���$-h��F�,�](c��m�>(�PX���Зć0�l���Xqm~�ő���S�N�}���_��H�����z��%�Ut.��_��bD�_���Nb�dpNr4L�!Z����ı���nG E�|�I_�3�23I��}0��)%M�v��D��9BAѬL�5�Yy��ۅ'.:�����+YM5zz�d���'�>lW�x6�ƺ��'�(��]��8�Z��+&�)i˸��|��+|��+gsm��L1������j0��L�� k��v�K�A�Ap������G�H����,|�����j��kxr��h!�{ eSG@����g:�U��`�k�BH�4LS��V}:����!��h�wcA��F�5^P����Q�PG��s�*�s��)E>�\��}��&r-HI\�0* .l'�X��N�,�� �P=�O��|�.��(�����J|Q����:7��ϫ�bk��xLɫ�Z�ʹT�����|9�Ƨ��l����wp�O��2�UT�
�L�Ɂ��#�f��|lg�c�O�)�R�C��U*?��nQ�<F� �j��\��ܞ���ԀI��X�0*;"�?ld�X2r�տgT��:�}�z���ҌD���^���r}�
��8@P�T���+@jGj�[���(��Д�Y2���������.e2>M�21�Pq����dZ�_�aÝA^�g�NH57���l_ZNF��'�0�J���id����P���P�����9�"-y��-ǆ�D� jL.'����2��T���{ Lk�]�ԃ:2��wC�Я��2�u�2L
r��j!t�f;
S�C�d�\p _�ضF�d%��Q�����������@��%���kFͺ��_��~����*#��C�t����Ɂ�=��zX���N%S套��ս����~��v���9��$6�h����gX�6�����!�**�Z�0�	�p͸p7M�n4�zĞC��]l^��>� 1<A�SN�z����	ae9������̹L+o�]�MFw�4�)�;�����w�j}�R�LFǧ�g~̈�Q�\LCH��]k��:N���(s/l��u;Z?���V�,�R!��q%�����maB|�%��s`���%�F��JG3�6�O��B6��$7\\*WN|G�-�L�CK`g^�OY*m�vPg�7�u�I��,��&�t�\=�s������+9�m¨���6*�oS!j�� 5��MGN�U�9��O8K�S�$G�M�|���g)>��$�tT�n�I��Q�X���)����՗��ko��p�hj��y0���w5���7/A�SiX�ڗ�V,�&��DFzAyM.���5Q�C���W��)�s��z^�3M%�����. /΂Ѻ��hu.��1��i��x���������$�$���ۜӵv��Հ�G�:b���zr@�+���j@+m�(�wU�xo�<S+x�͂ 6��+,�0�� �y�5������$>)վ0�=��;e�Y���0��	5�C\� �/�貉���D�#��) ��W��U7�}E�'�$x�XM�A�W~6E���$�5hd%��-�ٝ��U/�Œ�W�
T�LH�_0�9XA<4��|{����1��/ܘ[b="�Y�%�n&�-r�5������K�rF[���l3?�x��!�d���h[Hϗ����X�{O��b΂ؼ�'�舉S��#�f�({I��_�m����(gx����7�7�^�-�r�+�[虈U-��?��X��<��ȭ:)��+;�3|!kmZ&������$���2����9��ܕ���F�B�W6�C�ք������tnmvo�G��T)-��B��*���!ƈ��;,��,��U��0a(���;M>��/?����w�)e�t�R&�o�~�ʀ��.�6�Af ���~{_yM�ݸ�zՄ'����eZQ�V��K�J6����r��&��>�Q�i��S�8)�b��� .l�a�;�vPl �|�h��.H��;��{�Y�W�򘮴��	��Ê����p~�³��;���4��X�j�hxI��B3�j��(U�to(D�P'�lݒS
*���m�,��խ�-b:���lZnq:��c�>��w�l��޸tOy�Y����/G��+�a�"�WLX��JFu��o���H��M~8��j��	g����Y�8d�'�|F3��>
�p)� �#lo��lqx���Ԩᳵ��|aM���Z���we�ʒc#�­)�İ���_lO���E�D��6 �c�k��Jx���0 Q-;���a���C�[���!}�k���:��9P#z��_��._駫=������OЀ�K�(w�$D�+�+���g�Z��f?��y)&ZT�s��3|/�S͏�C���o�ʀ�]?+b�CR���zA���5���?`�~�����Cy�5�8�~+��W��Լ����W���}WW�u���qo��DSPt�N/0�����]��X��s���7C�C�h��(��G�}�B1P��ڈ�ɺ�H/�#��V��As�xן��*�2߬'�yE?��_:�̳�p����|Yk,���p�:��fIS:�D�C,Ǵ����W'A�~��_��Nȹ�Ųt���POz��j��W���j�u�v9�CZ��Qk��>&�{v�.����@�����`c����!)*羣2/�Q��e议؞�s�D�����!�Y��?��&�-)�rW�^��
@�I-Í��;�*i�2�+j"D �/"TS�q��,�u����8�o_�0U�����YS?2S�Z�k��E׏�˛����Ũ\�"·�Ew��1��9.�U#���/��D�qG�DEx��ߓ���UG�<��<��n�9�;A��%o�\B@����=�=�P��}e{RB��p2�0T�Oz�J���Q��y��bީ�7N���B �H�z{g���`������-�B���ԥ������_e�t�؟�ϋ��X�i��4-�Њ�����rlH;'�]rQ��إ��5���v�ЉRYQ�0m!����O
tʁU1��ܡˏ��k� ���lԌ�g�u�XN�tQף�b��eR� �$�ǹU��	�����t3nrܖ���t=�U*ۣuCW~��U���{-7��Bw`hm���}�画L�_��
Z����;}.�,��?���q�y���1 �}�,-"��H�;�^�UCn� ����I��o��_�$��ǋ,���2!ٜ�]-�I�7{�2�/�����'��V8�H$�=��{p=���"�K"�(��
�f�\���k�sG�A<���=�����z���iu΄��c����QT%��G�{�sl�FǈM�M�N(S�9���a��Tѹ� L�#�f\���+l]��f�UӐ/A�[�h=�@]^U��4�����k���zX�y�^K���!/zI�g�h�<!q^2p��<e���WJ��y�!�(�qF� �!]��p� Vi'N�J+%lkﹱA��,�-O	���*��n��JG����2pt�h*J,�c;�bCc��D��?��=�4����۱�g�5԰,�^cƊ��0�/��ф(Q����o�KJE��f'���n)��+z&.�63��l���&Lx�$y�w/X��m���(��`���Oo��#�Q��$��AP����2*��v7I��]�fd	���A�w��G�L���ceg-��(�H#2�s�i�P��/�A�(c�tC�7+��
�3�b���\^�Z��ף3��)W'[�����
��j�t�Z��U���sf�8��-�����dܦ(e��oa0+;���H�oL���������jc��P-��!��J(�pP�ȕ�6F�51Q�C��F����&�O�V�IT+ץ�z[@���,�a�r��0r�M��Ik�/L5̓	>N���9E������qL�~�ANj�������X�E��;�"Qޯ}��
��P�g�3�Y��4-3�D�}Yg}�JU�C�CƠ���Ոg����[`M�Vcﳍ��~�L��7������'���9'�ER=84�b�IF�F[��S.����R<��gF.��Kϰ����E��ؖq����r�g��8����eJ�Y��ט���]���T�++�)*4e�.
6�Y��ƘY�YC�>CO�.�{�Q�$K��vꯃ��&�XF�8�C���d� �3��Y��gB��c��2���&���"H�+a�̂�EO�=�y��m��{$P�!<���4�5��Od�ǲ4>R��E{;���?>��m���
�e��w�	��e���H�m!��^ê�/�*��H����뾂+�s�m�Pg.v�3LU���m0�Ps�]|�.�Q�¿MXg#n�B����_�i��8?��2�k�9N�7�U�IP�Ƕ�\���uy�T ןY���5�(\���M��.�m,��0��Ő�]���_����s�V�(qF8u� �|�̅N�w�ږ�N�ȃ{�*(�n��n8 ?�zղ�:i�D��l$��"��<}�a���
�m��a�u�P�I���A�sv5x`r]�g.w02�!ht'�����:Cr�S�<r\�� 3f����AP|;U�����+����#�е���K��6�[�g���򬆁��/w�),.��M���D��v�!�������?cܛ�)V!��,�%i`��k���/�8S*�>�VPp�,V���j7�y�C�a(4�#Z��D�ռ�Yv�4~tn�zn�ㄘ��a�'^J�������K��r�G&�
#��#����ee^��W�Ժ<�Ұ�Ɠ�K��u_�ޔ�O�GG�_�����dBؐ��敜>��$��TEG��*7���w�(��3��X������dk}�����X&,XD4Y$�
۽Y��?A�&ˏ�<I{�vS�9��8�����D(�� ��1�H��z����E�O )/�~���Z�^
b�?�M�1�9n�,jjl������C1�����d~�9h5()t?�geG���Z���x��҇�Z�߉W���N�}J]Ѥ+�M;�:w��L���[��թ^�&��Z�V�#@��!��x4;�����:m� fznwh�w��V]��|Zm��2ӁhBŅ�;���X�0q�nעa �4�(Uo�d�ȱU�z�xϴ��x-.7�^��۠�������Y?�/�p�Y��\���UZN�G8K����MY#Ym�m�qxl"=cl��n�P4g���C-��9��&�S��d7�w�;w��E*�(������Q+1?(/�j��5��2�?���&��E}0�d�`�?����K쫦ahA��lsc�wzq�ud(tځ�!�ì�)���yqقÝ=�'�*��h����4eA]��3k������AT���5�9�٠�C��T�8�]�,�=� ��y�,6�e �m�S���Ror��F![�ܩ(K=D�@-:݋2��$���]8A��@t+(-��v�_��g��k�p�@<�S�"$�3�(�����!�D�s�jQ�`^�M8���&;t��=c]n6�������=�bA�L<�q��39�h!<?|�Д̉��h�,��ix'A/$!�;u[T;�q\�5
��STF��j�o����mC��,$�!G�qr�aH#�	�:��B�^�4͎����&(�g�Q��]�q6�.�)L�^o/�<��M۸d�n�l�')�o^ �mv���ć�y>ZR:����v6�]	MV��=������D�� ^��S4���QL��Z,�}A/�#� m ���T�6�0HK����������^MA��9]�!V渭�3�ф��[Q}3:[*w�M��2����2Dػ]��|Npɔ��5�`�<�� y������SP�g�e�Do��h^;�p�c��b��4�:�밑ѝ�ǅ*�
;P�L����ƪ���K��,z]w���E�Q���O��Q����p0���e�Y�q8x�i��@�IJ!���ޏruַ2�O��ylF���/� ��ލ)� �b@��Tu�N�w#_�<�wʸ˪�����#�>��i�ՐE�hQ��ܜ�g4%d��x.��=�N��u�QQ���j���#*���V�P(]7P1n��	Q%>�]��y>Ѽ�[�T�Z��j[�'].�]��^�gĩ@�&R���>/�
��%�$b۬����]�RKX{B��l�5 ��9o�MAe���Q$�轻���U��y
�q�O���<(]˹Z��_���WED�r�L�%1����?�|!�ѻ����,�J�8��;hX���Ωd�#�dv���>�W�WJk��p��39���IOx;��z����,�P9T�y��h�)����"'a/yv?���E�;�ь�ƥ��[df@������K��܇��d9G���{pc�!�h6�tz��5*"�(�����4��OC��@�岊PQy��2���Wfyi�. ��*yH�\fos�!���]9�vԲv��O#Qn���, �#D����E���j:�mn�k�{����ߜgv,�����*R�@�t�!5,�[��}���*_��T���F4!=�矺RU��R����Ue3k:�����Z(�9�;�Ƭ�q�߂F=7ח��q&�5��b��+d]�Z���裉�������!)��d
�i��7��W��:9���6u�%��ԿI?I����ш*�2���N�P�p]���)���իޏ_� ʱ�~��A�������il�ߪ�y��Ǘ�	��|�B�Sw��U}-��E��ꂎ#��R	8��SI�ǦP?eN6c�V�ӫ�J�r8�2�:}Af��_g Yz���(��I	R@^�y��>�gC���E�aH}VFu�X/xt�n�8pF��0��Uѻ} x�󱊸<�^��@���;���c�0=��LƼ���A��óqj�_~m�,���}�M�P�Q
�A?�"���p�+��L�}�	�`P��=�?�
!�w_��>y؅.�:����?�B��h$�0}}vQڮ)	ڝx:x��m�qc�D�%I�v�ʊ|p_�v�j�_z�U(v�<b�^��I��:a5��-"1�)�Xd��j�W��e� ůЦ�9�{̅`0U���M?��I��]�7��Ɛ��� ��1��!l�D� ����L�m�7�V󵲺4�x���5��Eomj��;�yϕ@*^�	$���"v��]-�e��B5��H#���)��b�i�5#A>�,�J���$�b���v���(����j�ϳT�ѝ-+O���z�t��P���!�e�a\���r(��籲͂���OCw�u?�ė�X��~�9�;�r���9qVr���w���1H)�)3�[��D�M����_����Z�ҝa*$�k��@��gg�޳�v� t���Qz���땭T|�Ha���N8fX�p�'�WIJP/pT���v�{�P���j�#�p��]��D��
&M��:��ӌ�J���;�j0h��Yo���K5�ŊE������q���=|h�"{	"�6N�]QAF��Y0�jy��%�s��*ps���E�,�`����iW����]�H�w�<�(O��C�,g�7�~dF�K7�~���Ď��۶ٹB<��~���)D���G�.>�B�q�����Z�x@��.7��ƙ��yOx��cv
7G��(���M������A����DQ*��_����u��ڻ�?6��<A��m��X_�s��:��aX6�x*Ciy�c[�NS�E\�eb��5��+�w8i�"l0W	�*���FP�Lj�}�>�q��,X���L�vz���"���I�3Tz�+%�Ӻ� Z��sq�����gR���3�/z:�庥��Z�k�����!�z�S�����Q�`� 	kW�hk�ES�\�7(����Ǌ37���O���� i~]~�H.vs�G�m�e��L�gYd��3���c��3�.(��T.�S��Owwq�7�QZ\M�`^wP��s�mcE��Z���O��1�K�V��u�S��H�AԡZM���
�P?�10�2�Q���/K�h�̛�j( �/�\_����k���Ӈ0g��m�`&��<<"+I��)���jp9Ј�����^⏹w����3�W.���wze����a��+��v�.��q�i��_W��(� X���z��&�{X:�ť�JtF�;\Jid��Q���g�Nh���F��ٔO_{�iC�X�l� �:��:֊�ղ��KE���)�{b;7Ȝ�o��Ý�Q#�Ƨ�`���w#`.L���Sax�Y}H���A�	{�d��_5_�����@횓�U-Fzf4F������&{�5^��2��ϠȘ��ܴ���?� �I:��)�~Rcf���[uϽ"i���r�Uífu~�J�m�S�yS�l�}��p�S�)�,�y���JY��cb�O�:�B,�怾�mء�b0�9O�Z�(�����B� �-���A_
i4���;ԛ��y,m��\���D�:�l&[��B5��B`,��w�'��.��-�=\��6"*j��F��[t%��ܫ��5^��sdv`�M����r9q�k\չW܍���iۋZ�}$X "�����[Y��k蚚4��0��8���!5�<�49��q7�u<:�W�is�8q�X��~1l�4�f��J]/:�`��k��I�a�ӛ�v�w����H��b��vW,��~��Ƥؚf��ր�����3�ʷ9�G���8ߩ�O�vu�8},�g�ïT���SZ��TN�w�>����w����in���`��YL/S��{e�i�%#�E���:�#�~t� ����1Ig4 2��p����&�b�Q������w'yêZ?<Fc������aD��xB
Ntto����W�K5/3Y#�dƇg֕����q�<ϩ=��qI����~"t�rT��f��t4g��H�6��0�ݐ�CC.���(!�.k���j�o=n�Q���wr4�s���0EJ��%�K��]��)��h��D-	��wx}#��9+�9#g�5;"�b��q�P�@al;V�z��/݁���3�fs>Q(�i�2�#G J۲�!�����7G�l�m�{��t�q@� 	=�=�r0��#�^�]Vոp�s.;��J����f���9H`�q�'	X�:�Hc����y���8\�
���|j����l皜U��(�ie�����T�x��Gw-߈ٝ��k/
��o~>ێKD	�Ə�L�rX&�![�5Lc��:���0�����,��۟�yU��<�<��>�S�>gW�b�>��N�on-�a���q/�g䁮zj��Ǯ�{Q�Ft�C9G����=��(ϙ��n��
��l������G���s㥈݊��W��m�����0�TK
�U1eg�fc�W��\�AITH�F��S���ZY�cz7��\��~-���2��,��$�[d�砺/��+���:���ؐ�U� �d�ߓ0s5��iWU��҄Q�1�+d6�L��U��	Ƀ -�]�^9!���X�,��w+��Y��%P��sCI@�6,��(V�J�	
h���4�	�`�mm<C������lsB�� �d4�t��Bx���Ȃq���2��1Y赱�M����.��Ҹ�NSf�yc���D�4�ڂ4��K�;b]>;TaB<��[��%��N�9�[�W�� �+�u�(��nӅ"��a�b�1z#�h�ڠ�(բJ��IH(޵�4��^�?��M�Y,���YR���)5.IAq�n�0���0��꽂8��"�=<�R`�rE���RFy��Q�yˀ�y��� `k���E<���2���Y\4Ըk=��k���m䀝t �j?�/g$y��'�8�!O�����6y+Ur?9�"Hv��:�^%$���#�k��L��Ij:�A��Ӧ��Ż'�_�-��<�@i�_Kc��9��[<�_�$�s$|��k1���f=@(d-Ne*f�eC�@��7�_���]�RQ�w��A�0$6��B���l��b��D3Y ����#��˕�n0���O��ƍe�}˶��@-$e��&�(�aklJ�w/S������NKǇ�>�>3�=Mw�<�XF��6����jn �G��������MH�&q�}륳%�h�j�$b��,җ_�:���v���w� �� c�?�������h
C�����P�C��xa��"�.�Qq�&|!�H{�������xow�x����is�����ۈP_R]g�4fj��_%��}sZTPcʿ}[����ߜ�9�%��W}��w)α�='^ި�~b�Nf�:�cjv�]q���fK~V�6�u���85yX����5�K���8|n��i ��E�`�eB�}��"C�VR隺(!��%����H��J�0��J��E#	h�>8�%���+�A:H�o�c^���&�͠��E$3�`���ö�WiJ��}��0Boi�������"C+	0 ��Dd4A���Ҍ*�����AQ�� �	��T	G��=�,�}a&jU�h�֭�ov"�
D��T��_N���T�i�1DNn�_������Tx�hG�eW�蘪B���L���/�r���?��~����<��Tr�N�J�� �y�ٖ.��Q�:d�WӐ=�.ɞ���͇�#�4�t�
p�çڲ�F�~��##R��F����V���l5�:/�[�7 C"�C����c4��Ů)���@�(��nU�EM�I���� }��;�j(�*��߂>W����_*�/�-��*MN���.�4��?�7��?:�<Q�������}���?5�ᗾp��(��F���q�u/��qdh�4�����K�S"�C�t�:Kh�u^�?����l�["�r�$�K-s����5�Fg6`��ʈ)k�p����%���`�G(����x����X�ݿ�Y��#���X��W�MV�*)��WM���{��P���@�����F��~������H��dn�9C`j[֌�
�
��>ڠ��0>_@��	����5�u�?�{%�b�a��tRF�%�_A#�G,�ilN�����⍫`�G��(z�Fs���rH�hqJ�y�5!��׫���^1]۽�����%�mVG ��D���,��5�
h!tz�.m����V�F�*��3N~�}�<��82?�i�sW��DhɁ�ZV�R*&$�4
�Z��|g��}������<�s�BJ��8�g���0�<���Yn���~���Y6�I_#���SC.<HNm�{}6�C��]�Iv{zt)�\m��SQӏ�������h��Z�g����� �!�\�\�g`s����tT�O���_�9Jߤ��Ff䒎O�����u�7~����~���N�>!qL&�3�`���1����d�V� ڣ88vd�)��~��K���tH@#e<��e@z�m�C��}J�}�;%��)�
�B��޹#7`ɽwӴ��ψ�M@$�uLv�����О�k-��CQ ��7��?�.K�#��s��8���X�ݪ48��_-ca���_̵�k�� `C=* ����DXeYJ��l�ƃ�߶V}��L��̭�aOe5ۂ���ؠ�}�t*��3#�Ѭ�:����y���C�x��W�~Iz�A�n�>������a��Gߥ�]�S�.SZobaD/�u����eQ���Rl+�Əf����f��;��"R�E2cJ`9��4��5�-�����j�Z�;w�h!���g;"��WE�2jU�������۲��xX�sa���"fR(@զ8�ǽ����p���з6�ߪ&?c�C �u?HDU�g�{�6#�+�r����V�2���_Crn����U�_vX|���4$�8�zR�{l�ʄ��|��4}G�b�4�m�u0��pC�y�N����\t8]:�����0n�j�F^_ޖ8]]T�=��h�p�qF�k��^p�
�2���kj)(�I4=�i5(w�g��t���IX/2��2JP'+|����|aN����`X�n�3�:y�T.�����f]�i�A*F��	��\.7p��*��|��b��**H�Ɖ�.��'�bq���~��P�z̴<�qOl��y>RQK��Zذ�@�@����\���Z����_�j����,D~4,�lş��&D�?��H�)������bv2~[
p�R�J�M��	�)w���󳜞s�ui���f���o&���嬾�v��K�(�R��h��灒���K���G��c����+��=�+���̮�h�ܭ#/�Ĉ�C�?��r���i`.B���ת�J��������+�0�|��`�#�;:����ad�E0�Uh��5� R�jm����۱����dE��c)Q�q&U�x����a���:�l��a��+Y��q}q�ᗊ��չ���f�3�0��\��c�Z� ��{c � ;��$��_�67�Ii"���*
5�d�"0�b�o� U������x(����s�i@Q�,=&�X��(�>9'Ά��i�p�V�G�������h+���w&m��t���m�qV�Xp���ؚ��<��fs��EoW[li��#X=_Dߑ�����@�C/n��4Y����hH	&A�졲qU%kj���$cC����  GN��@^|x��r�?��&�e�(��S=�B�uy�|`u�aJ֡� i+E0S���'�ɢ,�+T��YY�SMH�s��h���F�,ϘV�FQ���8���*���l@�,��(V�h�^�~�?��4�=�g�1������@�r�aہD��*)z�\�b��w���9�p��Jo��{�,� ���r���j�b�0�1�+I�D�	���\'���N�4u��!���B��o]м�k�=u���8���-e�j������yd��*�i4�41�n� @X��z�afUј�'A�Z�B|T"-{<m!���~t���{�Oy��S.4:��u�f	ꃬ_���b���f��7z[ɗ?fQ����{@y2K��\�Q�ѫz�&�BD:��σ���ݘ�6��[�����{�G&�?�ҏ�xY�<�>���P���p%t�`>h�-R���v�2R��ؒ�>����8��~���mZJw^��-� A�U�묰���{!�W	�c��W{/@��1�6mx] �Ү�!�����N��Z�u&���6����*,5i�}=U(j�~7D��C��xIC�����Mk=c�HL�n��>p��D�cfˎ�Z��F�~~�Ƣ��*��ʋ,cx��{�F2�	m)�3��&��HD��Y�oN6��)լ�.���,9��j򟒦q��`S��Z��An��
�0��t�k��)�K�-�3����I\AK�@Q�j��������;�}Pq�㱺�Z)�O�Ѹ1���A_�e��<��;��i�ɶ��.����Q����g����7i����1���8���t��M�(��c��R�Aɂ����*�������PX��@$n�&�ӈ/�����N���"u�+�{)�)[�W��GN�@:���U�~_*�m�����Y`�c��U��=~���
��>$`"�4��Ca�!<F	�Ϙ�J���t���
����M��pM��Ă;Z2p�e��>��G��<��tZ�J.�#8�s�zlQ2H'���Z�,/��I��3�и���xp����I|`����1�yV�O�ˮ���TAek4Bg2��KZ^�t�VQU\�S�'{,��Zځ$�+��%���XȀ%uO�O�
%܊�6*b^4�{��~ �y��VăP/�JTc��5\M��m{�i��b�]�#�Q���)�r%�1Po�%	/#J�| �D˝O�c�Fɗ"�|�-}�lۉ���::2EW��j�H]�::hjF5@-8�����C�J �l�io��S����c��|��`^�F��*�g@�"�E���܊�8�Kl�� ۷��<�~$�=��--��{��q�8_]����໹Ie������ �i\�Fm�8�Y*�r�@��5�c�µ�nKq�G �m<j����B��j�$� �Tw��A?��
l1���=��dE�}Lxn|��DOA�}�S�¨�ݳ�I���r�媣�4̋��[B!x/bj33x7������NwtĲ!�m�����1���&po�;B��=�5�%���`�ש����q�����v|P2��p�E�9d#�	��r�|�P�SI��g�<T���>}F��ʷ-�2�1��ʠ#��MR�@�$����|�hnR`�!��5>r���#>0[j}����hV�T�i�xQ�����+dq��r��{��m��u�0$�_$��_�׃A�*-����Y���;���~"�������;,��xzٚ��Aq�ݚ06\�2�I���.�j�
D�j�k��7����Z��/�P-�t�Dv5z7��"�.IxN�ّ���q�C7�Bvz[�&���tG�w#@���g��1x����S�#�&�LC�{��M��m2@�:�j�~�'��_�&�ۻ���p�і�Y��1�u��߳ �ǵ��"�J���K7�Z�t}m�UI�%�<�3� ~U}�����$�����N+�{tu�=��ru?�%r�Ē���)I7w�]O�k���]'��/��q���g�_噧BH�����$�j$��I:�g�qH��hγ�o���ۦ�p�B�:0"M�[���Vn����@�.w�A%SK���7G��{����9�2�-�'h_m��.�Sl���dM��<E�}�\-v�A�f������sʔ����o��/����z�t�<���.M.��<�EZ��a�RoH������}n�������Y��P$^�:M��mn�W��#�|Uΐ�o��@��_tLM5E��f�˅����^ 	��	{
�(u�O��W��,�@����W��g0��lIl^z����S��R#4�<{���f6N5@B�=�'�bi`�#�>\�]�_u���<(��(֜� ���xe��"ic�D����Ƿ6�~2���%�bF,O^���ZMA	U�`�H�~�IwuZ1�$6�l��"W�{o�xV���.l6~7j­㽴���T$�(�����@��N����	��Z�Cu���� ���r�D|U��S��-��܂��DZ|�}���s�U�s�*aD Ĳ���R������B�S�z �@dȺpEy������ �Cr�T�0f�rT�*,|����Nf�����b,o���Y��mۚR3���b^~`X�� �	�����'Ɂnb�-���3�AZ��&�G�LFn�:���0xI8,�0��p�l�ß%A՘x�h���D��l93v���R�e�X+��i��U��8�����d�
�F�4(��*0����ݞ�10����LZV�C3U�$w=y�2)!�Ǧ6Џ�j�))3��:��Ju+�;���/C�t=L�#�j��,~��O���w�8sf�U�$�}U`*�7����⭳)8R��Q:�^��!��c.�e���nD�'�$��;�_��-I�tĜ���h�	�l��Z�pT�wI������/�bn8{� �Ĝ�n�m��Je|�u)_��rـ�rT	����I"J]��C��S��?��L=�Kb��4l.�{�m��/N۩�z�'�i
Ƙ�B;#��X�}�:�
m'�+�����8,7�L|�-H���'��ҡ�5e@`�G��1�ӱEBic�)F������>&�ſ���-yw��[��f��^xx��Q`&J�t�m3��6S�X��˙��5q��6��!F0Qwp\up�_�x�I%ﬞ~���s�F��
���Y��I`d����S�tr�9��0�}�s���bj��]}�N	��x�<�dKZ6Z���Yf�Z4���P����1Q7�&���'	�P�&<W'�9��J�Ͼ��Þ�ɐhi��"������t��8�>w�S5�۠��GD�CҺfn	��\�}�Ch���C��_�>*����i��V�	���N[@!9��B}n��GJ��J׹�` K�ڔ*����F��jZ�fa)�b0�j���hV����]����_���@2ۋ#�6�ގ_��*�����&Q�)���z�z����#�<����[<�,�J��?�z�:��;�$��/f���'`�{kf�CF����*�i�@��N\����wɠ�]����7j��0���P�-y��S�j���R��z����Qǖ�^�z����j�u�2��a6�"����d�i��&d䲐�AR=xV!K>V�{����
�����?��X�:û���.ѣ��:\X��%��!i��((�L�Q��'p�W2�>��؂�x���r3��|���IE.���:ۀ�&	�~"�^[k[Xg�A*�ҿǷ��
��v��ѸZb��t;ۧ#�(���m��Mm_OO�3Q���������fCi�A���}@{�Y��w.N&��?n�<b���,,����V���GUc�����Z9U�S��psš"��*��5"Zm����1�������o��=9"՝;y6PR<L�HY=S�p�#A<�����B���xoU��O�g���	p�ϕ��H�n�!RP_?Np�S�S�Ւ����)��1�L���+
Em����	S|��9�~E��TnjN%(�tj��YZ��g��4��T}��;E���$�Xr�`a64K�R1�ݟ~���%�;A��*W��G
���h*N<��M@%�8�����>����������c2$ڻ.���p��;9�g.�*�c�K��#`h����k��:wgr#�X<e�/��l�����3�q2c�A�g2=�7]����'��o�p������hp)�����eqH�,(bDh�\:�Ku]@t�'�m$P!Y���*�A�خ>Rj�7���U���lQ*����YD�]��ʓQ0��.�B0���Jr��o�*���)�1j�M�	�I�*D�<�"��I���-���&!ͪ�ڕN	��&��c�ݿ@j,�+D6�� �c�9�%dR�n�%��)���奪���,0���Ǻ&w,� s��W�Q������xHZ����`��?D�3S�pߑ�쐛�1F��J��*Qj��PB�(�dd`Nw4�:���kC�����&�lJ�R1�pp&w���«�u������{(Z}���=���"�y3�F�Έ�-��oHn|��)~��ˌcD��@��&\+���&{�UҨ]�z�a�ܭ��ɝi�V��C�[,�T�W�P��oӕ�)����
�I��\�|GE�t��D
�L=�Z�V�MnV�����O�n+���<J�u��Y�b�c�&��bTFH��Kduc}L"V'����S1(�g�\�8B6 �'����ݸ��C��0��;4��s��S���nstգ|ɏSl�cg���AZ��+��^Ww���P* ��d/�M[��@��nX�\_��xFVx2F.mKY)�"
^~��O��^
��o���GE� ��m�9�vba�OE���`ם�K�i���记&#͗�޾�7?�<qr�wM��0G�����ѵ���n��e�CK�
�VA����-gj��ڪȹ�Ԁ!񶺳"�v��3�!�sc�"����M6��P{��:<[}��[��>T���פ�%��7Wx�hDZ}�S�D2d�ZH�H�J^O����0iA}E�}��?a��6�U+ࠇ��D5qbE�����ֲ�y�[���~_������-����s6Oc]�5�����ĥZ�7�P��{n���W���c��a�7�֞�����̒�'��}�V��{���3�Yh+U?��}�&�&�b�i�w���mA�P���~���� 􄭙�˄k�Vt����~E�}���3J�U�`�O��T�)�!f׫����{DVe�;��e3�݀��IU�yôT��08VW�����l��=��
�	v�2�+��b���:�%��US��p�7�V���>0���aqg�������LeE�1M��l�	d�5����A��T<�<{~�E�^�'�:9���a��)k���q3�Z����4y��O|���#N�`\�U���*u�������E�������Y0��c,@??xo͸��*Mj1"u�Fˆ
zt(��	4M�����>B#_�{�|s�T8�v�e�"�HG��ў�,�bT�&���j�ɉ�8<L=9{�q]1 ��^��y5fm���}v�z��m>�-�;�8Qz�C�=�zc��k�M���[�� ���*lT���#�#�N9_֩gIg���9ݷ��4	K�ĩT���/�D�A�ƨ^3�~�kW���z��x�M����]�Ώ6��l�W���_"α����<<S�E]$����z=��t����u�(�̱�@>�P�C��JB�^���M��2�cw�?xo�@-v���D6�J�	���x������ C,�>�h�����}j�95��:g8�gW��a��{�.�<�G�}����	Mc[����a�Zz�݈��H�t5�ѧ_�)�-�@��pY��]��v��5��#������	q�l,n�����0x-[�FG�v5L�O���L���(/O�(��)�VY�U�>��%}3t�)p��W�'9<���e<��~�_���uZ��zD�l�T3>�L�+q�:V��ߪ%U~�ŏ�����P��ط�p��y�ഢe�|�'U�1���Ϣ���4��{� IN�I�R[��hs��\P14��)�=��ho�Q����E.-_�,w%�v���AC��".e(�*��ڧ����Z'�x��Ê�O�2c)�������Q�K!�/� ��[���yl;�;����/��m�Z�ý�����6��Ii�f�wS�L��`�%9�o�k��/�� ����b �z�6+�ls� ����w��X��M�IL�E���ȑ' �ˢ�������ei�&5
8h��B�����t��2���ꍠ�:~*{2(��X|P��Ԥ ��T.�=*���q�� ��หd��&��%-`d&�e�IS�+�e>�E��b�p9��d��3��QxA�׃O7���XJ�b���r���=�Y����1b�S����l)@dH�����ά��:t}�]�1�0e�x
K(�+# )P��N�\Hj6�,SoQ��ˠp$[��v��Y�CU6e��w�=�=���t��q y�U,���(�8������v^ɿ�-rg;��bq_�Re�`J�#i�-�� ��a��F)�z�}����>�i��/X�m�>1[�0+_U_��(��n����Q��j@��t�W�L?i�k~&�'ņ��6p/q�U�N(6�����M�}έe'��= C�6���L���xXy�o��M_�r��0�x�HXt_�~�	������A�����sI��P �;}l���Du�f����=٘^W�o�2�chc��Z}�}�=Sʩ{s`�{��-�� @/T�v��\*WKa�_SK�y� S����Ϲ2�Sa���T!����<p�8F����MV�e�c+���[�R�sOϫC��s���L�I��Rs��ˏ��g���������?�^?v�85^XK���о�{�y{��%X�x������I�4:d��Ѻ:� �I+�%	q �؇#���8`x�z�Z��gVch���?�8n���E�LF��X=�����>�+W�s}���gƬ��Ѱ�^3�ۚ�p���jR��<- x��;$�a��-OP /	A��AOM�6�s�Sg���X_4�� n��g_�����K��3tC"f۲�#^����O��P����S�8P�`v�u��i�Xgotc�D Q2��T:�[�L��h3Ȥm��bq�
-�hK��g�~�]�Ճ�]�9'���=�8	@�4��:�C��=�&)�Z43?�"0�WF����O۶w�*����&��T��:�*��L�EtBXv�	��B΢#i���b��(�2isҮŕi,�fc/q�k`\2 �~=��D-&�ai��/	w3֘~<4ȦI��L�y��d];L7$6OW���\��Œ�U{�*J���f,� j����b��H�I�湅��sV: }�fd W�);�hBZ�_����	�V�����ۇ/S`�;�8���}z}�p�qJ���M!>]LBg�M�I,�l9R���RsBY�k����j�#+�r��xy��� 8\@��Dp�$kC�&Bm@�f���J��puy��v��е��� v���Xj:����H��v3p(a��7�G~������'\��ܧ��X[r�Nk�|�vV/e�`�z6&\t��ɖ������e&j��2����$
=�嗤��A�PͶ3�b���8���
yS,$��9��7��"1Va7��&Sv0���Hv5썋����	�W�@���VQ��ث��u:F��e�g�a�!���;b��+S���'}3e�@�N�^�?�lA�B�����I>���>J�C{�A$�xW��������O[J�2Y4��w��B�KXC�mo@1Ƕ����Db��*�����R�J.��-ߵ��c�tr����Z�Vp~͘Z��^�$n�q?��+\A�6�WT�S��_�/�6����'ة���I@�i�e�,��Ϲ��Q26Qw�O|�CKS�Y�i�������0=4��6s����ڮ ��<�[���B�[F�!_q|��pd$��4k4&?��8��_�RG^f�jj�.hv�e�F���E����S��6.��5����J���/����Qip�/[��87+',i¦�0���Xyq19� ���^�?�'/?�k� ���<�����d�-�Ȣ���x��f����b�f�[ zic_Q<r��ab��`P��h���ˀ�z%	�e�y��-{Ly��D������/(��)�z0=_��M��xbH|Q�<5"�0�ڜ�Je�2�ŅW��r�٬��C�6��P3�4l+�v��b�����-��2��E��z�J�1!�nE�a�$��]x�#i�'�;������+mv�e3��0lK�0�20-1_��_��@��#W��,��/}M]+��d��k�>Q$1(bc��1:}[%�^-��;�Nl��&Gq<ޛ��n����s3'<~/�<��~�_���X�W11��h���ǀ̈J?Y&	�\���u��{������� )�g���Y,Oe�|6�x���(\��F��$�m�^�W<���8��{���HN��I�;��GZX�hF�4�> M#ѽ@�����T��
 ��Rn�C�V�ct|�*�q�;�@�.��(g�RH��7�Y�DA�+��cS�,W�>�G!*�&aΞGV��F���H(���AF���\����_�IV4��Ť�H����j<K�S��G���`T��+���О���se��
�K�i����`�@C�����g���
ݙ�c��=�����Ѫ�|���$T��� �����L4��Ʋ�f$T�h��t��tF߽ݿf�̏����1�_յ�S�M���S�\(a~Ec˙���d�Ra��qY��xA�R��)'�#!�lc��i�=�7��zȾ�qZ]?�L�/�L׶o�/�k]q����݉*O�{9"M������P������	��:�&xW�o9��Qt��c�:��	�O x���@>v����}�H2���c%Z]�?����i��A�II�� 28o��NPq�_m�fv�^U{����S,XBGŎ���dae[ڢ�wy��Jm�����#�����C3��9JR*�ea	�j#A��u`�V&�;Okf��7M�TbKC\(�.͏1U9$܃�t?�}i3����!������
%a�q8Aвͧ}pD?'J�ySYQ-��A����-�1Ä�1B �[�Mi����~HE�P�a�k��j��P�?�Y</b���kqJ�!�/|�����x���
l�S�S>:�NxUock�)�b�.��0�\�b��RɃ#�f����hq���A�֖�p�����������x5^�p�1� ����׳��F��I��N�����L��J�M�Pi�ejgRc�����*��/߉':d5.��r�4|)�W���<0MJ��Z}���WNi9%���~��*r���͂�?8~�A�{}6��QP�P�I;B_0e��cQ��I۬��ZX�F��j��qY K�@��`�(�>'nef3Ǥdf����M���H��X[�� ��uDV�D2
O�H�E�Cc.��c�ZyN?��5z��~��q�"�x�Z���!���<G��X��EЊ
�?!����P�R!��X~" �m��" ���Y�v+�� DX�E�h7L���M'`�x�y�����Nȱ����e�EV��q:ǂ�{���2�r����~��� ���Җ�����|_~Y��De��#�E�t��L�[�(�p�=�Y۞F@e�;�ʰ����r����*ӷi�C��|$-����V}�h䘇�0k,y1�|���v2���s��&�б K��V\�4�$ė�����BI5����vЗ��;f���b��6�V������|O^˫�U�����6�<�m�L;��E���p�t���W���.	�؂��q2��z��K���jKP윭Tף �[2UE�R<7u(���C���W��6\��"q���q"��,ɫ���g�xj҇V��R�Ǥ��5
`v�T��0���H���C/�����k����n+�|��E8}R�w�i�?	9�U/!���I����pC%���$�$,���H��o}=C�f� `�}�-i�5m��cȃbO�R,��&5�<��*$J��E�_N `�D�� �D��h�q~8�}q�>���P_Z�MI%��P�	��Ɇt�'���-�V��<,���(6q�]4�wpn�Y���+\����RO}7�Fi=���[��a���8�+V�P�>[F�����Цc���
�!�z$��,���M��x3���O��#e2�٭��we ���q[R���sQ�j,�F��p'�eKh����y,��!W*+��>i ��E�j���g�'�j��U�j���:����>�V����@��Ȥ�/�������i�����ֹY�=dJ��{S��j��b�qH��j�$7�m�p��\$<�M�l�@B�I�~Qމ"��GN3��ze�7��2��D��S1��*���VBG��a����|y��y����s{D}��I,b�#�Z�'�u
�_�ȳ��y�ɖ9����P_�w	(�h����,j�<��Z���Qb��12���Js`P�H�|*�H�1��A�8��>A(O}��܋b����#�Ca�BH�&e~�Ip�4I��|�b]�͚4�G�	�D�[V�(M��zx����t��q4,bPjH���'&E�1��YyU�0�'��?���7��#7Y+��3���P{lɐl����9/\��OET2C�UtR�P<�Ag?g˖�����MA�{ԩCJm��ڲʭ�q�
��Ы�'���o��+��S��V&$_]G�������UtN�zQ��4o���'��*��R����R�Xw���lw<r�����꽑-�ؾ��V�4#YN���ķ�&\�(a��/�A-K3�"u�H.u���13l��¤�G�p�g�lX�(]]%��E=!)'y�؎�%Y��J�@&��Q���O�f��3K?��ڍ]�����z�����1C��	�~s �*��RbO�L�-2���@��NH�;���7�;�#�y������G�4�ͥjpT�O�� ���*|9y�\���8�,��(DSUA�+�R��/s�LK��L|Q���	
0��-�vl0���kt��}����']�\��}	0�c�X��wb�CikjLF���x}���.�o�&�V/G�ǉÅ+:d�㓆f��fȲU_�\׫s&�k�{���/'m=��=A�vU���!]>�����=>���"�_{���#�_Aw�X�}"b@g�9N�hf?���u��i��^fp�����.�pJ����9���	cIm�dKC�n�����C�L��u?�l�{�H�i��"e�f,F/ٓ��XU�6�
`����E��K��օ@��jІ�9��k.=雕8��U|<�o �ol�[�(���o=(c�1P�3�V��U�&��(��o�?�[M�c�S6���AT U�h\�<Z��6�y��9r�-��Ԛ��~���K�0\�s1uz�E ���Hl���Uz�U��=e׈����^O�@L��VDث�n�0�x#�њ�߂-��|P^�*�4��l��P���Wa�}k'��ۏ���2}ˁ*ӄs�t��J8e��\p}����5�e�K�޲d�m[�Px'3��b��V�/z����,�� ����i�����K�TA�[��'_�v�f�g���>K���k�����X��*X�` 7��=���0U��V*�V._�]������z-�`�
w 
I�kN���"���� �	<�x}��`�����R�m�V�p�~<�C�#&O�~[�V��7]"��`�@޳�g����W���tS�q���nLͰ�p�q\������۟[����`S��Ť��e;�X�oU��L� kH���O�g���9�P�Q�Ha����?`u�;����j�I6kl%����-S"���De�=�g��G`��o^^^A ״R�.���/��$ݯ�b�R
'Lw-8���	`g����Rc���X6��k�T
��X�t�� �^��Z�o5�0e������W�6�>���������R�gO�=�wl�����#8E��3nˍb�t?W%a�Ȼ�)���Ȫ�Q2�G����x�Y˽E�FCXXEd/A��I���n��er>�`����ٮ��_J��ܘ��O�F,��y) Sw�I;[���㩳�/X4bAU���v�+gN1Wr#�'�������;a�Q������L���ݝ?�3j��'ǂ:G�W��8.���Ae4U���ǔZw��<":!{��7�As�2�o��2���cI��OZ)� ���p\S�
U�}�3���멗�e�3�g�Jmb���]�J�s�-��'��$�n?2`��);Bob;�0̾�~���;{1x��1�[�6T�Yw�s�o�ӹ�#"��_�RS�؊���Eä���g��2�}�(����=;B�3�br�µ�����h㍊�U��ɫ�L��S/p�+���!c��|]P_�]x�i���.-�b���@��[&6�،��ol�җ�=%J�`�t��|$�j�(���#K�"i=�;�����=�o>��Ou�'Ba��DOoUM�*����T����2vk]��k6���W�߈9���rfz�8��� ĵZcW������^S�ww
�{������X���֞"�����vCj��U�#��ھ�g#t�ݯ��T}Y��?|�j)Ĭ��X���p�����C��o�J�Ƕ�_fڡ����7w�b��Ǒ)
��`�t�r9��i�]�V1�_ղ �٤^�砈-���|����Y���+�)аi����P,�2�P=�:�@Y�Ļ���� )K��vb�ٍ��\EL�dS<MoUc�E�퍅^l���+Xj+���V$�/��M[��X�q_~g�����2J	$A��v�M����<��ev3�"b<CUn�����O���a�Yh�+'G�h&��'�7��f�Gz�N����U���흯,�}��$`/w��$�x'�@�ehH�z���@yi]y�OlO����f��^�PL�>�^!T��P�����a�i勛��$�O��=P%7c���s�e��n_w��oL��2�ǛE&��N�b�Fc2mf5��/¢aogjJ�7W@�	�q	��KEJ��Kv��m�qK�j��y��O?au���Zc����d����QWv�-ȅq��2�����g��P��#]ӴkF9�� �\hK�V�E�,��n�,u(J�{��I�q�������Ac����(��B;���l�w����7h��k\	��q�6a;�}Ͻ�}�GI����� ���)�l��B �z��[��=axQ
�����Ҝ�t�<�(5��j�;�_�E�c|R�Jn�j�p�D��Cpf ��!�y��DR���gIX���N"}p�"��/�y�=���*������E7Y~t�J��� �,�����,��e�Q�7�|?�� S���ǂ���V숅�0S%�ͬ����0��g�I7�]<`@\)��?��Sz?�����'�|��t|t�<Q�QmDm�z���.�n8�~ނR��Q�3�V�T�jڬ���_�h����x��(���q��/����k��|B�����3H�,Ze�$G��� ��U�	�jTTp�D�N���l��2��C}������[�MLƂS���fl8ZB�j|�~�$҃��e�'��[�
],������r�9�	.���Z����U�}\�z#k�E"G:1�<��Z���2�:�Då '��/Ӽ�=q�Y�.z�;#Jk
�:�/j%�b��e�s?�#�]t���At<�V%6ʁ����B.�5�� ��Ր��~�9)uZ}#8�;��LD���ӛ
L4���&A����^���z��M�� ���c,�t�����zk�/O� b藋�v���r|]p��mv�W�lMy�/��-�xm �5�U��x�h��㸁��h�i���O�G��sq���V�f�2���!4��f��cΉd���s�y�6J����9o;�y)�jNê�E�!�X�}#H˚'�����X��A����kb��^-��S�vUU���t�X����mfb=�髄�oj��L�|z$ele7�e,��c(���il�r���l���B~��y�[���d�HtK�0����LR�o�Grd,�{Yx�����J���l5���
� �n���%���g�{�c�	&(����}΂���l@��2�CꋆA�z$����8<�o��T:�^��+��@��_���o�f�/�1ΗT�c�\^�@z��<��� ���ׅ��7�u
�[���p�f}��ޡYTUه2́��Zg�A�O�.7�w����{x�{��a�F���$��
<����B  �M#��#�P��#�l4�2�Gt-pN��^ZE�d���VbC]'8n�):������A�(\�A=�8�+�HP�*��S�
���S\�䏆�(�����_Q���ءtcht`D���y���_"�h��zv���e�� �sR�1��M��^�e�zO�� ���:��2R��`y#��b_yb�f&����w!�f4f������Ui��E ԧ"��� ����ݣ��!Wpݵؕ�v�� Z��V�CIv�r:y��Y[l��78��\�ؤ@�%9b��EڰC�r�g�Ü�u�q^�h+V����m�r���nc?�p.�G��27������k�1��怐��*U�d�+g_c��g��xh��W�<�݇����e+���|D���.�|Q���4Kڥ�@�t��C�Eu�:p�h
�&a��o`��4���~�ke��]=U����ɷ��بGQ��S�}��r���t�)�u��0[�dh][�7��p-�e�M;��d�Y"A��Z\mJ��2�z\�>�[�֧f1{qzBjuc�(c�0E� ��!� S���W�qD�&����l?坙� Ǿ�F�={�c��r��r���«�}�������Тd-��Ô�>����X�I�DnM�����������	uO���p �N\�>	�J�w�J��i���-ֹ��)�ۊ�έ)o\V�`h��(wֵLw�҆ʢE[�1��6���	|οRz���C��Lu��K�����D7rDT8L����j$�2j	d����5HC�ò������f��n�g���A��m�8n�~Eq��Ih)Cَ����/��������h���G��i�b�2'P�{�
nKx'u��{��9�'�{;w���Y�1�H��~���	��Y�{�	'����cu��=r��&š��n|�����a�5�/#OQ�}�w�agѧ$9�����M�'��[�ص;��������P�2������a%�|P�m��n�9����BT����H�~R�T0TVZQ]Ҭ^�+��S���K�[&]��_2�fu��ߨ���t�6j	ar���D�t����x(�������-/�?�Y����QC=y���݀9�-#��0��&��U�C��f�$��궚��zb�$�ܢ���BVc~�T�'�ZւK�[I"�AO�H�@��8e�ݣv�q*UĿS��o�ưdgG=)��a�'s�����jǇaB%��!n!Z����U���n�d��y��f �� bӤ��
n9W��yl�zt����`Ƒ�D�<��W��M�|��(����ĺ[����׊�b�z���MҐ�rK}č��T1q��wQ��Y��T��خ��f-F�`�І�B�|�;�O��a��"��f������%�z;���M4O���Ͼ���]��1��&��q�VP�9�a�������7��2]���;z7*=��6[�4�N�A�C��~�l�	]�*\6Ë%#l@� *?D�wݲ��+���jr�k��X'Ύ}��U�#�'Ayٔn��<�>� 5��B�\f`ED`�<W�f���!���ms��}��=�f�Z�6��r��n��S�>��n�Ȝ���x��T=T�=����Gs\�uPLwMݝ/ ����B�;��6ED	�� qO�EM�$~�����&,�Y��Ҏ�����O�Y�g�&<m��;��Wj:��˵ط��$�_9�����!T��ꍞ��F����ߏL� �Τ2fN�M���$Lp����pbr��'ϲU���e0��%�:�ȼ��4�B%$4a��C>N�B� ���%\��#-��6����O�-���j�l����ś����z@�����R{��_�W�W��ʦ�7N�Ӕ�
j�CS 1f�w6�O��P?x��"b&�4����rF]�eQ���_�)�p"���Eŕ��0��<�:�C�x��۟�#zu*B����c
�?!#n��c�����>z���"�B\�@p]�|(��#Wj������ē+Y���WT��+gW�C��AoB%�ٮ�me`O�U�bR��Q'��G�4��)��Z���ND�5���UpԌ���}E�4�g������"�'Q�MӖ��!7n1�S�>IɄ'a��|I���� Dj�f˲���Z,��]�����+?KH&y��\�ſ��]ΥbYQ��$�1�����V���e]� �YhQ'��WLw��ϓ;a���Fh̓�a�� �؝=yk��C���Ff�,m�F&8eef�߈�R�R����EoK5�8C,2@��Q�i����}����5��㬱V�����N�{�ʘ��S�x=��?0��%�x6�nch�>�GO���ց�κ$ d�Ş��]%�����/�c����"�-$!�ތ����Ln�m5��=���Ju��Y����\��xs�r�q3� @�C�Z�M�{�^p���?��K�����D������VU��P��W�D�F(�.n�} Q_�K�iK�3HAY����
���m��,��١��Ơ-I�Ni�J��ͤ �L̲��Qȕ���W	Y�F�+��~�5P/�-s����WG�u�6�m�����:r�H���G9�|~؜�w?ŋ�x	
��M3��Ԧ���8x���c�ai�|�&|%T ��v}Ve&Uq��7�[��Y푩I��_ �Ғ��[�6� VOQ�}�@�f��:��5�(��(�3���2T:)ˈu�҆N�]��*�ӣ;T �����*�-�{�,�{
WR\8�$*�!eG��ߴ��W4�֎ݾ�.�����ٯ���{'���jv��\P�<�/�$Li
E����:0�I�՘Лܞ
�k'8P/٠X�t-S��'���~ٖ0�%D���Й�e�X�F/">�ǩ�z�\f��'�7�ZQMe�S{a�6>���ND����ϳ�wo�Q���\%tڝrr���۩1U���f&3�����.}�~�%KU'԰$���{�^x2G���I�t�����ӝ^/S�������S1"��\j� $�t,g�Ƅm����+�e�Z'�:�����3#����F�%�Y�I�+��U=��Ѹ��b�#1q��Z��w�/�g�6�3CW�A{S�Prr��Iۇ�W���ZpbRȡd{�|EU��Ϛ��l��c�]�L������
�e�%֚͒!/�l>��;b�Un�Z�C#f���(՛Wן���8}@ωvV �|xn���v[댸�b���6e?���ߍRCp~_����
�]&��ei�:�\�}3��p�t?�X��Nhr��p.�wx�/J] ��h/��H�V�/Z���1Ћ<�k��"�S>(��F��W[��uo�$!f��(���]����>do��|�>e
����+ Pɸ�6���Ȫ��~�γ�j
n���ݹz��$TJ-�fHIOl"�vOV߇���:���`�='A���+[܆��e��Cu�-V2����es�}[i9�M��h����.��G����(j��$�杲��Yu��	�h��5粻��E_󴢾"�����E~��ɡ������Ncl��tQc�n��+���k{��W�LL�F����!]�%��3u�����\���K�]1;J|�i�_��U ��X��dA%U�P��V�_�&�Wmj��X�1*� ���0c�ɖu(΂�L���v:�B��}�q;F�	:���*�-=za��K;����ii�̊T%sM��
C>|�`�u!3��������{jS=���9?vg�j�Bm��d؛�,��bΊa�"�k~�g0p,��J�$/B�A��LC�S7��\�.�>ky3�ϫ����'��]�[g�]ֲ3� l>���'H2�??�vs&�G�0�Ѵ[�~�����gOߕ�Hז�0��Y�nD���VeS��`���}�W%~:oM9��C&��[1$�9I� zaG�����F�ioG��X��MbƊӪ�TS]����K'��嫸��c�r��a�N�V?&U�A�h���tX��7�*�Ę�������!@�Q��/oR�/�;2��K�W��c�;�#%�M��^��?�Y�O��>���h��6c�h�F<ꥄ0�4��Z�&2>�.�iA� *��ky�U<b?U 䝚KfJR5�~	��u�'c�\s����u��U��E/�y����:�<�<v�X�����&P,ZHv��P&X�u�:�!����F�g��55��^���-�V�x	����]g�1|3�^Xskyyv�	�ЈʝT�ݤ2pz�>�sD33�0x��k��G�%�F<�~���5R7���8�L�C@(�^�D÷����w��Ƹ��mQ���� N]�n+eH�U:����QO��D�	���9��2�*Ⱦo\�>��b	���7�Ѧ�;
�92��9�Z\9j��'�_��0�~(H��b��nɴF,$��XO�hR|!���D>=ZK�B�x!iq�GJ{i�AU�$<�P�o��1d�۫C�'�R�<H,k��r�N��R��-�������:{}�9b�)��{� �s�\=O��K�:GP�|�א�ܔ�v�I+��5��J��<sB�YzPB	_?\fI��&�g�`|&F!U9�ʒT��_��z�=f���72$֐�Rxq���w���L~�4w��~`9����"D|��PwƟ�;ӊ�7u,�,��ԯn_��"{؆�1p6�������w^�r����}s���HK�N�e�^��y�K��TV��#����6P�)�����0��[���ҙN���[�}�'��y�Ch]������׀�~�]�>^�!ޓ�؏���kM���򗻹�+��d��v<�J8�YT������c�:;|�d��LV�:[2;6���%K����T��Sw�eyM�q﨨�,\	9ç�O<�+��b�}�ͻ�m&I�����@��}%�� Q�XPoح��a=���'Ԙ� �y�\u�`�^OI�r�H{���Z^GyBh��F�5�4e��$��;����Dy������V��=�o{2��L#M�����-�
rnnn���3��f!8����c"�j�,�"��w���ŤTw���n	���ÔO�h������ ��E"����� θ��q3���bbd��ä��IFWPw�<��6�������b�����fdޥ�MF3�4�흇��ې^*��]:6�}Xc}u(���Ţhλ"E�BQ�+�A��;�Z�|�f�hCC�F]^���U�?o�Rj+��F�f' �!�c�[f����q9�R�C*d�JF���iFg�Q/'����R���۟��ȧ�����3��uzs#��i_��\�@ǝ'��
�<\*?�.(�J�E�%�sm�A,�"�-�5�@���7�[Y_a|����Y5�J�+"4T�H~�A�8��&ٸ�	��>�)�*z[!>��1�V�*�l��%�ۼ��[mR\��g�n�}�Q��mv��[��_<*�'�2��)��ݭ�y�Y~�~�!�Ę�(x��2WU�"�_:&H�{JG`{H���;�|�T����P�P�d��Mu-{������F���g��Vu�/����B���� (�Y���(;�,� JM9j�3~<�g����a��`C����2ʿ�D}�e��Q'渝T3��6��3(��Yb��E�@\�$�;Q-�	�nS�@\�Y�(ܟvms��g`��,��(깋��6-���ǳ�t�mɲ�J�t�F�*�Mtd
<l�)�mm�4�C�sU���df�<��㌄Q�xB�X�rȁM�0,�)��;��@)�q%8�%Bf��F��3��a�Ul�Fnr6�(�����x���seҫo?�F��/f��0��K&���$�զ��|R�ja�5���0�\������vp�� �A��Q{>�xU��uk��Щ@��<�>ɏ/����
�h��9�齬��n�=������c<����ZqU�grK_�R���տ��&7I�TN ,��CpaE�g̀�;J��:��?{q �D�q��\&Q��R�"��V��Jdw��M����/ãP�x����]��g;�p��9��/S	 ����j6 +@��� �տ?#�3��ٯ��y�]�Bc�;�E���^�Ëj?֋c����'�r@���i�7y�����-��z��A�@(�8a��? �B�0g��yY��xaԪ�b�͘!�A B0e"�|6A��<�=Ԥ��X oq\�3lUFt�;~��U���c�d�ء�o?��<�S����_�K��\��}LB�AZ�!�i��`"
 ��\:%S�u�oX9�|ȅ��>�OM\�Ɠ�Z)�� �7"֎`:��bd3��	y�")[PGy3�$JD~��BN���m'4R���G�����~,�R��P��dZ��rh����>����I�S[�݃�Y5�lR�e9��gwCl�{�d�{ɴ}�r2��+�V9YDy.�g@�.���tq(�oZ�褉9n�O�
�m���W]���ҭr��A*�y�0OWf���Y�1��O����7"EVQ��������ʣ(���x�ނ۬�v�Z��f
���o\��k�.�OH�9����J�E�,`ѝ��]�C��Fo�.ؒ;܉΂s˴���E'b.�v�����W�������8�L����GXRe-��l�(Ͳo��¯CE�]�q�=G�Ӆ8�FP�#b��!-,
��l���G�oz�7S7D�ǭ�wF�����(*M��2��j�����
�����<ZP�����b[;ȅ����J5��v�����dw�U�������u�L�8|��rꮼ� �2ŊM�x��د���[u�"ޗ��NZ�!{.<(>�;�b�Q� F����HuU�.������|�b,���x����	�������Ôj��a�O!&�m�4�xū������N�����d��&y��,�猥_#������"߶�>(��(�>��vN)�4 �A"#��(N�J�!ϴQ����E>��B�/�кi�*�~@+���;2�� L?�=^
���Jv�`�G�7z��0�N`�_4�ھҊv8��\�({~��;��K���2:�|�q0���`����CaC�T��H��
���I��q���`M�I$�~$���	 "{8}�Z�'��3��8,|avڪW^3����1����x�#�.ř� E��"���h�����?i!��5�o��ؿM�:(?ATlp_�}���z��ͽ�X�E�Bhp�x����pMk�ڸv��d��
�zk����#����'!3@��JK���J��8@��*���-L��/~�D,jw9�֒;@e�ٲ�mΜ��F���jD�u������:a��;��v�U*��2�*1h�O�pJ%+��88�-��@�������j@�'>]a�K9L�j]o�eXP��1�sN'A��D<xo&'-�[�ϖ�}r(t�P�#z>����*��@�k��.�N�`Uz'/��@/���;<��6Y������zR^�A�Raa1���S��O(H�,����r�W��G#���+ �[$?254wwk�Ǫ��	��?�CA�]Z�.�ѣ<��%	�Hj�8X�(xxU������z���.����v��M�N*{�s+�����Oɺ�����{!r�]��(��{F�?:Д,�.����pE�Fl�]n5Q����$�M��&����7Fu����4{y2�|ю�qR.�0%L��|��'���0DM����w��h]R_>�"�����|1�,D�Uu�"���~�m�������A��NOJ�6���]�k�h��N=��0ΗCCő�;`ק�X�b$�!�B$���=��=�r��rJ(x�+��6��]�N�ܞĔ�]��9�S����gzI=z?��H�^g�1#,U����fP��w��n3s�1�����q�0��G`b��;ty��K�
9��?xxY�.T���%�E3����Uő(t��5��'�*Һ>�I������UT��w3��񈞐�7��|�(]=�����(�Y�i�{��ݪm�?��59`U=4Yӧ�<r� �
��Ww>�Y#��y��BS�\�D�M��M"˨ ?I��ʢ#Q��,�1=��}�e��(mMe;@'����Mp���<!K��+k�&����g�?�uыpd�:#㫳w���!�r���A+>+�x�� {c���8��R�y�����r�D���0Rʎ���_b5��Uިׅ��������ܿ�a�Q�*;�ʓ�a�u(ؚ� �'��-��k8`}>&�(����9貴�DN���)�f)x�h�B�SKa|��`{Ǘ;�/y�L���Q43v�OpT?=LJu�C]0�`��*� �<>gYo�S6�ߗ��WsZڕ������WƩ���ؿ���Ω��B�Ll����x���d���:�'m��{6#��K�$�G�kKm9��)�Z1��M�9M�֬���z��m��y�3�_h�~s�WhѠ�⯻g_Qb2�h�^�b��c� �y��ҏ��\�p��5�w��U����ߟ��彻����J  �u�i3�� �T0lhẨ��Gt��,oPpDh���3�N�����?-��j�fx*wW���1�)�9߀���D2����z��~�2�ZV�x!��9	rG�6�V�c��{�z��T;�8�,?�-�hB��ē�{����	^oC�%2���&d���+�w�l���IB��H��Mc'��D'�Ύ6{�h�;�Oo�u���k�>���_	R��z��W�t�ߒp���r?l�a�������w��o� �S;�@���X�(*j~苛W	�� �I�.�짨s�E��巐ҫFC�h�}�=�%G��#e��2xP\��e@QF<0|b��nv�Wp��6�R�'o?֧�T�ky{>���*�5O$<fz��]��4M�M�����L�M�2L@8k���@�����A�	��N-�kN�����b@�T��]�[��	v �;$��c�����~�8�՟��L�.zcF.��o������6�(D��ӬA�&�0���;��?(�Ru��Yg���0���_�Z�?0�5��!_b���nK�bǰ���
�^y�S�/�Q��l�o�4���/�сN�� B�x��S�������'E���/V��,O7�S"EX~d:_�ރO��±�ⶍ�����z�����yb Cʪ/=
�$���:g�Г�_KX�|��Gt�奷؄J2ˇZ�H�o�@?�O���J������^qX�����K#hX���gi�U0���������;1��=#��ؼ�#�{�H�vA��%s8q+㋈�h�h��Cij�\]�f�k���D�"�����q;.)�Q��F�33 ��K�3�+�Y�j[�l����1�1y3�VU4��U��r�h��$&/�|���<�A�t�w�w<�������=Y�]�l�Z��!�I����1p�~�Xyy�5��'|�Z�$<k�/NU�\s�S8AO3� ��,���k��׺�$��G�7���ʷ� ���kC&E���m�@����v�0[te��g��&�_��CPf	JrĔA�kн]_j����P�_��:?9�p�o�O��;�t��#��;�AX�� �,@.7X�ߜ��~��6�G��l�ԗӱqY�r���t��q8E��!���1����ب��E��z&�ۘ4+�p'	ݘu��n�di�bI,8���t��[�O�"�u�h$���u�r����d1f9ԟA�|R?������D2��$v���M*J�\�� &�\I����\W(S�xvvy�*�9t���#�.ϗ��~����d	�.�Z@�R~���7�^N�A盝�"mK��Y��;��{�������T]�V���0̏]��(�y@q�t���h.��<�#B�V�.x����.��AC�������E�K�`�p�F$�]�Q�9[J����F��;�:S?��e���c&��*�?�|��'9�{Y�csjߤ�ڃxK+}�s��nS��<�=A��P��0/n�8�k�I�f��4�<o�ϓ ��� \��w���]5��޴�N���Pwә����I��ӯ	fWtƕ��饷�6�W�f����w��Xb���>(28Pa��$�+��#��>\��|���7f�wHCi�ɡ,[���_=#�[���]ܵ��R���⿖��죀�w��BH+\�ڸD����e��R����'���\l<��qK��}�A���Nt�8��(F�'�ܶ�O5$�-Vw�\�o��ӆ*�3֨�f�?����t*���B�P�mmr4zM�Q�k-�����jLUHf�hG��Y�ȝ��Q&SL��V;釺����^�I+���dgq�J~um
#�;S�a�(�y���s񨐁�LXup�N�������J�jVu�"��E�,��������K�t3���\�N��5e$��_T'��M�;5T�z+�ZTJ*���HVn��i�������p~�G�>�Wͱ\#��a�\JL�������uP��ߌk���������z"1���>�f�ej�i;Hc��!��(7�~��F!g+b�LCG��DD
́c.��R���$ڈ~�B�)r����M-��ƔA�.�T�F���?��M'q|���Pe�q�6g��*�)i@�0a�e=n�~�DlR?V����5S1z�lD��Ȑ�	-��jbn���U,c��`RM�W��ӏ�{$�-XgcZkt`t���U��#�����Z��I˯����(��O�+�/ţъ7��[e�5��G�c
�ҋI	�oM�bC�2t�M5���-�WfO��À�ߵ�icK��HjJ��s?�n6���S/HƦ�'�����i��uԙ�:8�q��`��HA�����._k�Q֟�^@�r�$iKng0�@��������PB$�[���p6tV�_���nI�iZC��vy��	�j�	^ ��ǡ���gd�@������f3WȦ��)=^��W�m�����`��+�8���-	\9h�F�F�`
=����ƅ���W�7=W����yH��h� ��Z�@�[i�x|�*ĜY@7�� �x�%Fo0�IW.��fޘ|�����	�^ӟ��!B��n��_44L7lފ�����l��7�Ѽ�L�*��^h6Q�Y��(���Dծ��3��v��(���K��?ᖷ�m[�+'�!^��m�sDQ�> �9��]l�8*c�d��${%�3 >a��D���(9�ך��`�l��6 �Fg�#`��~�)�ZP�t��U��:'��:�>�F��J65YZ�
,��_��m��Q$���iIԩ��8�Į�*4!k+!=A���"���,f����gƋB��>N_<�:3ڐ-�U�	Ǿ]�&MI�v�ନ��Mph�/��o�8]
X��d,sV[��%�����.]��D�5!j�y]S7�7qz�C�q�����^N=�-���2˨�LI:G'd��pbq���
�_9?����k����y/ݼ���B�P=f.-+��f�����'�����@@N+b�$�u��?��7zy��:�����d�Ú�w~��ה�4z������0z��)B]Ԟ��9�L��*d��x�6�p��#��/��^����W�<�E����#Z�=���]PJ{	}vث��ͫ�e�"!����Z�w]E�
\���b��$7������ob��U:��5)�|Jj�61#���l8�# �6��:�I±9ȑM�Ղ*=�,��O��4�ݦ�
}���WD����H�$Kġ�?��,l������?��*E�I�k�NN����cWhJ�Y!��Gh�R*>J�I��R�,�i9f�\��T0ɨ�{}�9�N�/�*�_2�Y�;13b%S��}A_�v� ���cm4P��v��:?�%�<����a�p�hi��y�?�	��̟��w���UpwOU6�0�M�1aV-������2�c?IX=f����.ji[�
4�ӻ�a�ϮNY7O'�ʦ�x����_�J&a��R8)/\�)�� �s:"��4҈f0�)�1r~�ƑP������5�,��VY=���iH~o���Z_�/&�Ռ�F���JxP����
�d��EH��L��;�� �^ĜCz��њ��x�8G�5GRF��,��1�,Pe���;�!H��&��cˉы�of�C6̫�aG��g퓂~�3�cf@���e�O|�v�Δ�
BzHZ�k���A	(c� ƫ��2�����$�!r6�W�p��jx�КX�yB����8���:=�"�R5 ��h��P�	F��7�no�5��&�Ǳt�-�B�G(Q8s6�o��~D}߻��;���'��<.��P�ض+8J�4�:�����b���HZQ�oH��w�8p{�k����Q�$,�r-t �0���r#�B��w��̭"Alq���0�vokoKh�}n$���A,敵n.��ǵ�Ԝ�욢:<�����@���9X"0��\�>�|䗱�7"c�	�c���2�)���eD�M0.�]����դa�dz;+;Y�D��k"��ɞ,�� �$i��&��:ʂ8]EYP�V󧦗e�	)���J��:���>���Ѵ�Eq�R.�R49� ��e�V�~	A!�h� Ncv�V1;�F��M��
*������P�oP��������W����j�E����	��Y�7�����υ �����Ǣ3'�?����a?=����M�Ļ�YĦ#}Gz?3�;z�8��S��,w�x�)�n�׼�>Đ�lL�`T#B�@�s��9��v:�Q�bٸH������
^Hm;\T'] "�\(���et�G��W�Z9	7��~�^�[A�~B��u�j�3��/��v����ȧ��`� �i�E7ͧ%��͏��ٸ�S��!ki>l���!� �e��qs�6y{,_�Po"�CL@�]�>�j��ޟ\�����Hk�գ.���a���<���&C4ʉD&�0���h|b�;�f<\��le�<��:�r�'�:��y[4���@�uI�O�}��P��^� �S"��a�D�7.�n����<�P��0�0�O�m�^���f��C;�Ɵr(ʃq�#�-es�~��Lq�� �-��x�-�����#�[��!��iOH�=Å�G3�l�����)R�+v2��:��KuN{��X��՝Uc�1|O�m��h1����BG��#��Q/͂fn�aI��Bn�D�a[I)�����}3�[��L5��%fJc{�Ύ�3~���6֙� 4�����L��;�cuݐ#pC�Ma^�L�8T�ި
ղ|���_Wu�
��9��>�|ʲ�vZ�u�I�F��y���k���Ĝ ?2� H^bMm� p�۪�&�)Hl�ֵ��O��/��G8�m�ⓙ��.�hUĊ�Mؓ����@V ��o����F$d~�#���#6����1����'j�Oօ�>*��rs�?BE���Lm��c��-A��Of��&E��^�A(��~c{���BC!�=h� ed�j�#���]-�Q����{hc�������Ϥ�eGʌI�8U�~��#�_*�k�v�ꔦsy�2��B�q�l��
'�qlhœ�x'}��E�T��}���s�t8�I�-��������C��.O���Cg�ˁ�� &"RԸt�1�>��ĩ=�.N/,͡6���^�3�6u՛p�<T��#i-�4b�)ۊ{Jt�g遀��b�T�l���� 2�tM��_Lf)Q�O�7�t�Ss ;��*����sgkW�6.����ϯ"����QxGޜ�H���a���5�nS IJͩ������>�%��y�P���I�мȬtg9��]�� 	�✚��������~pc~F��(cd
B���@��]�ŜU��Rx�`�,M��Z�ҞB ��w�݇�]-)�+)��zS�ZyzJ{%�%����i��$����
�C���_m�,I��kjk�]U�]#mQK�m���]���0�J�+ו�;T�`�A�ut��N��\�\�J5�Z�S%�[p��i�Ǐ�O�Ӣ���*=��6��v���j[��L}H�_$�z�A*�4ӥ�eܰ\dm�zΐ5X��zfmR`��7�I�!{��]��A�V�l�Shے8�`���#�i�G�z�����IL��:��a��#α���Fϻ7w��SP� �A���(�����T	u;��G*����bX�Y\�ϊ�S�禚<�_�����	@b�65b�����+��#�����T�e��nұǺ	���j���M�tɝ�s��6ℊg��ɯ���kn�(�ƫ�hF��X� x�m��(���DWl��������[��?C�4����Fa�~�
o�2ͫ�no����x"�?�5�xh)��E{<���qx����� W��}3�_=�Nd������cV�ϒΨ�&ٰhI<� vTh'��Aäa�����t���\�Z��$U�ۨ��2�],��� t�ړ�`a���d�
Ul�%�g�	Ҝh(��]UOqP~,J�ٱ?~���GPL�z�nу����TdR4ޥ�����l\)�AU�X��Uf�B�,�|9���֣p���/R��ٌK��<؄��p�VnM�ij-Sx�@�����ּ�?{\1�![Z�nx�>��Q��Dԫs�b�f����篪AA�����-H��:N{i���Z%L%�!`S��.�� 2�w�O�tǬ\$Qz�Z��CiLpǰa\L-�q���_����ZoSP�xf*�p^�!�(|�eҮ�2��kJw�=Q�]��y}�(����k3�-O����p	,���p,��jI�{P��[]EH��+�kz:�l�Ç�ɜ���-f�&^�IZ&�Ox	�����d��o��3N�\�$���p���Q�F�\�<γ9�B�o6w+�b�:#�7�_nN1}�+k֙�CI�/��OΕt]����_��OY�)6�#ީ���� �E��|<� ���R���%b����Sy��uuJW)�uz��W!�aP���-Q"�Z#��t����V�o��>�*���tM�\VY+e��m8J���ϑ�gG�[u�Z��v_�9�x�4�*�u@rJ�;����%^�~�<7]TtNm��-Qgˆ^���א9��vN�$Wn��Ma������+XoApx<��ra^#�)�,��>
zg��W��a�,���	
������_g��cT�
���$}�Æ��|��қ���_B�3�k�n�o��
��AF�4�L�H��`���r�M<��R��Ku׸1���H�f�k��=�Џ;Y|g��]DZ�����u�i���'56$�7 P�]ڀp���͠���	2�L����M� �1���B�c��Y3$��uey�yғ�y� �^��p� �D��fDw'lc;Y�����$q�T.��	�Q�QSaCɝ+}ڶ����R��v�QTܢM/��B�� �������<tA�@�W6-�1��&p+��$��k�շ]�r=��F���^��<�5�@	��6qZ�8���=�1��91��|�[�e* <{	�qQo{�PI� �j}Bn"� ����;˯�Qa�����J�m���F���hn4[\��~��4�0�z��j�Y"l�{�p�M�_����Ϛ�)V�
�g��?�|`>Ǖ�7��G���Tä�e=l�ب9g*�J51�7?79�e^
��2�j����G�H*����Q�C�.*?̜��Ĩ�9���P'��\ 0L�h�Kʃ�C4 N���)u���-�f�UCq�q_���+��U1i��["Df^FzD���N6\�������������^v	O�c�eA� �\�:E��_2��]!i>�q�g��0T�cm�ri3��ä�f�FY�C��	=�h!_�׃�@&�*�]��a/�q��`@��ܠ�?^��)�B�_�)c�o� �#���G,�<�l�}���~��C���6�-q�vq]v�����o,c���BK$�#3*�ޏv���݇��
a���͆�W��*۳S ��h���B����O�$0A�w+V�(��>HӼo}�W�(�x�Fb��ɍ&��Y��@`�#�`�
`S��T7~�H���}K�Xb��`#��ܛ��Ӵ�I��;���K�M,�:c؇,x-��6���	n��t��|�z�Ϛ�Ŧ�s� �u��ӢJFa&���W���&!u:�>�e�*.*�%�tɬIFu�r��P������d%�/d�mȀ��V��{N�ǸoyFր[��V�R<����~��F�ֵ���t8G�T�ƛ�2W?$$�>�Tz�3u�����^<E�)<�{N[�07���u�U�U��@ͭ6k�7�XV�%h���W����κ��V�p�0�r��������['f��������}	x�y����5x�> 	bm1�1m��k���>���/����/�2���,�zyAE�o�FW+��{3�̳ש�Z�[G�-�2f�}.�l�Ɗ:jvv:�3¬���;;������U=/27�[�!d\�y!j! �n:h�Q9R�}g�Gg��l,X�Y'��9�!��5b��X�ϟ<N�[:��W�3bw>��l��f�{MZu�-:�k�Z��� �P����	�p�htYl*�`������Ir���z�~���^$n.�a��/�n_�t*����^�=�W��(L�y��5��Ϳ�E�?ˢv�d- �7f[#�]�i�8e0�.`�f�,xQ�9�&�Y��t+G���#�V(�ﴈ����}�5c��a��)�y����Ke�aI���q�� 9���"t<u���<d�F�{�
�8fX�뻟FC\�g�8T1U��0P���fB�T��VD#�������!�E)�E娖��]N
lX��8�:�Jt���H����+��S>yIRǷ�ˊ|s�b�<¿Q ���J��t;/C����/���R�v�1�����d�r��Fj���Q�kP���Y!�Q5Ȯ�>[.V�maHQj��D�.���nɢ���ަ��-�ԩ�\�Ud��9 �<�}�-�#(&u"E�^�y���!m40쥤@4��u��w�m�wkp�˱w�����jF/�քh�#���Q 炊���8#�E�[/;�QJGk ����c�����|ӟ9�ɦ�#s���A�-����멱Q��c��N��s�e����X�-����;<z��9�~�F¸�Z�	��_�s���Y�FCA��4>��W��0A:�W|�����Ҵ4���X8

���xX�v@
5'�L��6�MF=y�������[pԍ�I1��W�tm��W�66������ ���9��G/)J�mGa7����{д�~f;�D1��L�Ehe�7sR�Xf�r��H�S��>&��"�6�Lp��9;)��O��i��!I�tw�0�}�1� b����h`�����Y�o�7T<��FVn��;�f���;����{�,������/���0v,! ��Z��FY�Cz辊_@P�W�PWW1�XC]�E]d�bKDr��1z�z�%���ka���H�4"�B�Uo�(�1��GG� c�i$[N�R�Db�'��}$�ن�"��`#[Ҏ�ݷ���?Ѱ�8CJ]�gp��j��E��,Pnn�/�)�q|1�cUy�,O�����[�X��Ȗ�7�k���`��l �}|� x�[I�VR:5�;�ۡz�� V��Qh� ͻ�5�O,���D~Kb<���m�_u1ŞxD�	�_�\׷
������Y4�X'S�刅���l�U���<�� e�kX.��)_�T�Ԑ���&��p�)Ν�����׹v���b���K�H�K�j��c�W�6϶j��8 {Fn�]��;�8���������͊p@�L9��!0�&��9m6}��ЭB��H�0�������F�K���g�H�穼E�����y4�!C�>�	�è�7j��4\ #zҕ��0�2�GH�v�R��/��j�ޱ%T�Ho_*)tgW5��b���PW�g'�p)���(�9j�K�'��{��\�r��>u�z���Ft
�����]Z���Q%�Pz'���N�گ����d��>S�R��\n�!� �=�I_�=Z�jD��,	�|ƒ������n3��o��K=w y�L��a�?i���,�sO|�M�U�/o�7Ec�Vv�⟘�\���?�+��Qu:G�~�>7��wւg@9^_��!obExg5s�lt���Eſ�e�H�d����gׁ��� �{MV��C��x��0��(��ʗ�|n'ˁMkfdJ�1����f��>lq&m#����	Q��x��I>j([�۔	�8�/x#U"`	���w��Mib�� ��и�?y�W�\��+��7mB�G�c��q9����[����4k��KLEb�k����q�n�F9(_k��k8к!����$ݖÕʨ�(wY�������S�w�g^������?��36�]�3� G{4��<���<���dWM���� i�J�y]��wYUIm)�-En�����"��o���.i4��dK�BVdƴe����]�Jo�O�
��YZьeo��Aģ��	��lC��G�iZT ���;���h~�<���z�%�Q?K��Mh�lĦ8a�Ph�P6�#�)O�)��AЏU��*_I�_c��ă�aM��|4;�ؽw�I���MRrK�����@�J�K���x糷��T�cr��^��$j`�'"osF�wH�b�EHh_�삕yRY(�1�؅����2x�G�rG9@�&�s|�����͚��st����q�y���!���|�%�O�
O������׼�y�$?f,B�ҟH��t���0N` �>�`�u����w
-��T��"�E-����,�&�Ҵ��w�S6���"�k:�fG��"��ɸ�	56Go"J�yYj�g����f�G>�Ό�Ղ����7Ј�N��qR^߷�4�I�7�&)eE�6��ܝLW_�?p`̳�{'�mk���7�U"9��?����_y;/����g��1�h�'��c�%�S;�钮6�&�kؤ�K䅬<v4T�m�>Y�n�hv>mO:���g���5�7I1�����a؜4�=�Q����I��П?���K�CDf~C���U������767C��[JK����^�y�qӘF�h.?Λ���[����x:�A١�[Lr�6�\�-k;_��iA������	�膺���v�-��� ���g`眿�c��J�*���Ӽ�V]�ż�˷N�����n[�����؎��;m��ek�G�L�[��WPf.�LvQѼ�ǹPel =R:��ul�*I���v�Z��z4�i���7[�Yܫ�W@*����x>ZI���WWc�e {��3Ud V���J�
�;�R^����x'9��e�;!���1�S�T	֟	|;���2�hH�r��B�Mf��ķ��sɬ�'4{m7P���[��۞��v�*w��W���U|��PP{|Hy��z��m#��w��17󈧚��Y�������j����]�6?�
��MϦ-�!�Eź�L٠J�G�u8k��K��}��|���=��.C�>�@%���A�ގ��7/�w�Ԯַ�^�V�e����?� �d}e9�
=a�q�w�F�$� ��ًyPn�?�I��OE�%/�\T�s����j�;���`���&�GO,ow�`4,պ���;����t#��J��sF�Ϲ�b*:+��K��{���8���өu�`����u�}��Ĥ��U�.-ў�\�M:54�)�s6�˛�ߜ���AM�y̻���v0@]�k�X�<�������9�W���M�
��G>8�Y�	��ҧ�ۦ60Iu���~p��wl��ܲ!����U�(B��\]��;p�V�q<T�^_�pu�z���o4u.�ѫ��w25� ��z�/1 �&�<�3>�b��1h(�w�ǋ�ې�V�eD	��o$�w*�F��^���YjP��Y��e,�m�Q�PI�T�V#"��Z��q���1 2S��e)�p�<˴��!�J}0t��x?/5�؜�S�~�.�l��]���z�}jQ5:36�(Yf��:�N|�p�6��(��֫1� 3��V)��d�1�Qj�
A�h����I![�AAN�F��=8X��@�Q��N���׎�(�S�W��ڷF����I��~C��IL�v$�٫{ӱ����Wڡ*�S0�ȱ������n����:�k'ц��zˈ�E�(��C$�bߚV��^�:�j༓���GO"n�]at�̟�q����ߐ�q�yE�Ku3S�J�jN����9�������YN˛ek�:E�(Z���X/?W^�A�Vp�y
�Tz�!�\��oگ�Qͯ��uh�	���_8��! Qm!������-^�L��	�_c���:,�p���$��{�<��X]�25oرg�PlTea:�v{96M����;���5R�]?o��&\/�-��h�/�e�_��&��>�M�,�p�h��g��%s_�N%��|�ݲ҃�Q|Er|�[�Q�_n}8vY���o	9ӑ��|����ܠ�Ol�o�ߩ����3�5 �f��=�����^�@_眛�1�%ޛ���
.y�x}SP]%��@	'��Ȩ��H~�Xw-�y8L
)�($�y�S���B6��R,��lcC�R&,��ٗ�h��O`��c�.|&���k� %C7��{����� ��-3�z��.v/�O'��C� �<;n�����T#�,J�4��r�¥u8�x ��8�������6�OG� R��%�V�a�i5j��Dx݄��s��L�`�rnHU��7w�X߃h�z�#��
���(�_!;��
 ���/�j�T���,k��mP�]c�i�h��)�v��U�t�'�)��k?v%р��Hv�G��A��i�,}��c�FU�0��Q���<AYp�`�����h�jQ��CL��[E�>-I�#j��HbϨ#롅]�=f%�r�RM�z/�/�5ܦ-%oZ�A(�=�#��'��N���J����\��˟�����/������9�EګG���U�I����ǖ�.��?�5-��r{��+>��ׅ���wY�[L8P"D��ɽ�:��c���c���_�_���xd�SF_.���&��˰��G񙯐��6��'>9�lHU���t��}֕Z*rJ�>J�s�8�u7��k冤)^AC���?a�����@].qG�޷�z�az��!����y�hԀ���L�-�,�f�4sJ*��N��� �H)��V�=�]�]�y�/�r�L8���ޭ��}���kHMD�]Yʋ[żN�3��9�è7�NL���T_'Ə
��YW�HU�YU�(!a��k�|�;��3@�Fy���,��֡1�¶P�H&�\A���(�S�����WbƗ ��~�����F�A���M������J?\�$\��p.�Ӷf���݃���g҇��ZN�|?���u�� ����Ȅ����t�򭨿�^V"�Ej�k��X��k5��9���W��{J��u��|Z���c��p�5��sL�I��ƪN�䎰��yt���:�& �W�7U�w�d��)����-gY�o��0]u�������db/O�f4���)D�Z���]�@��U��_4�1��h.��F]�F�pŕ"�p�U�,�B�$��D�v�6@X1�љ���ɑ�J|D-ȵ� �4�<�r�d�(�k��*c�4���e��q�V�ƃ<Cb�C���O����$�e�d�E]*�G�6[8y8(Xg6�1��)k��QH���~�e�g]w�^ݽ��@Y�Y���F�$޵�Z�mP��ɥ�8�����v�Lە���%i�:�X=	�N$EiQ0d佊��_��/�tkt����6���B]"�O�Χ��Z�W(Pt�2�����:ns�c�1u��]Lr����<s�2q'���lP��Kd�U������f0�E���j���(�z���rȴ���l:��v ��9	�Y�@�/�*�F�lw�Nb�!�=�R���x$����}� �n^F+�
��N$⃠�ZXE `�5)�̉��C�EC��<�_��1�^|��}�QHv��#��+nB�l�p$��x��~����l������E��Al� U��WӺ�a����z��= ��Å;"M,�g�>q��R�@\5i�Mlz�������P(�0(�.j�C.�p}˖��=�����a����Ղ�e�J��n�I-ZN��+g���ͤ��l�R���z��!j�p7��a>���O��==\=��!�]J�B��{0�~�[����ƪF~0�Ky�nnz����?�iHI"�U�P���:A��F��,6�>��@�&d佀F�p�����vQ��ڹ�Y�w�e�_Bt��|>�~��
)����B�lߟ�)Nbu#>��PV�9}(��&_ѠwW#)0F��L�mr�l����q��4;�܃�{z/�L`��We$����Vv�m
�2�L�H �$�e@��?�h������93����p��TQ2l��w��\���z�5{]f�Bi�4�J���M�G��Y�k46L�&è�r�{�7�ڴ3�jkVb*0=[?[�#8�������av��_�q�t�e���������ĵm�������(��6�\�Z]�$�(o��ԫH�A���#
?�����o�D8�&�*6��q�N���>$l[��F�p�a�0�t��@^R�?$���z�JY�h��b��^��7y�b�	�N�[��������q�>e�U	�c�N�HD
q���mٙՋ��?Iq}B����4�BN���:�[��Sw#���w�������ٍ�à[������T<���c9@�֪
��]�vF��]kQe�x��w"!W���_o���6+�D��Xr��<&��F���ڱFZt���²{�8�_4��<Ux����hI4�#IR���
	�����՛�H�e��=D�4�3�@z�MZ�ݛ>�FZT��WI��#7AK�M˵��j@��@i�u�F�0Z�	�S����=6���Z~��~����?�0xۤl��=����k���#�o���k8�@
�@�d�!g5�8���Mwp��$�\EN� ���ú�#�.jsf'�ܐz�z��A�K:f3��9]}YDI�q	8���0
Gh��BS���2�����C�(���M�E�Ħ~.�h`V�*o֔FI���"�T@ќe��M��!��q�}c�(���b����ȣ �M�S� �p�M��fG�
<�f`E�Ø��a(U���L����+��m�n�'�����rn2z��\�.x<n�y/���(�_i���Y՗�Fa�<�v�Q�_��D:F��_:��j#vĤ�,�GiW�*��O�V$�;��n��[�|��%�9�����J)f
cPCHu9�����[N�G���
i�mQ��k����:z�Ms��UD�����{�b��@�4�XE/ [�s:��2m���)���V9���_�������o	�=iSm{�G��҇���c�I�<�>x}�]�+�{�#6�~���W���t1���.����fY�z�܇���?�c0�<���	l�onr��L��Z݉.������]')�k������� ����D��1��s\���$p��m��$;�
5���B��ȓ����F�@z�S�Cj�z���fX��R��,j>��$����*���~̥�T�$tmQM���ѽdu3�J�17��!i
�:13�a�g�<T\�Q�7b�������pY辊�9�̔A&�u�) �GW؋�T��(�ӂ���ﮄ�o�]E5��uq'�'�D�1G�ֳ�We�P�W�vn����{e<�_ھh���Bx��&��Q������Gc���U�G�匲�>Q��jf�76��2�*7:���;%[�&y�e�c �f*)^i���C|�z�^pR�02VRu��O�^���,��bIA��t�Y9J�`ᙾwd��In�M�h��9�L�V��Tȕ%M���������ER]��1ZDRvzdpQ:!Zz�	��p��7��	�7�;�'�J��۔o4��.o)���f��_��ފ̇�TQ�\�=	��M���-P��|77��Z�=��k�'{�]o�!V������j� ������[�7�a�-�~h2��T�k�a*<N3���*';�֛�7U�Ba\q�=*�/vI�U���/�c���Xq{j����Dk��R���cV�j���OA�x�T�S��"�@���-*�BB��ʳʙ�!y�VX�a69�W6�&O�y�L�=��/����ۓ�#N�ճ	ql�:��k��Q���5�{N��P��(z� ���@�R^���<i jW�k �ǡ��S���'T���������L֧�*��v(�{N�s�� �:x?���zj��~��&�<�!��t(Z_������xi�)�zU�S���aW`Yp�WRc��)����;i�2��_�� qf��X�.�����Ͼ	�H��L�t �5y�p�M.�K�J���sՐ�
���=��e�Ny���t|���-�8]�w. �	��{&z6�ge������'�=Գ��]�h����X�34;֙�`C�bdN��8���pY�>��9@������X�{�ĎIgU�����^b�����ϟ�z�(�����OIy�Q�t-��Ӎ�6�j5�_w82�kq)(�e�;������jP��Ϝخd����x�Cִ._]�H��RgN%�5?N�!�����&ńKW�t֖i��<A{Xh̾�,��
��i�E����˃1juO�t�#sN��(Zg�2��R�z�'��X'��O��W�[�ԡ:�S�&]����dॖ����0��搅��5KJ�'�CE���Ǆ�ڧr}��2j�E��� [d,�-�80ksM��'q���׬IK�
�7���AI�,c6o-�zj5~;��d���׺Q)��H��|�lx��U�i�e��{��[��(����TX\0�G'^8�r��nxk�J�t���@�=¶�\(��<��6�煭�YS��j3��G�!V��!a�6>�����Ѕ�?�u{%|�Cn�#t�31d޲y�9���M��.:n���p�2���@�j����� B�����y� q��]):+&�*GJS^�(���v WBI���)�;�u�5��bQ�*���R�lSu(�9�8@E:���[�C�����M^���������w�vLA�0��k	<	}�JW���YV�C`�_ �.K�Ln�P�麍W℟"���Ň!|���.hPp,73���*��){���m�<as��E(�Z��Ȑ��#��Q;��pT�d�, ItL��SM.:r2Z���
�q�&����a`�� �� ?&n�VBv����3X8���x����8w4�3��I�|TO^�4�� �}ń������TI�� 3(X���ȱ��s[X���*5��~\$A��u�kQz�vZR��nF�3>���^<BWwO0*S.oY�֚�������0ߪ���d�ËW -V`�p��Q��\�щ[ސ�z�/�F\�S�
��A��y��c�i=._aR=E'��O��&��Qe�h>ٷ�K�`�����cѻ�]0��5c5'�2[:y�Efm��Lŷ�+��t��O
Μ�J�/�*�BV��j�gd�d�-�Pؿ�0��l_Q�b2ݼ��)`em^�VIѯ�<�>j�1�E")o/�K.����(n^�[W�H@��@�K�5�]����jA�%di�qb݀�&�֓%�v�h�YF�;VDv�p��5���x��A��q)9��#n`[��&�i`^�LW���D�I�T����8>)G��JTPj,G��JW�?�`ZR�&1.�	���D���ܹ�ΎJM�_��h��e�K%��<��QJ����(v��K�X����V� �+��bʅ���Pi�?�Q<J���쓾+�.�+���$d�;ַ�ȉn�Hw{��������_{W�t���(���9="F+���?'2Ƶ�N�>Aę� iG��E�oͨ0j}�,Σb�A�FJA������q� ���
�P�Y7��sAL�BU��b,��#�ךմ�S�е�g���YJC�z�:�I�E�r\��#�����wjRΒZ�=IQ���刍aK���J�	�q�����Y��|R6��[6������Oea��i�2�\�pKZz9GَΝ�ʬf9j�%��{\my�̚r ˶@rKu�P������S
C��51���]��K"�
y�Xq8�/��Q)��p���
J�kU��A�e(w����
��א�������1ϼO�٤�����CK4G��c�(N�D0�������)�H�jE-�9����Um�~$��h�Q(������:[F$L�������tu�q-�p
�U���mkOmҿ�5;z��	TQ�����W����]�� ����Vc����c@y>4����v5���rbp<+_ЅY���W�&���E��
e�v�>I�S�_;0\�'�D{M}t�[i��C/bM�N'�:GkqP��l~,m|�a�O=�L�ܣ�}y>K�WO7�a��S�cAGD���&�$���BX���T���Að�[����;z]�虬�Z"�q�'w��{�7�|��g=��i	s�i��7V�G�~�T�?��N�7g�\`��?MEC���͈�D'P�0���~Vh&]-ɴ�ʺtA�C�2�����/3~��Oͭ�m�7xB�x���a=M��<��v�T��9
�M�9��M�C�G��k(}�C���<���۟�fTy�M�W-K � |}��MySF(�ZDAJ^�e�~��*�e]֣�8"��ݍ+?4D�cY�ts�P�\>���/�vR��A .�ضM��ۥ>0F��m�2tX��'-�"�
B=�I�U\K1�y��������<��ru^k��o�׼�oNN� ��,�Ud��D���8�+N�"H̉�A��\�60�˼d���ηV�y+TvmS�p��ʿ�LM���ڈ���ݎ=
D[��$�"�FW0����M�����4%�.��K!7�(����B�<&�J�{���}��\WKb�Lֻ�z�n�uLܞS.1c��t���"��j�a�2���*��~����)H��+���}-��P�B�s��pKH'VB����j��%��n�X?Nl �8��=�־�q,��ª���OB	lOw������v�e64b�=�2K~�>�,��]�#v{�9�1d����_ݠI����F�s@�w�'�504����$<BW�my���e	"H27,��uǀ�=����wٺ�z��S@o�1���&*/�!��Kjϓ�
�۳�º�d�^`�e�Jay`F�P�F+7a��cM�J�>���u�gTJi+�ri�n�|{~�E%:?سr �^��-$
P�9k��^���+::\/�k.�$��1�� �~,u�76��>A�su�i���?�ɘ��dk�_�D�3�1��$����4I,>
�?�]����^�d�[�j�u]Ƥ�(��Q�Q����ay�*/h_��hy�9j�7s<��nۈh��ǖx���� 	�?*���	��������|#��S��¨م�ySU�I�K��$<�� ��èE]�E��Շ�M��#�7��cA�^|�{�c���Q<g��yt�5*,�a�h6���*L�k�Td�{�, ~�����!Y�Z�`^�-u�	���L3L�XiSCJ����@���c�t�7��"����Z)���>�
-
S��}*�ں ŜQ�+�S��wv�P��ǃ���i�uU��$�.�Y��1�U�~�zZ;-JŮ�F�h�p}�Ġ4�?�?��$�ef�)*��/�]k(�J^]���K�����&j%h�)����,��.Ng�ƺAK�M"Kq��+T;�/�W�����,�ߏ�Of�z߼l<�2N�#Q��P��9����\o�I�MZe8�E�����71(�k��+=�9��J�=�Wt��x'Q/�Cj�],S"��3V�G^ȁY@���UC��M'��������ʥ�U[� �"@��N�� (����_��kЀ��?��쾓2�6�`s���00u�4DdZc����31�d�>�C:N�/�u3&�%-�x�@;"�!��r��&�+ٯ<0�T�:���h�
!��C�Bd������QI��\ee�Pn*G�Q	�=��.=�թ&۳�@gCg�WWֈ�t�eQ�y�o�-�#=�)�~�=�����{�H��H�a����'�����D�M�(�oB�Bkn�$k6im�~y�|a�����x܎��l~�$�ϗ��*�_��Y:м�~KYX��T[cg��#�B�?l��1�7[�e����)���ӿ�����:�r̃T�Ö/�58j��,��h�n�%�>ÈF���,�ʕI�(�=C+�q�̗��]�!�Ƒ �&��Bןq���coH����:��Z�|�����s�q�3�ߚ�3�(��Ɵ�R��6��6Ca?`B3=DŌs+W�+��P�e�:�y�SO{�t��'�
�+�<��3�1��]3������l�4����#fKN!����M�Y6�Bڬ�����n�-8�o���};�f�-� �Rv��%?��oq����^��w��f�G�Fo�7�;e��0ň���q���1I����o^BM��}�G�K�f���+Ot�@�|q�VA�Y(���b��p�&!΅��<��q�2nI���qR�m�fK(�}����<��p�>:��vxdw�Y�;]�T�̠�OL�鎹��I����6U�x9��^s\����K����g.	����%�RN��G�Ec�x��_Uu���o����"f;�M5D�B�ޱ<t�}T���/�l���p.C�����Q�����M��or�� �F��#?}SVG#B2�����'��3�R�f�\#���='�����x_�T���1���? �}�T�{;�&����."�r�Ƴhݧ �&�PN�������b�b_�a���zǆ�I�}�Ԗ�0Ԋ�ϴ���l���8��EQ�ˋt���<_(��j0$Lv�u�]+#���S�����;�ǴLd~���y�]aJ��K��/_����Ď?Z!i���'��������s oV��w�6`b�:�>ô�d��)�z{��� 48���V"Y����,���7:}f&�"��y"���cI�	�Jq��kL���1���":�?����{5Z�<��� �YTa@ۇ����D��ɏח���9�l"��e��{���rô'�5�,}|#,Z�J�|���ɝwI܌�m�h*>;�g����;R�e���Ւ����$�D��onS1����3�ϊJ�U_�g\�����Ap�j�"��p��3���l[$��/��^&���eƖ��^6LE�-�S�]�n���XA�4\��p��y�q'6�Im���Xݮ��%,�'�d*�?ũ���S�?�ɛ'*;m��eq�u��u����
�����Hь8��Χf�Z�!j�%8}����g�o����ڝ��Y�H���8�\%g�G���� v@��lo�\=��@8��+���1#+-��dO�e�;]%�r}ls�s׼���O"��nH����tF��e�#$Ղ{P�+xO
�o|�=]Q��	�Z�ȁ͛xC���n�ӓ_��}���($(�<}�]�ESk�l� o������[�b���l�n!7/">�k���T�F���B��˙VH�S*A?�9��f��i����7�.0N�q�c�K��-���v٘�喥e�$z�+����*�������]r1t[��DI8�G��[�(��vr�c���n&! ��6B��������?Є�C�ٷ"ݑ��3�D6��݂��  -��%�v��� w	'G��mX�?���'��Y1��3��-'��=w�gW����[3�D��D��9E�O�m	"���$�g�m�T�w�GGн�OO�X�AB������}]�7�bE�py�����u����iߝ-�҂�̮kEw��w}U��-0�E[~%��i&�����>�t��@]h�]4S�ΜI����SZ��?;o}��{��� tu&�	� 	?�Ѱ嵈= �z��|W�&���j(6�;���2Ʋ�w�z�xtS�zb?�4�j|��!�`к,��mB*Y� ͘�ZTV}K2*��u� ������lDvJ�q�uV��S/T�Ll�Ϳb	)�w�KQw���<��˭�z����L�)�o�@a�y���O�;��\�;FI_$N
o����"�]&��U+����gt�Ƞ)k���r\���衲Rj,�����61H��U5JqРf�k7���J�#������w�v�m�wۈ�5n���.ݎ�4���`k
B} �+w�EXd�n��{g�$~�|��L��S.�^�d�ܸh�<��6�@��.	�z/U���Y�ߛW�8Z1xH�0�Z�P�8\9�)q��AmT�ܹ{�@�O�Qә���M�G�,�	��*��	
�_�rp��4��Yl;_��=�n�f�q����؝q�o�+�E�ć�y�=�)�
a�p=�9T��4?Ic��<����*�}j����J�N%�֕�ⅠC��;�w�UdQ����#"
X�7�b�s�p�i�;�Rl`�5K���Dw��RF��-����N�ߣ�<��Ê-�3J!~&|.���K�R�����9j�|��mŚ��rm��¦cx��\�9N\%�s�U7c�h��L�@ya`�5�;)&t'66�e��y����L��z�Vv8P�?���	�����KZ'�L�G�@�� ��+�	�<���P
�F<�/��yr�HI +���Xj��r���td�d*�x���g�C�w�ˁk oB�Bt�Ɨ}�2|�A M�bK��:��W�;�[�Ț�ۅX�G�6�������O̭��O��OS��P[�S=���4��#����"�I��D�*1���˜��_W�$J�i��r�\p�!�g2�m�op���  ��i��B�o+$�ENaT��7e�ɞ �%����o3�����x j����3��gN&yn?of�ʼ�=zP��3��!S��#@�������2�;]Oc��#%����ǮX0Qʶ�5M�)��Q�.(��湤���J\I���sHh���Ai4��
L�$��!����K����}�í��&U���]%T �1�Q3m���X��V��,�q�9Ӆ��|��������_���^�>>U<pA2�+�Y@3|>Un���3|�׭�v�п4�U����5���L�Sy_�H�:seMɤ$�
�(����cz'^n�R��4hV�cL�y\{[$�R��?�Q\D��/�%�ѴD ����ȃ���O�>`�v�Q�e8�NSlA��Lk�j'�J��a��&��p��y�mƯa�EYݡ�c�m>�a�yş��~�}|��Q�ӷ�v��XW�����X00%E��+5_�9GuY>����؁8GQa��e&*���'d�
�2a틉xˌ�߳�mTHv�TZE��8Nǋ� �	�}����O�>G�\iqv@O9��@��v��Cǘ^\�H�y�*x�援�J��ą
�
c<�bۂn��1$��dr��X��v�'<�x�#��	<�ٶ#�,F
��ЋB
�z��ɘ��+�y(5����/�>��J��>h�Ԥ��d��1�I�J,K)L�H�X�6�r�B�o������%Rʶ����E�7`��cnN[Ȗq k�b�<ћ��tY0��8y�M�'KB��W!����S�Z�ښ~���q�hG�h̍T�)���'�('��e��(M�����U�w,��1��O���C�l&�L��1�5�9 �:�	I�(�S[$+F��4�E��ad(=����#>}��
k$	��v�2}��]Hf����[�(����UxN�D��}�a��6|T#8��,g�΁kq�o�R�6���!PGn��7��erzx�>��l
��I�!�2�`$����pK^�X�{�,G��)k�����ʲ\��TP5gT�ؕLO�!P$�j�N�{qg(��C�����	�O�1��M�"ُYuٲ��/E図
��jQ�%4>v#箳����U |���k�S^�e��OY86���Z ��xk	�Ck؆0��`Z�b��[��r�5k&�]3B��`��qd7�2V�b�4.�p��\�.�q��Y���$���*�l���T8�6�ѭv9��j׎/�N���JϪ�e�ޏd~V��.}��裗An0h�A�6��,S��L-�ɐx����L �ɔsݸS�h�{� As7"�9����2c��K�i����Oh��"�=� ����mI�Ea���$N����i����N��w����te�*������L�!��C~�����5I*��_����v����SVv���㵆r��*ۚL.�)v�h�jaP
�e�y_�J�k6��^_y�[�яX��K��Е!�ם����qYV�b}�"*�)��8���V�f։�:w�B0CA�B��9��:% ڕ����)��v�0h�G���i��i�9�9�b%B��c�\A�TJ�4���?�5���;�b���)�f5H�O��-��j�1v�[*�|> }�@�'����w^u�W��ڸS���&0�q�5�'E��q� �>b� ������/�Ē`�����H~��X��\��80p -�^�����;�m��#�s[4wP�2u���`�ّ����VVJ���\�(�N�'I�:ˠZg;��2;&��Q�f���oa� ��zߗ��P6Y�
�g�K�����6��h���.�ދˍ���)ёIm1�WD#���)���Y#i:Zɲ�OU��X]�`�9&�!Nz��u���z�>���m��./��5r˥�Y6�<)[*�P��xcPk���,���;�����gV�Ϲ��ۆ����7c��u���� Z��.^!�!%BN+�BE��X A>�'f�ܳ��z�:�Ӎ��yX�_��Qķ<�cTH�h0����׻���	ڑ[�ǟEEok���T9�Yw���e�?!+H;3U�0n�܂2
����q
n���1`Wm�I:��#�&C��"�Q���9���+���v�
�
����?�1�����^#QZ�e ��"�Ue�m��=ꮲ���3ٲ6�YA`dr_��n͉��k@"0W;��^D����s�=dʫ���E��
��C(�Nm*�7F��UxoGLx��`b0��&������y�+A�-(���xT�u�����0ð�����g 1��-]�7h��ᅯAI�U�����v��{t&D	BM�|F�-{�bɡ0�囖u/��U75�7�FD��dG��lm������MV�i��=�CŞd�FC)aa:�����K���:j닦^Bk�b��.��iDq�T�C_�5*��K^��Fǝ[>؊V&Y����?���V����,�I�����fǊI�S�Y���U��hl�&�N(Y��M��YJjR���}�3��*������0�Aq��3��#W���[���;a�}���ۧ?���ז�֙�N�g�d� ����������6����7I��UC��rZ�ɆPBg�\Zd��sS�c%�3|L1#��N������:���7z��𐔋Nr`F�sy��t/O��V$f�C���|4����_@��UBZ��G!w�@�4ū}��5(z���v��RW-6�����E���D��s{��~M����h�+2:��ܘ��@%���>����I+x Ȉ��Z����cw�0V!�e����T���g��4��,d�6)� lt+�,�Ei�����:W�
�~�����`a�p����ݺ���!���+/YvdBmhs �� dF�%Y2�����n9�]��s��0A�o��.��i!Dm���fcK���`)��J��c��R��1�M����d�J/`x�l7�C%F��<
��)��A�o������uc(�?d5��4��f2�����%�#�'o�A$�W~���٥K^���ϔ�;�}�1�AY��ק�.C�|��Z���g��y�>t0�H��!ݿb��b�E�7L@h�CLhi2��%�U�Si��-��4o4����/�H�P�	�	K$��^�z,����Mx_���yu�3%�C�(���>~"�Z+	䧋���퀚��v�
������#�=�5�p	�Q	�6�J(NE-:_=���T����I�~cȤ<<�Yׯ6G��p$�X�Ȍ/0+ pr:`d!=rr�B]|R�8's��4��V�W��+7��r��OU�(��.���%F
[Y��/���Es�x�6���㠾�^��i�,�e�s2���z�2EbP�c8bl�gL�1�`���րڬ��撰����x��_f��ĜV�/��I�_��/�Q���y*ф:�G�¼=�$~&�a�F�-���Y�ɗ��O�W׾�� �)w���=m�O$�D.���n��Bn

̄ܙ 6�U�!Q�t����Nar�)2��b
67�凱A%�68uL�Og#�`�MG�e���@Y�3�������������#gȲ��KޤJ:�,+��� ���`�H˶G>X��佰�mDS>�Dɧ�A*�D�I|��ŝ6���+"q	���f��(�pt`�bV(���h�"~fE�'۶"!�L�E��<��O�����2�ɰ��4dDXX���������v|$�S�u��뻺���S:J���EO�٠,�>H����������_����<.p�?�DU
���S.1X���|���/G�[�*y3gc���&��8EyN�F���{��y� m�K&�ʖ�c�?c~7��K֢�-�rP��^�G�b�Ҙ瓽�zF�����A�a��@��(�,ߍ~Ÿv�h{#aSK9V�#���,��z:`���/���z���8�56A�R6pi��dZ�&mD��<��u#2i��O��x���� lfz����I��MiT�k�����]�O� �7٭y=;Ǖ�:�d�K/SO��@�Q[��P���в�.3�Y3v�>"�ηa�b�� ��%L�?>x�8x0���h7��q��l�]Oh~�z��o�%]ǫV]���F<"���@�W��j�텱��pW	�����L�7-�}�17�8tp�Q�i\� �� �;Mx�Zȝ1F�C�;�ڝ�;CU�D:4c�Us
������V���]�
*�������nyP�K�xjX\�SN�i���;���'Zn �I>W�{�)e���o)�2p��ҦѮNY)q��X9֪�P4�� &�ͥB�l�^��{�R�]�<�Ed�%RFdAf���L���{#��E�����O�w�<��<�bPw��A����V�$z��\cX�7�o���T����E��*F�!���*��?O��Si��.
�5�hj��������n�R�6+���,j�%�x�;��G,��2C���T;(��ڻ��hB������~
^H�Z����F����e���`<
�,��%��#���|/]�ۊ"����w�MF� �T���;n0ٓא8Vk:.+)C�r�/�)�pC���N$��Ȗ�R𮃆�Ǫ.O%U6]i��<��p��uA����X8�6J��>�Ů�A��H�r�z���3����.�F�USΩ�8s����nLm��}�	��P<gWS�`k�eъ�#�Sl0���� �����U�p�ykx�Ќ��t�ڸ���F2�8��n��ŔTNŦ>�I�o�d��~�v�7e��	

�ls�!�:aSش�p�5�ՙ��G��9 �B��L4L猁?�@���偽G$-�߻��G�V[��D�7Ag�|�y�U��"��
Gp���أ'Д��ځ&^ƥ��k��4�B��{�����u~��\HĔޱ-��_�R.�
|Ҩh:B  ,�	�Sug�$��]�����1�*���j�|�]�F��M�Ž]�b��n��|j:������Z��^�,;DY:G=� Ĕ��zd-��?$�]�m�s��R�zf~Ψ�������	!�`��BO�]�|;H\ۧz����.`���P5���k	�pQ��P�[�`�^��(4dP��5NUW(��Gq�o`@c��0)W<9�tß��-h�8d����J9AD,�L�`��@cl�zk��Z�]�e�-WKI� �{�F"j�[����wx`z6��4�$����=��s�~4(���xuW�6�AC3;�a�g�"AiE��������=y�]ip�߭���r�` ��]���3�JX��(�U|��Б����y�L/¤ �.}�{�Nu�����:L�ui��F�1^�v��$֪��KK$������B��$����M�sBP�Id('���@�drb8@]�- "?����܊���(�d:*(��&Ʊ-�/Ib%��{X��Bv�S[^�E�]L���"��P��\�UM3#���5��m�T�[#J;��E)^W��������*q`$�2��F<Ͱ���q�O���*Hp/�� ���"q��즓�~d�P��&L��fTْcV�QV���`�DFO'qY85T����}T�ڞ�Hs`��8� ��_~n�y�o�Q[����<�$�4@|�FE=Q���gsM]
	�Lt�.k7�����Ļ}�|;��
아+��H�Gnw�m7柏NS,��*0���G,1����ʗӏ�q�� �@�lNm��U�)J����M3�����Q��K��h���et�ڗ��/#��)�l���?�5q�,�U�o(�V(�}؞X��y�0 g!˿? �<�d�������٨�@�_��xuSwt[�ݯ�!��=���k��	ʃ�"�����6M�،Z���"�
ȼF�h��0��(Ň���'^_,y^5M&�����٨�C� ���F���P��b���!�G�	���!�(юF�V2hLׂ��^d�G�gz�ځ�7H۬ur k5��K�NF���$��
r��[�ڐ2|	��:�y;���`���F1���.o���:���U�_�		L�3-CQ��:{:IZ�7���?T�6�e$����}���2�s/+�*b�ؘ�5FA�(c��1/m\˾"H�.���/�e��;϶6��$���*�8����N�$#�M��\��֙lR�-u��m֐�D���=�!kZY0ؿ�5�8��+ǖ��$��#I��Z^vn�#`���#��A�0L����d�{���òj�I.�O�Id �K�b�����3d� ��F�|���m@;��:��tj���Ճ"��].�����:
� i^�|�,/�i<2�%�}��V���' ��^�����c�	6�*p���y�$�an�o�ʼ%l֎k��_��}���]fMcE�����Ֆa��a�����������n�v��b0�DՏ�:�4f}W��'��5��xZ�}�h�ϳ	�.j*�\�-�#�'�Ɉ#�Y���jځv���a�+T�n�`ϟ�)��dP�H��~�hrLŜ��m(���@�}�m�rY�?cP����%e�O�� ����8� mB�N�Gc���/V��|Yn���8�����~?�%2���Y��"[��F	�U��Az@��Ș���D�I����d|��=-�F����n�X�ˤi�Q]�E�E�0O�uZ0hTH�<�����ܮ0���&K�ʡ'Ꚏe�Ž�k��Q����&o�~/��SC���<5��Mh^�Xv�����/�i�ZSS�|�r:����w�{v�J$BoП���⯜Y�U����l=��W�!/܉�8��N|�14�hYy��5���jG.��Jj{��}AA��Ͽ�?�[��Q''�U�8�;X���bx���U*��:�,Е���P��B�����24a:�C�s��&yR9��N�Q�<�ƕJ��YVE��]��!����aV侰riï�V���%�u�I^t�,/8b���jR���p+��%�T��Q�h���㉣��sxh��g`��f��H�E�}�ڨ:��p��)�f*�Zs�������\�W�צp���:R_$��	��¢��J���G=�7���uN'Sf�~���*h����zK��Q�6T���n�ⱗ�X�41�+��d��y��L���d��������S�=^v~%�#ı�xTƔb���g�DVC������<���ܾ�MrqxK�w��&����̞����m9��0���?�-�]�.�z#!�4(7t���ۑ�� ���3�*����W�s���f�������GLA%�R�b2Bg���֌�1�����~R��y%�f��ݣ�\��q�&���&�&��<�X�&d&:���g:��x��
��@Eუ�>of[�iQ�����n;޾׆���\2��6��粱�w
�_zQ�7��mN���DQ'ݽD���a��1o��kr�z��$�׸}��3��k�g��/7&�_�D���l�C�s��"�������N$��(E#�_� B�� ��F=܉�^U��R����1+pZ��@24."��#E1 l�b�Z�cS�A9$��3{u��c˟��*c������c�(@a�
7��Qe3ʅ�;dU�X�.ȉ�*.K*׬��yfѵ֨=-�n�
ջ7���+�������/V�&�?�*eO���zA�;B�1���8n�2�$K�yN���!0aT0&.ճ�5Y�q٦�Ôh�m�<R)F�l�;|3+�8H��i�pC���#v���D��ר9�W��y"��ý���c*�'��

���}H�f�3"����MC�A}���t}��1Z��!~h�.�[7�����p���c�|i	�3���9�F*��U��F�v�9�ۦ�~��4����6��߲tBI�&�޹����Y��uq���@��~#6PhYa�s�����6�q֛��j�r��M�p�xp� �Y{�7פ�f�*� Rqsچ�Q3�DA��K�w)�^�>e��Q�T͞@U����&+"���uE��_�<���%��2yݧ~V%��=��9*��;�\<�33.�lĞ>��(k����4:@As)��U�U�ӽTtB���_?�	��s�0s���~v�=s�Ā	b)ǛKR�S$�c�4����ˠ-��5�Y{?����J1���(3���Z�,���P��d�	9��k��h��0R�Xi�y���̌���?5�e���7e�p�r�eK����nփ^N<2��H�^��%�>���~��T���s�����_���tw���pD4�]�a��2���?���ޮ.y��KЛ�,��N�H�M�F���S����,4�N�n�8���D��m ��^�rhzִ�((J�`���䜌�p�(��[ق?̥�����2�t�g��|�n�i&	�}Ѣ��4z�^�-R��#>���Q`���ڀv8;뫷�wak�c�������j�;<�4���H�\�3���g.���k�����H�١��F�FE�a ������pcE<v�/
A� �g*U�7�M������E���2B����x�C��ϰj�����v����Тr��l��#s����
̈́�ZR �E�b�g�Y7?b���f�JKAg�V7H_�o�ݐ����a:���2.����ǡ���sQb��@�<�1��I�c����w�_&O-a6���cƀ��Y�E�������.�ny0A�Rj:��?"x��}ĠsH��D@V�]�϶�:<�H?j�`�>D0�9��yR=T�
���?ذS���H.&B�]%E��D頡���F��*A9����Y;�t��{�kǇ�Z����G�{�T8�(�=r�����) �e۹:fR�7+��f���)��3��R�:�]��gC�:��?a�A���k�N��5W�ag�L ꯧ