��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��-P�${GIW�?j��g�E�ضsN�ˊR����MH���jz�
P��`�سm�����0�N������S}�0��yt��q�����Gx�kM�U:�Ř�ɳ�,t�Үo$2̏98��bة��=�j��M[����nr�!>>�����N��⊬,�fy4F&��6'��*:ˮ��<t�MmpdI'�.���%.�B��b�˘�[�������se�й�����Glױ�>k��%���S_���F�7I�ӊ�uJY�o�~��
0y9=iX7(�w�Z����@L^�������4�(�ƀ���! �I��nZ?S������1Ș|��9�M�@� ���j���,Ĩ��crP������r�QZ"�ck�U��5��y�DKj�?#��r�e�6��@�(�t��h���U|�{op�pve�+4���zQ�>�'q�V��s`#��S��RQ=�W�&Ը�*�H���<���F�\j�B�'qڰv��Y���%ߘ��[@S/�Y��("=��y���c��e���o��2J(������U�^��a����_���=C�[27֨�R��|� �\�O�l�od
�_7oЎ)�sox��Y,���*�p�Q��~������o�������(��Z�eα�W�Zj@�<J&<<�s�nOEewR�a�=�b���\C>]I��;kW����G��D%��\.Z#�t�1���ioRD^gؘk	��v�wOfύ���l ���]�nO�JI��_Xf�l�'�C��_Mw�Yv������yE�
���\��5->A�E����%~�Q��B*���.��|��V����F_�׌H���A��S�g蘊s��nx�l(�<�"��S �i�P�����{йB���@GY�I[9Ӷk�/L�2d�țs.���Fm���x|����ŵ�6�Ų[`nʫ�b>�ʨp!�[���L��A�,m�x�Q�1M�w-��V��|�N�l� Oʩ���ʝ�������b�FUv���?�����s�f�)��%�Zg���;�R��\�L[�jq����M?�}��C��aP����X{юu�
��֋�Z�`Œ��ܮ����X�C��kS~q�A�}��O|��������s��������� �:ۋrOhg �Suj�;��j3}	c��ⲺY{KrɉEУ�.�ei4%���v�@zs�Q��26�'J�_����y .��J�%F�D��X�z�Ҡv!��2F�4ZV��M���ۆ�[�R�8Ɍ=��Ns!@��3�Qb�bg2�g}j/�'��%}M��H�9?'�tZkX;�$K��s����\�`�@ݼH5dk�]�݊���7�sm�܈�
�� y�Ҿ$V	\H�syK����w�Yz�:B��]�FCG���q�����"�%/�9}p��M����h�_üa�V}���hH;���JNv�{D������#K���qРzE�!�X�>��#�$�֭�ɟ$EF%��" ޏ�9��B��_W�"gI(�M*�sB���b�,��#�i�-F��Ń�E���5<k���~O�v�S�Q���A����9e������������/�4�$��� �yW���>�Ș�i� e��H���|�0k%F�����2sf:��x�ǁ͵��Ĕ}��A�LF����C���p:^�u�Xԃ�X����ީ���	�?��F�5g̪�
��/��[�H��{ 86j�xѼ��l J^J��Ԣ�EB�����]$O �\���*ґ�Ϛt�GQyD^ǌ����p!��.��D�M�/�Y\�ꩢ���y�n��h�0�5�w5s=oض����`�*��
<K���$5Y������VjP���'�J�-�	�3�:��a���8�Bƅ�0L���������$����"n9�O1ͰC���x�d��ŧD�E�����K�lbؚ��;�C�~�^\S�;>��Js�E_�?7L�����i-xy"�����C���������$��M�ph�+nֱCޣ���]~o��ֈ��v�u�]U�X����i�tB�W��$C]5�GI�x��q�?9�Z�:Ě�6�q�w��\����4o�3�,:�;���2?��B5/�9�/%R���-��{�̌�Kł�Ko����Bv��Ř��x�,����l��jˀ)�)��p�F�(�j�ޔq�ΨdBmrV�bc�Kݼq͕63	m��,�|$�.��9��}�����V\ޥ+��"�R�=y��cT���ַ��b��K�a��wP���|�G�j�k��%+���$G�N��' H*�@g�?�������=�b���S�P��^��m��P8t7��b�ȸd	r���/}�΁��匴����߱C�;2s���Bd��d�h��8�����@��Uj[�|	9���+Ӳ�]��� 2�{d̆'ԟ��ʼ��|2g�#\�^��SA
70R`��f�>�ìk/L�-�A��aM� ~�<<o��`,����4@�Eľf&Eɶ2����H.����������lf��}��~��`�|*3?B�%MeV�`lsZ��KܝC�4q;��݂�\@y�{�dsV�[n���.ۊ
�3�bf����W�Kl�����2nf-j�w��d%07ו蝇5�2s��s�c��Jōr��m���sx�R@�2���5��Lk$�A���л����dew��F�qn��(��K���:DcQT��	a2�N���@]v�E5mǦ��*��J�:zO,8)����3�CY�B��,��'��Ql��
��$�H����,Z[��ߨYm�����K(�$&Y{��j�n���p�Ȏ(����+�	yMg��"�~���ޖ�Z>��l l(45�M��t�-5�/��{���L�俛�8�  ��#��)0����e}���%�z����]��0EȚ̀����4S8^T�����nF��l�=,�nZ!�A��:��f��@��N��D��5TJ���')0�~QY&�����ie�D�]d��{�D�~�g�ڋ`�7kv㑯eB�*y"�u��%,$T0��x�\���otC�{U�䡃;c�^����ٴ>�}����B!�q@�甾����}�p��0�������1��)���'���Z�,�R�!�W:='G?K0Q�2��Gj)���D�z�w�4�h2��։����yV�So�An�Ə�L�G|H��5{�&�2�P��ch �.�a�[9��C�J|Xa�ޜJ�C�eb�N�w��Q%�5-�Z�މ�rϞ�sT�����ޡ'������@`�fC�J����++l��P̞�9���g�	������"�K��sDhm�u|�Y,c�=���@$��܉���l�?����xsv�/����L�Pv�H�OH � a*���S� �8�Δy^F��=���	*0�rx$��|�f��	F���SL>Z��]�wa�}G���v��8Wc�D�p������|q��k^n]�n�F��"��o�-�?EYW�.����dH�Oq��x�(���r���Q�Ԉ�AGE7��R�u\�3{ �D
��AA��,=H�(��� L�Ű�IߋՈ�<(��$&�8�I� �oڢ�� ��>spz~�s,(@u�g$������<�R�#GX��W��p��*���׼�K��.ҋ؛���om��ݛ|%��!(�w���{4r�m�b6Q6.w{l���G5Xv���$��g��5��=K�Gh���Q��K���ػ���ÈÅ��÷��f�� ag
��%Ơ�Ք`ylX�*�Z!��0��ό��N�q�q�y
Xz�ay�6��'�n��a�����B� �	
 ��l	PAk}s[���,>}77+�j��N�G�d+�7w��LO;�#���	���ޘ��y�X}K��Ĉ��=�\�V��������y�'�U>��5_جc��+<�����d;���8C�s�� DT�e_]���I9�xߎ�Q��Hz�JI��Q����$F��+/@�=�h�&��6�L��ysr�tW�a)s3�h�1ϙe��z��)��0#k�~�kS�y�ӿ��e�R��%��Dx�A�?6e3Æ|�j�==�L���"�w�~��Q.���)��(O����,�e�N$�m���f��k|�u��O��2b�^i����ڶ�M��L�g��E�@�~��2�^>�H�K�	�E3�w#J��OuB���g��FCT�V�	���]Ae�OP@�q$/Ϋ}��g�6�t;��2֒�Y��(?��r����1H����렷�:%�tw<�sዂ�LͦT)�ӯ�Yn�uZ�y.Pp�Otn���ΖB�-��k���͛d;���Ԩ�J�����|�֏8V�S�{H:�qf<��k�z܄�޲w�f���|�ӣh�T
�<(��	������P�=�=�o���k�G)�wI+Ld#��Ԗ��F�]l�T-'�ކ��/�C%���T�[V�r�+�'(lѳ�g{�Mcb��,R>���s� �[q�C;��DIR�d]z���D�Ej�A#���!��5#��0���Z݇�J�*	ќ��+�O�Nr���/AE��(��j]jA�����d��}�5���������B�P|��է(����O�ҭ���M.��Y7�����¹�YIQ>�-��-����hJ�Z�|���g��5����]�W)�w��8a���dN2�5
�
6G��[�.Gsפ��\mxrՙ_j�1>�q�ۍi���2LV@lrZtw�}*���,!� �'��ŻC�?x��$9�'8_%9k3#\�z�u=X�aZ�"<�u��>���K�ҁ)��2Ԫ�O��s��\c3�5�P~���E�8Hfӑ{bk�)���Βk�}��*`_gF�n����.X�F�ǀ��A�s�AcCGZ�}މ|�YS�;��^������K]	Æ�?�򣉓�*j9��;k{!���i��x��W^ܴ����t���N����j�{;���+!BSv�;�^��p��0G��}Sҽ�{׹��'����&,h��p����Rh��p�ϟ�2.ѕX������bQ��4��x��_F�Z��n��n�ľ�B�������X	�҅��Q�yQ(L�p��M�!<��m;U�9�|���N�!��J�Z��a{8�t*���`	�i_t�wƖ,$�sK�uZ�{�GV�#<Kc�9��}��!�D�re�2ȋ�tI�'b9�P���f�����̓?�V�h�d���A�Q:�|�y����@fiޮ`	����r8%�J����1� D�"el��U�(#n�͂E�9mk����}i��g���F� ����q�M�c!&�xs�U}�P�kRq�|�󜦡>�9�:&~�Edv7�s~e|�-�����i��Wz򈲅�kݦ��Qӕ:j�8�X8.?�;q�eK4������e]C�P���I�����\<�y�;ު����ཀ���XlԈ��!J�pNR��h.�����0o��wf�FW}{���&��E9��W=A���T����6}�X��٨�����Έ���;�2�ۏ>����<�P�i�A\k����>%
m[�z(��Q�q�k����f�Fu��%���s�vI�}HwXfjL	���x�E�{@K���*/�5ؓ9h��k���Уmt뫜#|�hI�x��ۜ��p���I0�J̈�hV��>vD�eXT}����è��5p����∝��C�*��ﶊe��)�nql��\Ұ��{��z�� ��_́vj��J2,�-���{^Dݓ' '�0p�����`|��?AuޝY�d�����w��9��l�=!�)C��R�6v��K;�a�>�ӏ�d�׉���/�)�K\���M�5%N��D�_)"�7V��K��՚)�!'���X�tBj���0���`��]ikA�w38�(�UW���U�W���`A�����B�t.�i��2CNx[�ż�;;���}=B�V8d���Y?�m���l%^.n,���	b��5�Ϸ+�mK�b�wڬ��~��!C�Z�SF��iV+�B����H��=0k�@����k�m�����6�����$�釩�����e��{ɘkX����B[�2�l����-� ,�]�W�8YZ�W�1e����5��d�>1���m�>j�˔p�@������ϱ�V���k~�׆��j�x�}`��Q2D~?��#U��Ҁ�K(S��m���c�6u(׆��������7�,;4��W�và�~_�C�q��`�J��W|�E�;i\���T�w/f�k��o'n�(f?]]�i�lz�cyؖd1�,o�S�q���OoL/����ʆ,���;���h2Ҧ"T�x49B'����
X�RA������{]�q��:���o��A���T3	�Q�#'K���T:�t��G��I�vڧ�o,�p��3e�w)_vD'�!����S'A�t'�W�E�V���c^'��noӺb.����4a��G߁"�Jog�#6�������\�7�l���2��r��[Y�/��XC�9�|0�įQ6�0��B�3�s�3jH7��w]��$�;6�l����H���y�FW��ɚ@�|cq��vU�{�	�+�i�k+����t�gh��e�Q��d1ڴ�{k�܍�|��`�X(����^��4���fڿ�Ѿ�����)]�a��s�!F��.��\��{��>��/�ѹ��k^ ����J�(�jJ��y��K��H�|r�K6"N�g��[)� �Ȏ���V��#8���6fk� o��wb�s��+<ɿB�(b��U؃�攚4U�n���`�p���Nfƥ�ڱS�d��c����kW>)�<�� �I���Ťi���Vgp�Z$�+����E�A�5��F^���O[1�2��')�U����劀�/	��.՝^����0�27��+���<��)mс>70��7�V�[��i�Zx��|����^2��G:��	[��b8����bn�&��=4n��e�ׅ"��c��%���6�;�z��E*u�5�QY�����[����\p�8T��#�«���`s�#t��	�q%��PIl�W�Q����y�c�a�6�#�P:4����C�=@��cAU}]��F,A��`�ˎy11F/lu&>�����d'�5�p����\>P�:m����=R�n�e�����������s?~H	e�˟��lB��I��V}jN�fE�y9|`��7\(��1ʲN��>���g�(�_&ֹ�j}��l���Y�N��b ��W�ڛ�����zS��8�XR���߲S���Ϲ�S�K�o��ͺ�yi5}ȊeF����BE�*/jqO8���g�;��5��K�V��)����m&p"�I9c}������s'a47Q�K�x�}.q�${�(j1�:�[�������P�N��t�!�Ly�9�����+_���1�i�5�opM 3����kn��9o\�_ۥ5�&&x��d��ѳNϤ|��K��*CUp��LGZr�� ^�t���M^��7��| �#�͊U��$Z�PȴAI0&
t.�}�@�};�AXJ�f|�g�R�^�a��VKsg���C�n�U[��y�S����U_��IU0N�H3|��J����[V_'��U��:���
qP�^��`������^�����g���J���޲���F�
3Qmd�0�Z@㡄X�|��}K��Nw�R���Z��N�P���Izh�`���"��Z��fs{�XPi����f��u��:�J�*��T��y`s���3�Z��v�}���~�Pr�mf�2�@q��nOb7S�]rx��U����.-}CjE��X����M1�$exF���w�[7�d�k6��C 1G���zԕ!�|h�A�W���L����-\Ey�Гn.�4k��s�g̀�u 2�	�a��|mKC�vD.!������T�A�H\*iw���ϥW"y��ݻl<����
q�sqG�nX4��"�W�rKc���s!�ɩ����K� ���E�4��&*�o��q,��^�5�8�+���l���^*s.��k2&��r/���wZ���n{�/;(4�ۋ*͋*M:��6e�>�3LhD���4��oR����1^m�&}�����f��/F���/M(�|H�u:��5A4-7�y��-��sd�r_����Ws Ӕ��X:"+*�������&:"=�EZd�� ��M��y{uo���"Pct�C��쎭�l�8�P�����}T�q�_�~�T��缄���_�a�n�2L�
oY�D
�֣fZK���Q��.mO���y�-$�G�t�F|�k�a�6����΀�}䛭�[*��� IdO�~{���m���u�32H�%��w�Y|^�؜��g|0^;xg�Y� ����ᙔ�A��/���&cO�?Ͷ&�!�&1������^���_τ^���`�P��-����w���@I���+[����,�����a_،�J`��v�񉅟qj�P�d�o��4��ů�a�I��-=lK�D�ѷ��vl��Q,2��qLy�l�"�$oQ4H ޞ������VZ���p�Rt[��+���jʻ�6#�T
`K��f�f�+C�:RxN�%�J��膓o��Ǌ5�'\[^����N�@ɡX�6)-o
q�kl��/�T�{?��f�l��m�n$%
�~����+C�s�N:�h�$�`"'D5-��O��$ �Qvq��HZ�y�Qߺ>�m~��6v��Bn�^u/�@c������G��ȸ