��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z��i�hW��1�%:~c�"N��˹�wG��5�H�
�P+����ֈ��Ŀq��5�d�TDe&2��xS�\"� �#D�+N�[�ZU'6��s�ON��� d+Һ�޵\�"�J�б�tz�����vk3�^M��q�T��Pg�=;|3ktB)�����H���x�-��Y������X��@kkHy`�x�N��3��9B��''�J������'�� �>X��;�;����J �6�{˯v�<?�<����B��P��N�E+orİ�B��h�`�2�-�K���z�H�l�E�	�7�H��MT�=6}��J]|h�#�����1���n�g��E���1� ����<@���k�᮱	��|#~��~Հ��H��< "�7��'�t�Ћo���:Y�C\-�<��C�ee�ë�#��ȽOY |�|*����=�H#�#���G�h'�/͢v�:���WL�t���J:�))	�v! :$�\�1,<�n���H�M��0��^���XM(����6��@�y�,�����$%��>�1����#�Rk8M� �F�G��iQӴo�����}kףl��r��oo�#��R����4�fB�@Q�Q���	�ϐ���P֑�_�2@@�b��NaV��NkW!6B���匤(�ц�%����>�O�H��B�P�a�Oc��a;�����^K�E1��������;��!�e9�7ڐE����p��,�2��#2�Щ��)�U2��Mv��ʠa@F�^?��!��d�sN�'�� �t����X!�fl�>���Zd���#ur{���gߩ��?
�i��������Ƣ������2%\AzT��bMW[7`�.D�Q�3��@R8à�-�b��Iz(h��|@jrQ��ƻ��0B���������m؁�_��~>s�ښ�;Ts+i���3���"���y�|�*�t���?��\	�We��&�
���=��YF��\�AE�68;h��.�"�ku��z}ε�'�>r~g�T�wx	8���|�@@ ˸��?�x��"���M���A��fgq�mR���@�6r@8��Qk����l��4���'�v���fw>�����o@�%vS�ū��{tO`�J�0B@4ՄXx���A����΁qť*��ky���2������ٸA�^�CJ�ѩZ�h�`~Q���j�ę�on�a.�A%�]�}���#�  ����p,K'���`s9:]�nzT�%�38�&h�Q� �;����T��7:�Z��+m���`��8Z��I��
�xab�{҃e�W1j�Q(!�J~@>�%aj���� ��j3g:�^[�����O/�\��h�^J<<tޥ�fu\U��[��lX�JI	��I�P$x�5�����N�20[9�S鱻�������FE�,���ɯ�O�&�s�q��Kk.��^)�-Ē�5|G����|�)֧0�ce�j���$@<�lρ��ڽ�A�N@��V�զ���]L�񙲀�4���k�v 
��,�Y�~p�-�y~~jw�@qFO^LtS#�a�%���U��w	�+�c��3$��ש�����T�[A��e|�pã�6R<xĿ!�R�j�T�ʟ�6rc*�N�׶�@zM�2�E�ۋh���GJ�&�K!�)�CW
�ʺ5�0L�O�@N���c{� �yz�\�UQ�աz�S�s`Cl.�?wr%��]@�2����D��)]Cp�ŏ�J]��Œ�*1��ЕҖͫѼ ��.�CQ̨7��O
������..���J|�%��#x��x>�;�r6 �җ�����k�j��M�p&:��C�U��8[�0�RM�
��Y����ŧ׻I�5̛��h!���
���ڶ��?޶��a� �(]�L��4�_%���Bwy�Ɗ�9��v�ND�9�Ư�v�h����^�+��}�u:8^V�G_V�74[\u���2�y={%�7ya� .�j��v^9\�Ɂ�ؠn;�$�(ek.Bo=p�`�yQl�Y걳F���>��E�r�����<�q�z�w����,��s]c�7(���V͕S��	>G���p� �}fs�*T�>��3U�����-aI]]�	!9�kTδP������3��������K�х�!���5��;�1R��	CG�c����������cH��
�@ ��	� ��{/{�m��ָe����9�>?7^��Z�L	�(6Y[(�X*y�H�����p��уrxf��l���|	�3F�0�1��G�"�:��4��%:�NTs<ƨ�zE�v���"��u��·�o"�m�u�����2�%�Z1� �4����R��(! S��&�+��!0B3��������ngo���!	�)�چ�3Ȧ�,��\�m�l���uƸ5ya��b�����5��G��F%)��.r80�	����d��'��6���g�~�2�U���c����΂�Y�4���2FG���ֶ�����*h�V]
}%����g*2w�����Gƙ��6�j���j��M�[j�C�,����_dUt��	�����b�D����mO�?����Z�J;tF�|l5�8o�l��o拀Z>j�����Y*�F���&�7�����|�1��}�T栥z2��ݮrJ���� 2����/k�[ث8(q!!�=�n����T�T���Ԅ�y���,p��(�g&Vc���1�_�^yy#�O��@iG��c�^,r&�B�$8/q2}J9���o@	:�޿F�+����5yN�>��Y&۬8��1�mZ� ��m)6��EPc=�r�'�c�ws4T�,��=�7��;u�%�N���-�'H@*2<8	���)�P��!�SW�Dh��qP#��55��|�;��6��=d~��e)�<u1h��B���Π��}�NɿZ��i��h_�4�1"I��n�c<��i��;����7ݚ�1L���Ѻ�=优� ���ln��a���"q�_�_C��W�S{������xj��-�y���8'	��������V	un7sFI�gu�͑��0�.���)����'��{3'�A�� ��C#�ڶ�ׇ�w�pJ.��%��%}�qc�:���.����V�:'ª�1T�e�� �6���gmX�k٣}��H����&Gbj/�/��Hr<���w��������o>�0�%�Uon�Y߯)	��qd��I'�oM���쎫�;l/�
C�߳��N:�צ�4��!�$7x�����;t�J]�nT�L�`-U�apa��ZP(�(����M��_ 4��M7��fpH]���O�(��@[mq?�U�p]�q�׮l,�%�IL1��^8�VT�(US[ ���jN���'��`�5��-��"����0������Jd`i{���d~"���7xOɳrH&��jtj$��W*�;��C�>�q���U��aϾ�4��{����c)�P[�eBE٧%�i�"�� �aq�R��IMق�qH��Ol6�S8a4��&�Ѳu94=����X3]���$uf�}Uf�t�pZT�0��)��g���h~[�*u��X����q��Q��@���V�ئ�^����d�����a� ^���;y����SI�jH��H�Z6�0�~�mb���D��m8��Ww�-
:^�$�s���q��8��[�aco�ܷ���NiЇ��6�h9t9��4�SȰ�*>�l�����U��0�qi6�օQ������"���[VX���h���P-V)WQ�\�d$c1��=��Y&h4'���)�l���]0��v�¡!$���7c<��i��\ ��`�fU@�h��{�q.�<�
�6;��"����x^�N�n���3qp��S(���F�NE�)�9��@�1ҴM�?&�	#�V�|]Q�����lJ���YH;�����)�X>V��BDz�i��:�%Zg\�-�l'�)���*�Tum�s�\=e��"�U)S?,L ����fx�c2-�hJ��ם�	D������N ep�RA�#�ifX'����Ma������j���m2��A�	Z�'�ײ|"9����r��v�} :�}��X�w�Ώ�ʹ˜�X�A2;��9����NK�	Y�3d��zJ��Ϥ��1����*�[�m%F��J@���[�{�����֘eu�l �r<���FO0���D����i�n���=���)u���<�}��-�@�K�E�s�A.�x!�{������|^,��Xʹ�^N�m��R��7H��d��[����(.ѲdP�)�(l���uٙ{*�mm�K�l��&贊���h��;Шq2�|�y�a�|P64��،r�-ʎ��aP���T�����]���#y�D����)P>��N�Qy��a3{�ɚQ��M���\F�+#������ի�3Y�'�E#;Н>M����-O{��~��>��uxœJp��zV��Od�y[i�+c6g��>�isC�@ن�e���:�i���-Ǯ ���p�IM�J�C�9ފ@-�'5�dh�%w�UxhW��V]�e���\��|��/�ы����hȲ�����q��\q_J{C�;zȴT������0bJf��MWzp����o�e��Y'P���Z���U�'�DlZ�SP5��}�� �Qb⽂�V�4�<��s;��_e���f|���
���G�勑��]��0�û�����}�m��8�~F��$�����V��0�V�L���Ⱥ��h��R��U�ș2B3��9r��k_}tK;�����{fu)��3���7�e����7���64�m�JW���� NjqUM�?.%h>'�C���9��PX�u'��W���z����4�e:�)�Q�v	��a������"#A�0��,_$3�$�/�g�!oď*�B��n]W ��M�� �����樇�쫑��s�V�A�T'dWB!�*<
iܕ3�X�����D�f2�6)Y6`k��[�cʒ�k�N�Yu��k!$ٗ��}��A�|�X���Z#�O����1YC�"桠�q>�y�~������BPq�j/�h�2j�gLo�L��������+�z�7Dwy��H��s�,���P�Y)?��}�P�F/�C6��l�j�)����l��%�A�:pVp�A��L)VH8ێ�h"��m1���i�/�����0��<�@Q3�e��a]�ˮ(�T��EV`b�u��m~�'jwLos�z�O�E�L�4{{�v��%�Y͗2S��f����"���$B�3aW��bٳ��|�_3,`�x��\C���F�ѝV�і��y7"ʀ�u�~AH
�����W`d�2ק����+&�/Y;%"$�cFM�l�z/��㨈��he�=���R��{�Y��mG�D��b���T�Q�b�?1>��M�����155�IoA�ͳ����z��������/=�����̠�e����r��lRF�қE�_e��v��яMC]!Mkm�Ah��NJ}�4g���g?G�_�9g�[v7Ө3s���e��-��B�����CL�J)p��GO������ʆ���&���2��Їm��f��3�GL�TE��L��$&0�����9Hf�������~&|���ߞ��8�,��Q1�.~�E�чg"\�}󇸏���<<�N����A�|iK���< �5��/}�s�&��u���N]W�����D�	�^�$=���/����蒯g�޻ ��T�T����J
P�<��}V`�B١�]7���,������3Yr�*���GY^�lڱ��v�=�o��������oK O�猇�l���k2�j��V&-�Z�7�`�A��ȟܐ�ƃ�(鞆�t�&�P��?h?6[�iކ\�)�J���bm�f����p���3���;�����R	j]B�b���rQ��>���h��+}@�\$���3Eԥ<�l��20p�&��D6��{2�qS�Gv=�Y�R~�^,,�xm8�$6A:�j���7m�pgUWZ)(t�.��$Ɠ�R���Q"r��*�y�4����~.F B���������CP�N*�:��S��\])��<���*O��{�N�T��Yw4����LpKB$)�\�6E���Cd>��|���e��%M^6{��v�<@��<��C?H�/V�(C7��]{G���9BeOmK*��]�K��}C�>���s7g�M/L0�b�����ᫎ)z�2�m��=F�#Q�k��5�M��y�l��5�9
�N��#�1��&�kKs����c���'P\��jx6��vj�+��_rX�U�{1�Y�ˡGa�@� }^�v����n�������I���T����EZP��m��뢆(2?>���+Fp��p���k�#@�e�IM����y�0=ò;S������� ~�ȦK<ӫ�^+O�JFhц��v��� |�3��gu��6��<+` �ˁY��l�=p.��W�6Fpp�2�<bD��@��s�CZ
��r�W�Շ���W���zy�V��<O�1;��2��e��A�]��v�N�}��:��&9�BϹ�rL\�\�YbO2��ND2�b���qgzB�yIڵ~;� ��ի��|x���Hl�A�j�'�����(�Qj:gy��/�qF�#��R(9�lO�kǷ��:ؓJe[-�Dt�p�!4�$%)̸=ca<��ݖ��	(�N���=������\��V�@}F�%%ý���$:��
+Wk���t=�F��sj��1�Je/.�ch��q�p��46�$�.�+�qZ�DXc���kQ|h�kp�?[H&ݭ tԀԔ�j�t~R����P��k2�F��򮶶�B�;�a�����N��cN�V0�	�~��0�eE��B8AgNݨ����A=�+s�FS��`G�o���B'�6i��cz!�f���.gT�ΈQ'�9p��O��|���M�~��S _z�5��H76�9�T�Vr��9)�'m#��!Ӥ9�ԥ-�����c	��]\,���H�h��Σ�����^u��9�<��&�i�ʺH��	��o%��ʖ��=�-��G`�l*r}Z8�h�%׻�	���K?�kr(�kоc���q¡o�
���Oi43�VQXH���6Twǧ��ɕlН�1�Ӊ&�?s��(_2b��d@��b��Ӧ�;|�4Ƴry('�~e�q�>��i���ma{�q��#���� >CK�Һ{0�u�ō�xĕ���j�RNރ�bL�}�1o�c,H;�i�r�cJ7g�ݍ�K��������d��^l�Y���1�'fe$ �qwϠ �_��l�l=q�>.�t��&̖dq�Y���W�������'�p��������A{�jDَ���*Ց�Ĩ�V�B����&��Y C:���N�\��7JޖP�\-��r�1I��� _��\<���?��V��h(N��(�������D�MD�� ͆)��F��w����j+v����XnF�F�e9�=��Q[<:@�=S����M����]��\�K���D��[&�����Y�{%I�S �|�X��3d(�-,�eo4���>��F� ���^��h�/h�P�\�����ڃ���oCV��,�ďtکs�ζ��	���a7��~� `�P�Ի�i���L��Z�k��=%