��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�j�U";��߽��$�[��4R��$
����e����?�Q�Cg�7S{7ف�?>�N� {�:���x���j̽B�����-�P��?ʰQ������p��r�O�_\f@��=�<"Iyܞ$�Pxҳ}�dmSsЅ�����,�&�'�����'n`��X��)���S��*�_���.�<׺~s0�����<u�T^�ᘭp�P��WȺ!'�l��"���O* ���d����"*>���r��>R�Q+u����S�G�0��K��П�q����:P�:ײj���k^��%#9�m�c��Q�_���,��-@l��KZ�d�o3>7A����/ ��yp:�oV7ŨT�-��F�0])I��&�+nN��9y`H�]�!�� e1ɞ�M�p�3���u��LM�d"sJAU�7�l�S�%o^��������Op���y�B��٤�*�tV��c{:�NC�
8�	�*����a���L�1��d�]���{vm4�θ庩�/N�
��BN��*�`;���������%V�k�<0��Z�i��zo� )���tn�̅l��)i�o��@uoL&Ƙ�:�=-r�%�|��9y���<��ert�i�A�[��5������Ʌe�t�M�i��K�^���遆����gT�Z���1�h�B-�Y_���/D~�� ���'�H��e>I'�6e�1��{χ������rW��,[�FCl���n(I�=��v^�ME���g�h
�UhO9���-L(��Z� ]-��4C�����H�8��~�{��]+H��r��.#i������k���p��);���)��ҭ�U�� ?�6p:�k��_�߭@v0/:�s�o�"ҧ���h�yz�i��L�-y��)]��6�	,L���K���&�׋XG�+�*� �l�ҏ'���$�ݘ�]6��`Z��0^R&|E��?B�A�-�͞��#�4���0d�$�26s?�>cl�A�1V�"��DI�iS���ʼ��Yn{��ᒛ-Gg�h�:�n(��wlS�v���7�h�ރ�b˄ê���d�=�~a��=*�m��o��JM����S19���xT�ï����#�}�����0�$:qL�o杆{�&�LSE&��6�v��"���",#���q}emۈ(:���2ғ�r�e0��(���?Z*K�!��Ú8G�or�w�M|�?S�~���xip(�Ul��Ņ5��@�[@����M��V}��	��ٵ���c�Tb@!u��22{�o�<0��hE���Q_K.�4� �M�h-��M7O %�6�@���m%lO
�tY�J����)Ҟ���Н�[���şo����/���[�@tzڬ�-�i<B��T=����ݕ����E&�F5�\��<���2E7�d/������Sjo˨Bz�� �v#�	N�tSr�E�B�����^������i,c�؟�$� 7��G
ܕ�}`V^�n�8���oc�w����
���Cɷ�!�y`m�&�uż;')�ɉ�hf��;��O~ڰ\KK���T;������#��oN�-�ڡ"���W��׼�Y�w�d11�H|ж����*�$�VD�m�$"����AJ�=h�;L�8	R�x<�C�N��#���]לn����5j6q� ����|�NUa��д��O���r�:֪�$k�|�^��&��|Ri�J
ZNHJm��y;9BӞm����.�����	��)��yG'��9uk�lH�|%�+����'!���������P07/�wHPD-X냋)�S�C?2 	4�IIs���:�������{�=�x����<= ���z%[ҩ�N �Ҙg>M�Do��RT�?}����a<����C�a6�a0l�8T?�n��4=H�s'��O���A��K�TLK��Iʚ�(�-_��@��#�ǯ�/2�6�#��^��N:Ą��^�B�`��X�Uf�o�@��an�������!~�,����Z;�lúZKjz��h$��G��^į�5Duǿ!�p�!��|#�A��u�#=t�dմ�C��"�(f��X^�:�hl����υ�@C��Iĝ�ln��9��� ��BQGpgX��U'�6�2��'��P�VBm��M��\�J&�C{ģ(Űb:�2�K���o;��س5��u�Y'�D#��K�{-g~	<��К���m;ߵ!]y)z�:����l�*�f�i�?�PP�/-�G����������=Q�XOQ�O���%~�������T��>7q!����2`����b�a��Cπ�ښRpKvn�S��0��]'��@O���AL���9+nᝡ��߉C��)ƽ�SG��G��J<�>��iZ��Ad�B�:���=�"�/�ۭ�W���8�����="=� s]�H�����@U�}:Ԩ��h��lX���]f��Y!��?'�^5��Ōpkl��� DU�:_��d�#e(O+K�/ثCO��x�qN������~�ӽ��ŝ�N��Dr�י�-Խ�>A�%X�P3(����%
��/r _Ԧ��Sw�S���t���.�M�`6|jӬ�Bm1��G��Ox*T��e���]!�c��!b��S_�]TZc�@	�{˂<l��T����� C�sc,�U���Q���i^{��"�N"֤|�'�A���h���S���C�F�s�%���^T
���3I�tC1��7P�mO�"�)#Sx�����	����N����t�/��]�,wW'<
kL���M�}]����c����C���o������
����g[�O���T�J�S�,��T��bu5��/9yɶ�!}��/[��%#[�,�)�iv���,�bRꎡ=���Jt���G�F~N�G,�	��e����n&4�"v��f0w���L����Ju�0@7=1��m}���"��Su�u������b
^��9������6J�>�Lm�=J���q����U>��'�I��֐��|�����%А��94�VF�b�ʎ�g�م�*�����꛳���,�%zKW�����j5�dHq3R�1`���	G!��*�BS���Z�q�}������4���Į�4Gr�����UѩQ>�C�3[����P��j`�