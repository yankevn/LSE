��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�U�|�=?�r�� ��>&�G�K�����������݋h�	��� F<�n�BA4��!>mq})�C��De%3,ȅ�(�e�:�z	_��-Ӵaz�4J�D�a����6�� �w���
��`^H�oF���{J�9����5���q�*�.m��������*n���?��%3��/�*�X�+�a�\d�ԩSU��s����F�sT�kI'`�.�C՞D��!"%�!yB��3����qy:E ��ӸJ�Pf>]S�O��x�]�1,p��(aT�,Ȉ^���ݿz��`�x	�E�@����vjf��P�0#�Jb_�*P|����py�=$C_ȵ�Kc'�\)p�C}���!�k@������j���E�P>Ixq�L?��1 �D��!��79��(�:�e\�`zI���� ��@�����wbqk���܏�yA�c���ެ�@A�X�/	֍����bw��埖�i�ޕ����D��E���^�ˉP�^�\h�*�� ����T�v�Q�d �*��˵����z̷ಯr]X��H�%�k���Dr�����.`�\�Sc��N�j��9�)Ũ�:��d�u�ES�4�R���m4i������?􀼊����۱�����Ƚ�f�X��m�PW��g�H����}�^=a�A|^� }\<���f;�F��R�t<_߄�5��/u��"TαJN1k݋+�������#Wߙ36��1�~<k��v�b"ٷDPh.������5W���+b.%�d;�젇޿�6�� %�D!'9��	
,v�iF.mO����ߝ,�U��E䦼M�ן���?�6����>������({���G3|��u��Z�H\��cd2J
Gj��U;Uf�c�m��O�\��eٱ𕉞������,ܦH~��2�`�b���e����7H�҉�S0�=^��iS�6����#0+���J>�f�� 6H�Uq1��p'9��=��%����a��m>q����C�m���Ǻ�u]%�.E��vN���L�!�S���q]
�B��/}|��`c�y���qb�������+`�C6�.�5�r�t�OSeH,���!?l3��9XD9j�n������w���R�O�)�Q�c���!�R��xE<��F�8�&Gx@�{#!$�}Z�_+��V�;tt{_K�_
ÿ*S0��i�_�,�h�4���A�#֧���AA�rQiHd'�����̀�Ou�7J�+��]�#�\�^S�Q��_c�94�v�<�^����VԈ ȩ�A���"za�Ͷ���)-:J~p�Z��Nq+1��.9��ŝ�Ay.ja�:4u�U5�B�U��.�yKa�����N�&�@=N���@d�D\J��w$��e�Ϙ�1$k������"�_��pA]�B:A���c~H�D7����������t�8��Fٌ�aR���G��?�'B�!�^Y���nL �?\3黎���G�Ʈ^�X­�UV��%S��ז�H����}��B�m1�GM܂�������֥7��5H�IK�!Q�k�-�*N�P;Һ;����4������{���O�?���=e2�6}�S�	'5�R̻��+��]�E�n FHt�b�=)K��`b� �?%l�Hd₤g,��SmS���4h �P 0��q�y�'�� ��ˇ�6ǣ�������kC�~�������yR�ω�2'�p�hn��L�`��K��(�st���V�%6��c�?7��dQ�I�i���azx|�9��kgY�)w�+G���vf���h	�tD���� CXCR;]����	Y�<B^����d[W��vz3��K'��u�v��^8S5�{YZ�T�+!]����>a���T�m�t�+��t� m�>��M��}6ƺZ�J���kcK^?l�#FzQ���rkɐ�G�1�=2���Vd��P�r�{�1d�u�j�gmh��_R��޺ӜƝ�R+��`��8]1�*��P���"��梲 �h4sp
f�dq�xY"�@��< �pț��O���+}��VJ� 8�W�4���";}:���F����u3�,fI����W�dH����_��$�c�.K��ŠA�	��%�A6Tp0���)70�w��!�4eӰWxz����Y���k�Ύ!Ih�+O����rcc�Z��'���f�u?F��N��E٪��4f�<�ba�����4�J�]l���m��j�@�},*+��!�ifV�b���<�k�v��WKY:.(�CY�R��:V�%��{�:���*���mzg� �����-�3|�����l)�j���4Mp]j%��-�_{��-�ً��B��~���<V��Z~��CI�>��=��k�!w�itoo�&�M�J��
J����sPݵ��K KA��*9R6͐�µ�1���p0<��B�na�=_���]�:ܐ%�7�4U��������2���e�T��m"r}�^�Ue���"	3�S�<��N|�����v7�&�ۙg.�yL;���Q��kD%���ه��P�9�%�ERIFF��y:���������r�$а�Qi��1ܷ�ۧ���]n����o��F�ٹ��P����MW*�E�A����4
��,�uS^�����:���L�q�,�.8���0<���l��"�ԛX������{��
ڢlҒ�.E�8 ��*����Xr���-��3��ڪ.�	��YV}*�Y�Y���4�}K���"3�+��-��)]Tw6�I?�(2;�;IX�������O�bW$��u�v��6|ʔ��dNW�Bokm[V��x&aߡ0��)U�
G�A/�q>k��b�.*���p���>@�͐r%��/�|G����vBZ^�^�V��
����W4�t�쏮�{�_��g�#^\�U.��X�r���n�%((��V�������s��w��I���U����c9Yb�%�D���S��!ϒU��D��ɠ���4@�fU�xw �KI U���N��'�%D6M,��X���|�� �9��.��A^��=5b	�� ��k��;r�l,���~g,ap�/5���&`fV�Q���[66Jv��"��\_P�P
�	mu���k�����g}�V6���&u@�k� ��{�Z���)�������4I�I��0m�'L��-<&��͈�9Vu���意y���uZC{:qW+8�2mywz��W��#�ѐ2��0���ky�TQw=�<鍱(Da�"(OM�P�[:4�t��Y>3��Vy�	��@X����)�V���ٙ=j���w��ȡѯ+q��z��$B#�dXα-[# ��G�~�H�)��~�7\�$� �o��[D����h{b;tW"��6I^g� -_&% S/�[:���B�zFO�� �MhXӤ��@[���S��&��#�]��FY�a����F�9��a�τ��g��+���
�-���p�/Sz��H��9 /k���6Z�񅘮��9t�'�+�%�M	�1ރ����X|�B��8���a6�b����c����Ѷ��SD�Dp��|�F�	����_�u���d���6B1�4-�\�Ѳ=�@�d��[�eXމ��	�	v]`��`cfژGo���y{̘���1!!��~t%��M۴�۲����bA��rۼ��;�wz�e���h�mLJg!�Ֆ\�����*oS������V�D	�;�h:��I{�(��=)�~kf�4	�R�3�	_w�A5^�* f+���Wb��8�ͤR��������u`�T�Lȴ	� ��S9*09{����_����o8HFW΂��N�}g��s9[z҆F!��G���k=ާ��9��AO�S�3ձ���Pc�TԫD䢰1�t�_+6o��
gY�:�%�lP۞?���d��(�amF%�"4�pH�w�*{@L�H`�ǯ�bT�-�(�w�ɮT��$��c:����t��Y���f��`�0���1��<j���7�a۲15���4�\��E�e�g�;1�߀S_�s|?�W����()��A�t����H��ww�����u/$P��������BӴ��v���WE�`Q^SOt��u�G���.�f��F`	��w�K" 3���ܥš���n�Q-)K�cވR��9�KѦen�ԙ��/��=� �0�XZǥ����&"�'Gh����D2EM *{�#�|��6�tdo��E�i��!���zIbk����'y"w�o�'��*��1Vퟃ���O�	������zз��;���ןSR��n�
�W�/$�C`�BP�qn��w���<(�S�%�=�����+��!��)@Գ�?:C�c���~<��]80��Ye`c2T�$7ކ��p��[��f�k�s��k��y:�!��>x��IF�`(v�{Y��>/kuT��1,���J+� 0vK��tF�C�b�&,�N9�0-ip���IP��e�?}dvAcN�yd�A_X���}E��V��	�d�����5�3�������
]������V)�[������C���!2���c�(S����/Ġ{M����8�:����$Z�p�w��GK6/-�J<H�km��-�z|&8����L_d^�ڰ�w��z/eT��O���2C4Geo_D7P�{N��Lc��u�T���%����