��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��?�I�J��zd8�l��%�;Z�	[��O��W �]��rd��k���S3.e:�R^u���.YY
�V�)`����j>t��{Ϣ�Q�߆S��i3��*}�fT��}�)��5y�G�L,Gf��;������X���v� Յ�M�#�KZF��P ��
	j��eJg �.!��ۿ�3�y�z,� �p�G��J	��Njڪ��I���CLm�G(�\)}^kx�#}��O�!�1b����a�ӟ��C�$�⋏Y[RR�=i�Y=�|����sD����*M7��A���$���>*���
���,[yq�������w��z5�+�6e�o���$I�'!ĸ� �f��N����@o����P�H @:�����\�]a����,e#�L{!�e^	QgP��M�#��T9Zi���FV�/k��7��#���.�υ�eM�+I���]21't�ɷ+����ù��gI�9�����.��I�����B��H"�&�G��>���((�{3s_�����z�NO��ʏ����z���4)	qCh�`��M^ ������,·^ɅJ2U$o�
��&�E
j�n�o���5�	�uF���;�Y~Z-�k��0\}��4�NpmR�������?�4�~����Ib�/��q�I�e(-���W[�`-������Zq�g��gO����\O�?�G<��I���;	�����/�,(�=�����/n��p��ÓS5H�3uL[���A��Q�3�$G�Lk�Jf��*�>��3?�J8{�3}��5`2���(��?*�����n�XIE���y��iq�G�^�U��v�ȥ)E\�ұ<J�6�:�[Y�ĳ\f�\�j���D�MS��C���	�������Ǵ��>a^>��Cx��q6&�RH4P2q7
EsD5��d����L��<«����x+���%�G<S��r�T��>�Z(�	棐D�'!��e�%jf��W����X��u������H �����FR%@w�#��MK���ü�n�R���E�a�bA��y�&`�ٻ���?^�N���ռM������|,�����13B�:�����%-c�b�ԫ̦L���ė[h0�x*��ҏ���U���2M�1]2�����%ro�B��<H���{�Je�������'2_q�I�@-�?��Έa����r��]��ΨW�����Y�e*a�φ�u���8S��>�:Sy�?���u�m�M���G���_�s���Ƃ��VgWNQ�U�C�p0Oy��l 4�,��	���u����{s�{z	��y<o�叇�ź��+�ܚ@�g7$�.ȻF�&��~MOE�.�GＹ��qW�͊�VN��9*4����82���OLD�z�'�"9������DyWH���v��V9�\<Cѳ+�,���R{�EZG�0]��#)\I��L�x�ݻ�*�����Z���I��~�z!<Tg��5dn�ʫт�ZO�Ubmp��o&�!�
l�Q9��@H{A*;	^��r\�H�-+W��&�4C�]�y3��P��>�y�����R���T�Y��L���?��6��:�b�h]���]N�{*<�~���DM"$T��l�>�FzRT#I�}x$'`w�mK������Z	*�,���9���QU|}��<�3rD��}b1�;�:u���J��@�=��%�58���I�:�d����ʏ0���E3�XDE�J*MY�[s;�׎��5���&W7�9���I�2?1�=N�t\�Ry�����*�ZIK�1���(��0�$]�9��C�5ȓX���w�?R�<����&��,I��jױS����!�����^f_���+�T@��<ٽ�W��Ѷ���w�O2H�z!
����:�#�"aH[__O��D
5��I�N��Q���v��,{=-�!HE�r/��6~�-���B��l��D�Y1
8�j5���)�C3̀�%9c�V������Weղו:M, ����>��hC���i�S`�{%�������L����ab��x%>��Ў���t�<�1C�T�:s����8�܀^���ۓ�1 ���už�N�yƍ}�'��7�)��_� �~	�>l�!�m �]Wp��O1�R�|"�u��#�#?�.�3��au��"f�+ Ҟ�����|��(�+A�����s�T��z�՝k5G1�����\�8��#o�ά�<g+#��\����4�����1}�xk���e�akσ��XI<ee��k���<���x������ߚ;9s ��!�v$����<��Iל1�&X:���":܆{-K�z��mg�dGG�1�B���խ�Ќ���N}um&uU��i�<.bd�!���7�Cbb��.1S��{����}���8*�$k�ZJ,N.���4%u��_�o��o3E�<���c���
��PJW^?��y��\S"�	�o��8]X��s��H֧G�����YhB] �i`��6���M�reD�wNýJąym��w0��9���B(�2u��k�d�,�RK�����H5Q0�s�Q"e<�0W�t���$A뒭]�û�)ޞE��"'1���]��P��o�\����|�|
��Pw��"���u��������mI��WZd�V��> c7QZ����e�����S���7���0<&寤�c�x/�=�gf�v��W���En77����Ev�hm``�u$�Y��I��QQ�[M��E�,�t���Y�"1�hgՑ-i��y�i]*�8��g��`6z�L+�SrW�T؈\V�ՏlT�
���j:u���!d=��',�Oj���ПG>k�����s#X�n*�5����0B �7=f��˫.zm�p+]Tvm+,T�<��w	
�b������#V\�yK
��j|R8����@V`����(h�s~��Y�͵I`v����1���+�ƕ�(��oe�����#8.��c�nF��+^���D,���o,����gA �a��g�J>M/�ڇ��Q����e,���2&�X�J�#������y�������)jH�d)f�$�r�E���"Ks���|
#�ճ��5Ж_h�0���e��*����z�����й&����2� �Z��2wX�`0]*�ǚ�L�j9�4+��j��_�BD�>�M�,��O���ׇ��xM0j��M�H?@�����靨�������ߛ��
��K���$M�xػ��_�*��lat]y?�G�
����en�D :et�<��P�^�'14�X��xi��I\�-������7��sz�2����ĝ.��V'����]*��l��[��~ ���?d�L�M��#̢ʑ*��.o&�Sl�iT��8Ow�@K9��-#�r��g�u��Y���m׼�]=&R�qZKΞK��r��:2�,z}v��S�g�׵�VJD�H�ׅ�\E2��dpJ-fUe��?G�Jު�u�l�+GZ��<ϫ'gvK.4^w�
9�~���3\ [
t��0RM �I��.
+L iȕ�RN�OE�}Ρ�`�5?4�S��aG�,@:��jCD���QW���5}@��C������?��BN*��3�r)Y;��Z^+��?�����u"��!��q���5� �Q�襴'���f���D�7���⧱����������W@��#��١[����Qm�us�{��X+p$��S��樨J{	]4�'��`�i���t��< ����-ngI��nm�@�'lT�hEm��/�ߴ�.�qs�X�q�mh�;�6���Sl�- �J�����R�~��¡�u�ڼ�F~����/8�h�Y�5Ga9��#��[����_}�X�NB�>��lk�@�A��$Z���~�x}���5[��$��6c�-D�L��c���VF!�l�}aS~1�]G�� �ޜ���&�U(Ϧӡ��_<?��ဏ�[�_��CĹ
��@r�h%�ʸ�(��}�ba\��*��9�c��~������&�V,ZDW��,#�!XP&y��Y׮�Ҏ����C9p���5�9n�v��2��� ! �D��X\���4���׃0# QЍ/���-��-l��DXl��U�`|��G����b)Z�χv���hĉ���i�h�3%�ɝ�����=�F��J V�<��lPj�k_�sE�HW�V�|���L�Q�d&�ꡲ�58�Q�w[��lz�>Ľ&��TPJ��*hr0t5q �+�Y*�ӻI���4�ܸ(j0Ǹ���n�'��������<�� �?�1@_�ß��5�~jC�YrX+��-^٥�FLX�sq�g��I���iF�? ��c��I}��Ω"*`>y���R:d����4�#��P	��z��69y���s�V �0A�Y&�§���E8��Cl(YQ��B3B&����cÂ^*~�D�Dvj�]��������X�]|�v�ڰ5�4,�+Ɲc�c����2L1�;!�:[�=�_�Z�S�3O�俐FVs�Bd�V��O���L����@�0:�(�k��+�܁z�T��MM����K�CP�sE����A����4���L�N���}+�bɅ��A�l &]��(����Y�̙�u���#�kQ�wGT3o�=�L��D��x����3�ly�̌� �Eƪ��&�^z�������,�'�Db�tro���[s� Fz3��u��%m�Қ���jb6�.�@Y
�	�h����.Gc�x7�I�J(�2�0�1��@�G!Gu��tV�����so��Kx�-j��p��Hs�p��n��� ���X�g\iDّ�yr��Qv�}iIWZ�	;���2�@lIʪ��Uﭲ� U�[���6�[�1R�e��/���]:���^�����>v7�DB�I��7�I5W�;�e�{�i�x{��E��ϊ���$3�:��wd]������6%4�nXYB������r-��pm�C%����K��6rɩu�����Wu�Z�:i	.�ܺƻL���B��Pԙ��n����.)F��:r�m��鸛�Ƣ���5�{h��t��]������~+��R~���	@P�`�dL�O^�G�!�/^���Vg���	Z������㞮>gYİ�I�<���]�
�1)�(G�e��ky9�j^�
�N%����2�mz�S�;�d�3�n~��M�B�׶�Ҋ���t�l6O`wy�[���"�j�`�Df~9�6M�?�$��%l����n˅�:�V�ZQ�6U=�4�&�J�e��}D�e��"�(����<m��snߵ�_�v���A��0̌��ʯ��x��_$dDqnW~�|$sf�X]���Y�����5"��pCI���(�������a�:�Μ
#�"j�2g'L
�d0�j�=���V��N	��lQʩ��^=��p�*а �//79��l�ۇ:q�N�x�E}�F~�2H�QB�&(vc��قCJ�S�!����vL�0��	
�x��L1S)7;"��o6?g��sr�&�]?����2�7J׿&�-�&��L��Z��S�<�9�A��=�3�R�F�IV�>ԦUyx�$��f�R7�T�3֯x���Ϯ_��.�`鵩�O���@��d 컣uD��	����v��
�ZC9�I{�kG0�o{�7O�?#�9*���%�I��4e�����\�hp�w�\7�
%�E�ʋ�r�����Qf#.\���t��(t�z4eu�4����mω4L�P�Dr�"�Y�u�#G�(]�<�-��"�A�&9�1R��L�q3��Yl-��ښ:3^Z��H�3��vrY�4�Ʊ�c��',����B�G�O5�v�;���Į�b��>cӴu_@wm��{igN�ux���p����gsi����?	�i\�zX
0t�%Pэ"MH�jwX&)+����\+�������� �d���_��^�I�ͫ��xN=�(����� ��(�g�6�xm�ָ��՜k�k騲=��x��+f*�.x�W����=�8��KU� ��@���t_��K��9�k�N�X��sI�d����)r���$�'XX�Q�7'����͠�L�c�;[Bc�]g@CQ���bS�B�p���)+G�������7!�8x`bb����r���>2g̣���mt>���`�[���1���&V�C��/@�w~���c��	71�n��އ0kt�$�,|��;�_�#�	t�JqwlCIu��)zoކ?b�~���v ���U��A��)*��2a�EPf0FPf+w:��TDE���M��y\��ԛ'����9ۡ��>���y�J�@���}r�R���Sv�U(5�68��K�����*�������K��d����9�N�
C�a����_}<�����i>ms����\��є�ko�+�g�޲�hñzml6:t~C��������!q�xPx �Alg3<`���W���❽���t�qo��	H}����x<:5="��Q�����x��^���>Ϡkѧ|b71�y����t�Z��=2s��Nf��˰�4d���{��Rl�w\���`��-و��8�]-�p�8Xw�X� "���" �a�ל�F���ד�����㫞��N��R�T�D��q�4��)��!���,�x�s}w�
�$�G29����k�������I���5�(?Kv�'"M� h�-@��z�[���X*(w�R��RB�Em0׻�V�*���M���ۀ|N]���n �f�Bk�+u�[��\�z�ֲVT8v��v�m8\��8 B��>(:�z�-+Q��S�-�).���@��GA��"�.�G6ըմv{6�����7���JxC��ܣ��D�FW�������a��a�?u�&�O�W#B���[����x�+rP:�	y�v���=�݉�\�����K��X0r^����B^s��ur)�;%���s�ð�٫ ��r|x2�������\�Ʌ��7%�Y$����h�'��󞦭�a���r�铜k�o���X��Pe�L]�ф��w��}��w��X�Y��[Av ��y�*G��uwRQ'g0V�7�J�`��6 ��KҌeQo��I,'Cm��6k3��J�چ}�v���u�D� #��*�Lg��e�Gl[��X�u	�O+�����B������h��f��=GH΂��^�v�P��dmB�Ɗ;�L`�X˝�g�#L�,���/v�.G����=0��	ΛG�5�=iG��<2��\�{1V��/��E�-F�M��^���5u\*&1�	.\?-r�Q� �Qz�+F�Ju%+�@��~� ��l�f���J�{SkC�;rhQ�k�7ߺ�M?��M�-^ߨ�b�5W��Ү'���vh���*N�b?w�UH��7"�V��
�q'��|�lO�2r���>����H��i����<v)���}��ɻ�����U8%�	���<q'�*������-�MD��M�k��#����z���Y�����$I�����ɒw8Ƥ�M��t���Z���Ї��F��P���r�#�ً�IJ�\
�)�z�g)9����fg[H���;th��}9��Fߴ㲬�D����s#�m������m;��CI��|�x�pR}��#E��ZI)��q�}9�6�z�i�Ӯt���λiX�զ7.t�4�c�諛����7�:F7
Jw��)��]e@��j��,���=iS]�JV5�P��x����"4��
��꠾¡����� y�y >Ex�~�{Hr��̩��$��A)�Su��a�8�<w&y��;w�֠�����',ZQG�t���T�:�(R#� �
���nkz=����MmfV�ʭ��_F�T��ٲ����_�~���C��."��g��D��ss���7��=*l��q�D��'s`gF?j��Ŝ�Yv�0F��@q>��/������]�GdέyX��)k�L��װ"���V��g� ��q���5y�g�,��f7��e����;b5���q0���:Jp-���6����ťO�uOhT r
������d|5��ז}�������{�D���1Hլ�& �5a�9�l�-� x���Z��4w��_�5;�#�,Cz���G�W�[y-ޞ�+�L��n)kOS}g�qw���h×E�)�?f{���Sb�J4�yk[Уq�F���7D{ �����̑�SYa�:�D�R:��}�F̣w�+i��,#�Cntk����d�Cץ�jYd2�!���j;���j�?dw�����%���7��i��%Q���u��NY�;G�Z�8��f�eG4���B�	<E7ҋ�-ϟ��κ;s&���#}V1B����ن�`��;Z�%�c?+;v�V!=*!Ua-�=l����;;Ee����wa��Ś�¡6� �7��[\�l��E�5Vg:*��9��n��.k��Ղ�1ohBmx�j��E�XZm���KU �K[�:rjH5!���`���0����	�s�\�Y�c-��,k�?�L�V�3��A�iO��2��%�bz��sR�%�;�
��IOWI��i�~�!-g�����4b�ǿIW0'24���D�|����K
����Cw�4aԜ"�OV�fY��OJ����/Na��2ʰ-/�d�j%��n��f�lr8�����ytF�����ɏ[�E��� 	g�lm.*;�Q%�P��Jڑ��ˠ�ˬ�"�B�X�T2h���04	�B$CG��a7�o�}0��������P�}HE�J�m�$<��7  X<(�ێn���qu��l}��ȟF)����/uwe
\�W:38���n� �X褺�tĻ�9%���$0X���`#Aqnmx|����=^�<���|�M}�j�!8�~��\3�V��a��,�K+�ϵ��zIL�7w�{|���ݶv�����.���}���@}'��N�V���i�/�9���'��X9J���J�Ǯ�)��^���7�Դb�)��Vs�i�e�<�?)�)y�f��������q�t@*mTy��9腛���ў�]�����K��Z��J:�G)#�E��4/�+� ����a����5ʮ=	���e��80�6�^�r��d��q���o]w��cM�έ��3'J�T�V�t�[�~ ��gb��'RB�~V_���^��T�d6I��������YI�v!:��J>�2�k΃�uB�*��Iy/-M�+�9�S=S�����X�96z�J�V��S5^�k�b���|oJ����tHP�P�b
A��QL�����y�I,0��d�i0mn��.�	����c u���:�<\3n���x}PVB�zF�hU4-:�@�`X�B�z���B��M^��u��n���=h&�v�y7#��u�E�⶟OWxD���(��9xv�k����,T��w�P���0�2E�9��W��a!�?��
�'�Tj}�+���ŝ3"��B�F�_�Cksɗ16d�^��A��ۡ��{��r�����wj�1r�u�Ĵ[�F��b�gu��}�i�X��Sԉq�t�qbi$��J�������΋in���a�߆1�c�����0�A�U�$^�,b3��AU/��G�`)���O7���V�=�ϸ��ߴ����;T���$;.�-�r������fm���Ƶd{q�pԕpH3���/��i%#��E�8RԼ���tK �5K���������\�����%�m��!X��L��\V�}��d=�K�����Ӈf�_�=�V��C/��(j��J�P5ƸqR�W7�"Ua��.�o�ZܽH��'j����djNWVI�V�:�{Bc �H@�i��kl%*��#��ם"���G��d�ξ�m�G>�)ɕ�d�Z�XǑ�4��A�3�`����kO�F�x�)b��Fq#y�sF��*��s�G�BfZrw�~�z(��ھq���D�z�����mJ��V��ʍ�ڭUĳ�t��hֵ�*�;�&��QU��c ��g�(�#�6�s0H)g���{xm��o�q�G����AJ/�gӅ6�&jl����]@���I|>�,�{~>:k����x�~�Ȩ�3�V����Rw���y�#fP�ǥJ����-O+�,'��FmH��D������Z����&P��
G�. @�ej�\����j��ANɺ�KCd/4L~��N�@�h��B�N�%�_-r��ϝ���B�x�hP�E�b��:�

��t��gem�h�� !�g��*&Ms���	���m�8cH��.���Ly��FL�,-S������ 0[M���[�!�1��tP����)�uMuKwnBl��'{d�-`����eΞ���ǜ�-�����)�VD�������' �92!WT�
n{t������D��Ec	t���������1����קkNB�j!J6���������C8����C)����K�p�B�ic�U"-|�`����舮 k�.$Zpg��M�a���a��Y��+B�2< �r�����~_"
[���H���׬:�Aǥ�ry�M)�Lm����N��2w�((�4I�I�3���4�t�Rڧ�I{�,�$y�l�
Ny/����q�]^�
B�98��+1���;d&<L��� ��*��?A���(���{��%[Ä�CI֟��d(�c{���8����i�����.R��n���9���
@ ������߱����u<Ĉ���S���FWp�ׯ�:/b~O~&���U$>-\�6FV����	T���[�[��\�K��G6`��mYοڀu-E;N�F�eWD�hׁi�'�h�T���F'D�^�o�C-��Lv���%jԧ�/�Ja�"�~ǡ�O�H������z��bd{'*�H�%\c��9(��J6�����	�O��Z��e3�Z���ز������AӔY�cN�3���ƷH=J�)�}G�~"])�a�oJTn��8�*(q�ѵ�5�����X�b#�����G�s΄$�`�N���P�x�^���sQ��!�����}n�=���@��W���q��o�����V�۬���}̩g�T�i�ζ�����9|N�}�|��--�����\��m����p��*��W?g��W����R�j1/��|:3��-G�5�@�9{�0�ӬPf�����^0T��T���N����ӟ9���*���} dV��QZ�2<�wj{` � �P2��S��&�����&F|<я�Ȓ�g��i�*-P����s�����9����Jg8t.��l���4�����^�O�� �Mv�}�)ȼ{`h癙��(�j�p(�mڨgc.���!Q|�q����3��!����˧����a9wV�?^⳯ڝ:�EA���w����M�"I�І��|5�̔0%���D�s�-x��'���˲xB剷��}�����$?7{���c��F�)��꩏���F+�_�Ɛ�k�W�Q��־:gW�.|�@g�en7?o8rH͂Osd1�|����2��S4d[k�Vl��ţ�Hi�6(���å T&��vԽ���f��
����1��r+����=�c��N��p���WR��汾���v�S��ldJ�4��z�}��K-�i)լj����-3�q�v� ��]��3�a�߾�C���{U~���3Z�-4q6�ŞN����+����fV��Dx*�['�;'֋�&�ױ�*�Şs�x�@���<㶚_�4�a������eP)�1�t������	����?�%Ab�&�=S:�MJ�6b]u@QyqU��e?z�$����<R���,�<e�����2�r񁳵�.ގv
r�~
w�Qը��F|
�[�Z���?��_%�\y" �����ϳ��E�q������;���|gh'�>�����mS���ߘ}rkMT�Wz��h��۠
����L���[�?S���咮W��(t�p��=v��j���2�RG.�,�+���J�T?��M�����r�ڧc��'�b �s����{C|�҅!Y6���R�|�#�D;���ۺ4�������<�����cJ�� Ƥ�uE�?�C5=���Kq*K��K:'�	N�^��>�P���^���}�����`	Nj�5�1��-�h�&���'
lM+�I2y�z��ѱ��r���5��x_#=u�|���("��1p��
��(�|]D��FO�=r�_�!* �"����]r� �i�>�P��S_-"������O�Z�xr�ݺWiW�q`��q���@��:W'�l�f¬�5� zЗY�O'�#���D�	��)���Jk����.��\	䫗u�3盿|�|L�m��L��O����HCl%�2r��'��Й_�|`6�� ��#���||I�Xը>�k�{�2}�0����e��+�")Q�tơw���q(n\eD1E;�E���D���v�;+�)�񟋔���+:d|]J@�.���~�xE���̠e{#���/�ag�ѧ�뒬��/]\������T��n�5 `[�	ף�N4�3�k�%U�^����7���j$�J�+��W��������5���9|�;�q�8�9�%q&�������m���꺤�k���L�`�JRQo"P��S&��{���Y��������b�H���S����R��| =P�_���eE�Ӑ'.@���6�+�nf��:�4��N���}���s���.K�������GR�=�P|�^���@�S�����q_H�1f!5��T�Z�Rj���l�%���B�5��s��,�V_	T���h8��%!=:��#��@SO��&��BVCud����������VpH�k���ׅ���c8jZ�W��ݢB��%�/|��C
��,9gI�7t�#�_�� yl��U��n�OY���aعl.�Ŝ�m^N	a�Tp]�N���>*�����V6�XLIp�&E���+I"b��g.YʦI1jW�H�� �Q�%9Ɵi�ؒo/�i���P�*�h>7�R3ޡ`�+��������=E���)�ΗB�A\jm�Ѧ��'G������^?�ōf͜,
�E�j]��̝`�~+�����}�y�G�G�!?>��i��5�b��. ⍛��/�@A���@�Z�d�_�U#���4�DX���l���`5kvw����L�D8��pF�<L�h_���D*�9TcaK2
P�_�V�5����_n�_U�r�Z:>�dW5n鋣�{
W�ۅ��B�Z�D�Fu�+ȿ�Ù���4cB�έ���p�K����� 	P+Q��V���~��*�.Y���1@�@��(�;q�t�\�Vå�͚��3���ѻ�Ȼg�3{�}(':��bӀ�b��m����hsbR�H��g�Z�S���m�d������!�y*S�<��9�}=���t��R0+5�X)gQ�+B�j�6uOq�{$�^��қ��"�Jb��QV�4�jȦ<���-߄'�z�%�[�"�G��G"����@Ez0n�^/���қ�m�,�0]�G[
IBa�I=WY}.$-�]+��/��,�QRm�:��I�&��݉�m�*F���<�VHHv�*;������@/ b��^���^�6����ݡA\�ChWP��XNcWړ)�Uĺy��@�_}�M��]c��))bh#���B�ιЃ��XLsB��)�A:����nv? ЋX�GE�Τy�|������1� uBu�a�:-��X���^/����tW�f��\qyH� 	����+ �Gn�]ݬI�ss]K�����a�G1�"�X	r	��c�Y�.�ŝ�U(�Ͽ}���Ç2�t7��j[u#=�7̫U����'�������9�h�G!�@�N*��B�ш��jƲ��;<e�mF7��<�J�X�jmp
6��e8������q>-4��H�1Z��t>��}$�������PIs�c��j��p�M��ތ��֘w��֥����r*���e-qeƭ�b�7=Z� ��&���$�2�+#*]
[�Fǯ-�~��K�0��f�� �3=z~��褿��66����=e.$�PԆIa\
(�7�ϟ�^tv)^Y,CJ$�ܘXP`S!U	���A&$Nv	.*W�P���7ގ��ǈv��:0U����ުK<�_ա�� #-�����vI�����Ն�8�����$OB��#R[����vB,��������I|w�~�Sze�%:�������k��s�(}	�X�G���t�WG��������D���-D6t.x�ܗI^h�Va���b"z� ��r�2��H�R���B���1��凜�\�1�b�N��v�w@�Yd<Su�EA��<w[�]�uyo�f���b�;�Qb4I']����-�=��>2��\���ׄ�;�#p��T`����a�h�By��.u���2p�;#L���z[d6��1�����!��}(7 �k� Utʲ�W(�Ā�Ѯ8�����g�B��0v�B}0�AS�c8����$����\��RK<�=/r,
̀�U�L�A,�9*��'j�SǍ���	m��y�����\ڈ���n��| ���0Kvr|���Kf�Vʛ������G��W���M�L����hI�T�bFظǭ)X���d>�%�<և����it_�ӻHE�[Y����s�H��Iٕ%���`1��:��U���0���K����`l�v�\��b%��d��&����`�é�Ͷ���1G�r�7ޜ6���/��Y�4�u"��H�5�_���o>�~���6sP�Ƶ�
�,�ݥ����c�y��b�0����"E���(A_�=5"M�D,�_�̖M��{R��� NՂ_���->Q�F���ޫ&(��;'�����x��|Ĝj��H�� ��E�T�J�y��H�Z�8(ۛ ��j���M�`���{�e`NS���=���֫�g4��];����3���%��hn�iBْ�q?����2v���H��o<�k�6�26���uD�Ջ��G�&���ک��1
m�kS,�~#��������.�͙�x�*�����t�+�̟3H��[HYj�yҘ�:U����R;�M]#	ㆊ�$���Q���6�Иx�b������8#���>ݜv*�P)\B�XuSFd�bny�S���Ǥ�oǙڪ�zߗʚM8�ڤ�6�`jm�!�)�x1\C�ꠄ!�_�[�n#������]	�F ������H=�F$��d�(x�i=��7�
.=y�PN��,0}����3�VK
�\U�$������V|�π��0�p���ϐ�0���0�K5����:��rP��Ze�Z���e��;"vK-�-' �I�[��Z�W�L��7=]�BR�x��Ϲ�M�|��G�
��l�K��C�F	��5�b$U�,��pc>>Į�CZ�;x���jt�HI�dǬwok@���Z�����o�<I�M��a�v�d��o�N��<�Dwof�|�� '�;��^9�-ڀc4u�P�TV�2� {��0���W�� �3�"�j�U�i�V���7�7$�g���cx+k��?�k��G�t��!Ta��p�{dY5cQp}��Qd��hȓЋ�XK%]�ID�W�DA�t&l�	Qw��P��ڶ9����R%E�ß����;7�.2K~���z�������"��L������=�u�A8.bD�?���3[7;��Ϣ��V����ӏ x��=����S�ܷx�;�YGF׏�^��-ރSÉx�lZ��!����r��ri���[r�((<~l �;.�r{>t�7,ư��&g�I.�h�/4盼�28tWς^m@3���dyS���ǿd��eT����H�+���B"��0k��.{d�V���.Kʜ��=�9�.�m��A~�<〆j"b��;b�R��>陴����ܳ×���1ʘ��@^]��aYW��&�z5Y��_s��&C�#�>J�	�m��4�1��<�3B�
��ᨒ�Z'̲^�xY�]#�x�2�	�3h�]���[ľ�8�:��m A�D`@c���¾/�5cL#^�x�<B�D�p�z4�8��_�]y�}(�]���ƒ`��s��������(),�)"��h��1`:�7�͏��Ow���('KcS]�{���R�����$��-!����	���� �DW����� ��2�=�H�F`U"z�㺩�)�Q�\�VD��0�`�e�-Pc����/ˤY9���)��h��m�l4�b^����y��1F�i;:7G��[�������l�`|�D4�[�e���er��y¿��sH�XJ�'�t��S� ���Ο��a{��|�yF�<^�u�ӢL�X+D��x�>��4m�U�B�L��Y�ȕ��y��.���g�>��!&*�V�)!e������'�����~��}�4�
1�vk��R,���'�O^߉��NT��_��{�ižИ��xXq�=���O��*. �~�#��;
>����X� @��W8��K��H�G�L6i�?�J<D����`]�k
��d��_Gr�7cZ�����3h���C�}��J�.�����m��<�9{bn�H��.8:��h�=���?�s�Cc�v�/����XEa�؋�w��I�\��i.O'I�ƨ�C�A�^O.�-؇�mֶ��	�F�����1ǿ�]M1��u*�2��KD��U&���P %F#~�]�X�l��O�7AD��GnP��'G6`fg�#7��M��>u���<�
�}�*v+�TGg\Úb&��g��>'p�����>�p�jn�K��r�X3�қ�J���B)�]�Crsp��ƣ�� u������n��S��.j��Ռ��1��ؔ��nǙs�[���~��F����&w.��V���W��Z�n�]�i1�?�V�E�3D��&,��tb�m�Hx G/��A��5p<O�t��3�í���ZT�6c��w���s������8�	��<����o�/l4��!: �@��%�j0 �ObS���αA�w.(׹���v��wS�z��Q����r$#����_�.s��PQPDh�!B�x�(�<N���p/�j��B����d���l�Y�T
������Q6���oz�A���)������k,2B�)��Ǡy���w������;�,��]�\�z�i�U�����/��E�8��7��4�}�C{�et��$kq$0��MG�nm����Xd��	\BX��>|�(� �*�b�������Q����E�
r�D�����R�wZ���֎H�e����b�I�����cj���:��Mq�N����~�-Aw�`�e!6�C�3��L�}e	��2c�!����}ϯku1�rS&y��B拎�6��j|c�8ӫ��m�<M0��q@�MEq�KL{��&�=z�nұw`�JB�^� ��義���f�*G'�� &��?HĎ�#�u���P���5��G����P�9l�S=��#&*�%���B�*N	�2l�x���-����f`H��'����w�Sf�J	7�7*�YG�17 ڟ������Q����m��t��lmn���J5�h������yօ$�<S3�n�.t=D��Ų���g��Y��D�lʹ�[8}�C�$~���]r΀	�-`�O�S�-;��J*�H����A����v�㰼T,�
��DS&�0�`�'����*���UV��Ȱ3-�'�L0֬ �(0$��-��8��JP�$w���d�7zer���P^����C{���7��\i]1��Ê�8Pu:.e0�aN60�ȴN���t�� �&��j�o�-H��� a�S��A4$�@-i�h^�����z~5=��Б�w��rS�V [N`��=�q���\�d	� B1��m���}�h�G%%Ok5�*x[f{>clBюz�����x� �0��W1{6�J���bȀ��'���)O��{���+�9v"��*��*�sa��<��������j����,�DC�� _裂g��C�'��3 �������o��?�t_���7I�nk,���8��V�	�˼>A7{z�!��M��W�s�"'��Ȳ�}�;����z% _�>e�|��q����C]�6�R�*k�x/��������싚'rѧ�-@�y|%���1�#�y����P'mA�W�R&+��Gk0&9$n�G�J?Ԗ@�%�ų��Z��r��E�T<$5��dQ�8p�>�	y�ź�o��m4����9h�	��k�^�蓂����+G�=bܫ�f'���(��g������g���Z�����]��Y�+���E�^%�^Dz��B҃������ǽ;(��A;Dw��;� $�F�eR+�9]�:Ht
�vZJ�6
p]#�Ľ����ҟT�^�Ey���2�0�׼	+�T�`��]eq������Vv^$�v�OI{���P�x�	�
�4�	�񭽽��З�,�Jʟ�#�Շ�#V��`�a��i�U��^3f�;��}��ƧV�u����+A���!����e�t�Α�Y�p��3�� B;&p,�`�j�C��Z�X0T̟J��2��Cȁ
�^�g,.p�Kf���g�_/�[Co47#C��sX �@�7����Z���blj��ӵ�;1�� Xڕa
��gt��P�<q��x?�_��q+�:�t�?�#��1�S*�9��k��rJ?;W�&�W	���y0I���ڶ��ؒ1	J��.昱җRŜçK��XT�)��(��������<q��~�p$ۆ^�F��&�z
eb	�[��u$`�6������l��o����	�����N�`��;��G�yWp���5&Ɂq� nc�9����Hf�d�S����x�$i��Uc���r��Yw���h���9��?I+�i���ii�go{K|	ó�-�6e��X�7�Z�A�G��4l�dʰ6,��Z�c�V!�ŏ��z2�9�[QdM����(+�{<z3#����AR=���A����MQV�/+H��HX�Kr�	՛��a�@��D�H.�ֆ�fv,4ַ^@=�I��S�"�/|��7�$Ҙ��$$�@������S`���5΀1�S���B�>"���h��}�J�M�y-���w-JuU-��}������|���d�D�F�K��d�=v��3���8���L�dƞl���CԔ	���1���*�w��$p	�)� }�� ĻU�t��e�<�^,���Kx���5����zw��_ ��R�����n�!?m��7��t3�l��tEWt FՍ)����@Y{%D��=)��1L�>3]�z�� ��� w��p ȿ��ǡ_$_��\~����e���o9x��P;@����X)�����_ ��qh�`;(�Lڗ:l�����qJ����x�����*�D���eU�,[bw4�N��p�mߊ0�"{�E�>5V�!�&���	�, �v�#
��05�An��Vۖbl�2��~��dR����8�
4*o6׸���2�4r9���u>j��_�=	�v�{:���np��,��J
��E��-�:�Q�6�IshYJ��,@���j��f���������ă�Hq����X���E�STę]����`[��A��l���>��q�9�T���V�$���/�(�/D��P�tuC�w��a`�%k=	΁ks���_Q��o��4|3���,|�ӧZcя3��'��h" �H�D�@��s�[��=�zx�F��I�I~����鱡;�M5��2�-�Ώ� HZ���N�Q�;8|�����&L�k�gJ���)�k3j^H�Q�Kyh�C��G\n�G�V4�դï;f�`��o&=g�������~�Ѥ�έ��ӟ5�B�"���i�B���9ژ�Ä2�����s�u��v�+yܻP�lQ�(={M����o֮��^)�H��pG�ˢE�84�i)k����ҹ*7�ƍ�?ݬ8��7jV'ƽ��/5�F��n�ݐ�}��EW0�<�K3�R�{/�뜈�K2_��?���Z����	71dGç�Q�`�a<B󏺢�Zd�o$kQ\������Á� x��+�� �����QK��<.�A��%h���r^<��5wC4�C��*�aw�˚fb�ޫbg�r=���['�c�;�A��c��+�]�&�ñ;�d���-BD�<�8����?�B��Q2I{���rtq�8�I74����*��v��4f�J����+��,.�94
z8s���E��Ä���We�d ����'<6��<���!Ε�\����1f�F��f�\8�ePU� c�FG7�{����1�${L���:�!5�}�k���	5��20��[x� �^�6q4�L���$b�TQ���2ܖ�UI�ԟ�10���c��it��RP/��xo���h�Wl2_�*9�Z��)a�O��Y�1{'�y�k�?����<+�5>�׽�#��JgT"Λa��?��5%��P�
�T���R)�@y�Z㞞b�r��{D+��t��}	�Q��B���8KV�%�(Br�r�cY��&�s"�zD����`f6����dd	��?pO��9�q��q�W($N�$���ߍ�O�7�%FǤ�ig��
��^��S��C��qe��Q)���& 0N�s�Ć�9�Y�E��Sy��!��ڶ�>q'P�XQ��B2Z���e�O�z�5�̓I�����>��P����=ǹK� �k��-i�7��(D{b�)-O��O{�I�U����􇍡�@���\ώ ���E�P�怠D��z�h�vAD0b�I��xj�6�
l����p	��^:C����I,7��W�A�Q�`�pZv-x]C�����^� ��-��b��up����~Y��ѿ�K�+�Ό�0J��hO2�z�ڿQ�xrҞ[
�����C]�$G���m:V���ނ.e�f�~*������N>���8���Dw̔]Y��F�,@�.(,��!�M: gG�`sN��'�*�o$v��}s���[O�h��%L�3�db��T
�e�V�)����Y�fi�k��ZZn�+p+Y�,�n�1��<Po��"��u�ش�'�BA�4�F���w1�J� @�ޑM����"c�7�X{ ��[�a@~ �2�{��p����)ʆ�c�Ʀ���g��= '�])t���':)��/W�
'k��	��y^l0*��+M�&�����߂���"H��6��E4�W���X�>א�Σ����T�|%���B�<Ǯ��� $NEo�����ūf/޲�0(B��Xf�v��;��ɭ��|�@���Dd�n_;+�QJF����_�����P8�g��zl<(I�)Pd�l�I;eA"���9׹N��-�(����]Y2EN]� �ݳ������63�(ʡ x_)Cn
���S$ �� ��g�	�wG�pd��K�U����5����D:N���w{�ٷ�ڝA�	�/��-E�+�JYA�`���a:y-}5G�`���M���x*�A�2�k�����7b?�0��j��w�~iKA��EW附����	��iQ��@��/v������Q~���^��n_le�h�ݠΉ��HћF�h�iw[ݫTl:�A�eUNQ`ˈ��9�P�k�S-x��"m��Ԭ�Dق�j`�e&	�g�z�  nE1/_2�/K��X��#��<ǂf����I�5}M����ڏ�ڀK|�<�欗gю#ɺ�/��*"�w��N,�VF0�X�T�R�Q� Ԋ$%;�r�z��c�{M��D��[:s���%��tO{���(�@�Ћv+ؘw�~W�N�Yרe��<��=C;i6N�$9m.��kc��f�;�9���S�ɆN�o (D��eP'�y8�0�4*�#�?�[�"(��6�������ʊ��Pv��Ջտ��}�ȷJG>�F���3c�2����iዛ��Wx7�}����}��f�Q�<�kj�h8V����R�x/�������`ɉ����G9��E\,��A3�(�С�Z��!Oa�P�r�'O��N�!-��[�2!���O{>��K!&Z�j|�d���Mo�Ϡ��3o��H��j��~�TLn�{��l��F� 6-�d���~8~�|d�n��8[�����T������o���T�2��>:�m��A�6��?!!2�V��DW�5"2[n��bt�d}�Fp�B����:�F�G�:U
�1�uiξjs�8�12�?������h2x���W&aʥ�ը(�W���L�>{����X'=v�*��@:�R�u�<�#{���F~۾)m2c��u9x�Oe�Is(	Y�2(a_ML-�`@��@��&���G�!�k��<���^��nV�p���<dZ�����lW;#����3����?� �#�ȵdߧ���tҌ�S/&+9)�KeZ�j����0��+��KA�|��'�$ž�߷Z��LV�59>$x�T ��������o�x?0�_S~����SKsy�\_3b��0����p@Pc�+�g����}��������Ə�J�?9����'�r������˱���3� ��Z6{�����ܿ@�Bh���Su&�4�(�X)�2���ۙ_�Kqo���y
�O�	�q,c:Nܾu��n��I�~ᄎ�`����p�ī_�b��g��~�P.�`�D=!
��,�N?K4r�����#υ��ƕ]���Bp�)�˒�IŲ~�A^��'���2�vR��MK,cO�1�K�g"�py���F!L�p����V=�a��B�uPa�	y�M�g�������gffإ!h��~��oG��k����L����"� E'�U [e'�̟���$�r*2LR�E7z؎� �2�G_���w����M��yݢ�g�@�AS�bz��S)��ZӁJQ�`;��9χ}�-b�Qt�U�\G�4�L��$�7F�3�8��^<&���̭ˇ�MGCR��H�b]q�=5�դrG̖)3�g0�r�/nuW`�|ŉ��zp4�`�nhy�J�3�����b��W�M��A6���<�"���|C\)���z:N��ѝC]LQ<uѿ��P ���e ���j}jotI�Fm!��.1r�
�����޳�o�Uñ�*�����`��=ȇ�\�碍�F�L�Ùl��2cn�eN1��f,����D/]_�s�ɕ�;�h$�ie`=�v���\`��َ��A,����*�d/B�D�Z��0�$,�㇉��?4��9ϩc��g��;-+�ƒ����G� � Km	��٧�P<:uə[�*�h�u�L�����
񡕦;�6^�ƭ�x���xy�0�q0�\s
+�<q��pP����NY��A��B<G�Ne�]�o:�ܕi�+�[���� rB$�q�fa7�IWn�"�I�&B�Q� �I>4����:����������0���9�|�Ip�T��K������#�_�nkf2!5���Gc߳��������$1�n���sM
Fʐ�}-�^b�4��]�_$f���H�:�â�6G@�R ��T����')iU/���E��>7K��i�Xe��2b�c��P��a;�[]�Qd���P�W�ek�&����bJ(��H��m�I+���]�N�,���~Ǽyd��.۰�}�����Ae� $XAACʨҊ��Zb��݋������n���M�L��nC�����=��!���$�����%!�5u�L�嬻��5+�[����x����_���񶍲	�T+t���8Aj@ /# �QgX����C�g|_P=^�7�S�B*�Ї�f�ҹ"��υ��D���v{��?	ti~U����rpf���ߋ(�34 ������v�q۝�O����%�r��ux��e�h���T��4? ���D�Z��A��l:�::ک�y������]�ן�^
]�<�rAZIT ,-Y�1��,�n�é��E3���tͤ���bpT��Y1Uu�LS�	��U�e���y�g:�Q?�y����W���ۚ��+��a�Z�r�u �N���m� b��B�Wf{������? �|��N��6]+�=w2���v���HTg�����������p	U\LT����rBg�2�2�Zj��C��i��,�"T��yTSC��V���)��o9q����G%U����1M�S�)xI3P �X!��r�����&��P�|�ZS��w}��-�w��L���h��CS*�?R?L-D�w�H��"�y�P�Zv�ó�B;y����H�4��.���s�5L8n�#�7��pr���N�W%�k#�f�j��>-y�`�!`ٖ�%�vk&9��/+aWU���	o
��\g��a�N+S�D@Hw(O,�i��*,�);+�u�]|8��'!�4��Ww�Bf�Z��	Cu�XƲ�Ii����z�d�	ӫb	7�لG Y�5��3���%��Іfh5�������.ؔF��c�R|F�<%�#�vm�lʤ���|ր�p�;*p;�)��-��q�����6vj��}���GD�8�gr�.Y(���֞Jc	�94k�,!�|BjN�O���8� �1�{��}�v搩�g�>�e�n�*�h<��p