��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� p�X��Y��!�����j�V^�ʳ��*
�,���I�)/��� �����{�4ePs�Ҋu�b'��j����Bw�>Uug��q39�NPU���>��Q�~�pC���ڪ�- vӏΛ�9ȁ��﨧;�2p�kq̭��cɇW �??J���=�#~�$��"k��,�Zz���h�;��89q̮�b�d*6�5����Rd���S펎�d8���)�p�qfƻ5��Nj{c�I�����eTo�5��XIID����u�<	�1 ��!g�nD�%A��
Z-Cej`�d�.��oN]&s�����d���?�L鐩��ԟA^Q�vn[T�����w���sN%�H���7Z��pz#�t4��0w߫�S�'�]KJ���
���>��u�����u��h"s[:	�G��m�k�w,����1D��i�r�b��zꃯ�, viW����]��ɢN�S��z���E��aTO���5�NZ#�2I�s�J��s(P�7w��lRy'�<�?ӵ.r�ĺ�5180�`�"`=�h�ې3�n�˶O��F'�8H�I�)��]a59��wiﾗ�F�1�ZE�c ��ӑ�ǉ?�Ҹ�3F{�M���A0���_B\jB�Ӆk�gm�?s�k�p�μ[��i�����H�M����ZH׮M�՝\gU����u9�,����q���L�Z�����;�G?",	�:��mSo~�"�<H����7�<�\��v�\�o�@�a�c��ݷ.��])�VO���\���6\�G�P�w��'�Fr��� /U��^��҃�ZP_�[)l[X3����\�+hd��N�L�C&�~�]i��(&� .$�"6ku6�`�#�ec0O̙P���?��_pW�y�H_��r�E*�$$�=�<�"�SFW�ӣ�7��?�M�.��p�'��I]�YB����X��,{i�wz'��jY o[ف��=k�:J���t K�MҲXq����m��x��◌b���!������T��73����M���&�3��ә�l󞰱�����`EǤu{n>�"�HʅmK/^�ˈ� �Le�~�H�xO�Hf��G��w
�c�|j�'ɘ ){^�CAla�!��ߨ8��avу �������������
_�/���	{AV|�����/;�sOs�|��x�
�H
����>a��]?�B4�tട]�"��ߑ\]0��k��:�A=l�ċ��z���#��L%T'7ݺ~���2�j����ƒ�C��!�9 ��)���������� k�V�V�TL~J�{��/�U�,�o��i�{���+�?Թ�{�{l�܋�O�HF�Q`G_�NӢ�z+�_x����<ʁ0~ۛ'O1�*S���)�t���יr�i������V��p��4Q�+��"�>�=���'˙0��:]�#d!��nJdg�
H��HE��E�X_���������3q�����X
�0ek�����Y�N�C&5JQ���誘̬58�<-��\S"bD9BxAr� �{���6���<�k�C �)�`(��ڌ���Rl����^J"뚛>�:L���KpOd��K�����䟂��D�ZK�G�O�σ���$�oM�"���,�9�����N�� �+jS)
C�C�}��Hy��>U�#�6Q�GG�2Td�w�_�y��
�$�Z��iK�ΌL=*��gё�`vVd�2�1��S,�V�D�V�$�]Zs>�s1B�u�_ϣ������W.�?�������w���;���u4�������L6�*U�����׳<-�Ų�
V��K0*���ϥD�R�M�Bb}�9�S�����m%"<�{�n���zs���?��qo���Е�Ҙ�*&)l��]]���?r�����9}���*�e^*�a�U5��[�2ʕx��CL�<JC�K���B�6ҁ��q� NU��t���� ��ʽ�����O��)S§h�v{1=�y(ЇjRi~6�8�$U�+���é�b���A�3~m�����M���Y�&�\�]=���<��)]�'�k���J������k?�#Ҵ��Q�D&ǌn�Y=�&�jG.�0��F2�C_��WᕵM��aF�B
���Х���ڥ*��wl.[�t�JE<�V�qc2o�Z��@�'��պ��׿ɥ/�r��+�)ec��C��ZJQ�.^��)�޿�|	N.͖�Ź���DJ�@|�~�P�zi�w�>�)�5p��f�{��*�����G�fxc`���,Y	� Z�5\?�"X��[i�A!rWM j`��mV<�;L⺣�Έ�4��F�m�aM����^�>+��B	��{����`��
���#i6ݳ����B0C�}�fӵZ���V;�g�;g���֡���6�LU���C�S�V��h��U�I�W2�g�C�����c$�Y�
<7���/m�L���{D��P�sz�r���9������^���D+���tb��cK#��w�N�s��ZTu�2�/n}�R&�E���VU"K!�7�{s��"LR�[���!�BoMI���ؠ�&�6+c��);vy�{�4ؿ��3�R���*�s����[x�o'8����_�M�Aec%�޲g�m�b�����di|DK^H]�n��_����7, �ZR��u��\S�ŵ.L�XX�Wc5k˂LI�`�Lp"L�@�
�X�;�3wE��N�{�l�Xױs�gn����Vx����EQ_�,	mG��J/i��z�b�%"�y��H�|$�6V�,L��j�C�y��#�E�āH�*�f�c��7�!�:��%�Q�_M��wA�����2���K/.�-�W�O��&B,<2��?�a\�O�A+X	 d6F[_|k=��s1�k�S�`�:[_	�]�q�ڗvpջbTB[3|�Ua���}7 x��hПTm����ͣ�b��� ��gv	��?���d�]*�#�-�Q�|��\���O`*{�$�9r��v2uBn�� ���U\�4���� �ٻ)صg9��m�#���Q��tD��QJC��C�W�M�*ɕ0C����h;+�]C�S��]�cs�)��B�\9w�����uO�)����%!�)
:@X��c���'$�*��v�q^m����kR��*<�Hrd�N�9���ǟ�������dz?�"=LX2,R�<	g&��8�M�).�<ٗth��]?�F�J5���!_M�W,gB
�,�*��7���0�Ul��
���f-�kh���n��{�9����ǰ�P�����`�S�Q�Z*��J�գ��$0��*:�|����E�5w;U�C�B����*+��w$ըD+�&�$�B5�|j{
3�T|wx1��NɄ~�8���]��|�G:y�Pu��aR6�羾�b��q�'�A�9�q2�3ǀ����mah��ę��"���u�jfr��T���������d��a��09��YnlȺ*�Ua��AҮ���r�1���5F�b��l?����.�ڎ�t�����:�z�R��^,.P�M��U��Q���c2G�ZL�s��>��E�O uG߿hO�÷����@H�6�e_�ҵ���R������Y�0��R�joG��{�B�D���������
$��]�"
)�2�`7Q���S��>�ސx*�~���,Z��o��Jb�k��'�l �N�C�󷟁��%�64A[�1�%D�?{B��	�����29��S�?�+����� �׫�֮7�ܩ��ݓ��;b�8h����_�}�����ox�u'���}��=�W��1�4g�]�d.x�.��1Ch��n]�Yp��N>	[@��˰�G�Ƥ��Զ���&�̔:�|�a)��q>؝�U��$\�����yG��{p�ĥ��|�Y������Li/�����ف3�Eް `�U6��*�2����d�)�rr��Bzh���N[;f
}1���Q�1�$��0�`��΢�����Y�F��S+�*�1�o�}����:��Qo���.��A�P�kM��5B�lz�W� �jrFz+�;��g�w}@3-�\���e_��}PV� A�U�(�G��U}o��!r]Pa_�;Z#��I��ުb̮I��VOjlɩ-�=ae�u-q���xP�k�tmR(����@���s,,A37*�]J;�Y�{�C�������̥]2۞�d�T��=�Jj�.ⓣ�LewR�Ў��YQR�(ԣ�'(��v��;ē{�2$�����: ����"��W�A�Џ�{�UuGo��v1S���̞f
=�G�+��kescO(��s�N�+�f�0#�Z>o����-^���G]�1���!}fK��'.�f�?T��9�sB���h�H(Wd}�ht��#�3g��0��゗&qv�?,bİ��B�ObH�2�:ш��[�x� ���"�]��R�r��-���\�1wm|�FUJ�ڹ/�)�-����dB��nA�n����D�������/�s�Y�G�}� L��2čT��d!���$a; R2{P��
E��TZ������yβ�!�Պ]�0�$ak�t���մ��+Y�4��8�l�α��%A*-��vCё�ab�Xsf�V����<����; /j�jy�"S�#�|�Nj]	�e�Q `�CPӠ�4�M>�!���N
a�X�ν�5|�T��$�����%�m��8�H0�tQ-ԏ�9�x-h#�$��>��^���Q�����6jZʴg�GТ�ǔ��dE�;�񅻶�J|K�ӕk&~#n��&�{xi��_����ʖct����\_���5a�[��W��Mk���ks��K�Re�z�#�����>�O�>�Q[\��(	7i����]늒���D)(u`�Ⱥ
p2n�w|&�YX4��C��S��9Ob襇� *��S�&��.9n5`��-�d���w����8x�zQʀ�fo�j�VL��s.���F��ǹR�����p��4$5G��ߜ���7WF�+1w�$��1v�
$��$~8���|{�H���!�!"][�p�p��f�9���F1K3(�Ų�U� �D��%����7"Ė+�=�gbV�t�\"�+e�/dt���R1�S*�ҟ|���Ȍ��6h�Ab[���a���}�� d\ȁ\��^�眲�}JO'���VgL��;�$���̽H��s��|mh������LB�=����Pv'!������_��d��of�(�&�g��K���>"[-p_G7UƱ��n�VM~;�]4�4��`E�Qb�i �Pi��IԽ&�M�1��K�D�C9}�6_o=d�XL�AW@� �跬c�{���؅i3	eقJ�{�!�(C���F�s���D��c0��K#��V�ߗ#�K�EבB��y��<�,�T���zؒ���D�ps�����}��5Eu��6 ���� ���H�ɴ�}��ڽr��:o�u�<����@iT���E@=�	9ȟ�#L$�Yepd�rb���F�&�mlb�~
*V<r��w4�ڃ��N��VG,ǹ�T��E��-=���R37ͳﶫ�yJ�^�kw����`4s@���Ŏ�0��EȌ����M����V��)d�#��f9�h���^X?����B��ޭ~ �u�l	J8/ky� �E���&GV�'s��
y���/d]*?9��`B_�d�A�?�t{1�ۯ����}���W�8�g��> .*ѕT�Ԥ�e���Fo47k5×ӱ�F��{ָ�<�Ɯ/�Bi���$���O�M�bܶ:�.6�5�I�DO�3tGϞٙ�O�����=k�z�)г����J�v�F�� `$j	h~t�ܟ��#�	ܽm^^O��kk���=�A;���IN�����+ru˩���&ܸ^]47��F�k�"ܘE�sPa���܃Y0�+��s����H���ZH@C�~8�R"H�F�Ie�L�Eq�a��5������(����pH�ϣ�;ިN�� ^){q�#:Q��s���͋�� ��᱕T,ŧ� 7���Bu��SC�aHa��^|�2�3���tLWJ�$�Ѡ�zc�7|mZ
���z���|1��Al�5ŵ�u�S�6:����N��'���]�nʕZ��ۡ2�+�,a��US�WSt�ҏ�K��Mp��k-va���k��?]y��/ܸ���"�����c���#�C?A<̵�|=�;죱�J1��p�;3�?%�d?蔀+q*�E�1�����l����Z�y/ ��'�'��ίf�̸s�#���TCR~M���-?��.���bS�u�w�,��Q��o��\X��~W���K�#.�_�YPd%��b0�W�T0��B\��s���j$ϛ8�f�o;'T����[�DQ�O��p�
��<27�U��?{����*R6��2���Q�N��N.0P���dl	!�T|PԨؾ�)��_f�;~+�T��W�8y�=U��ed|f�5:��+���N(è�T��ev!���n
Ώ4y9O/�渢�p^� l�� 8��A+�*[�)�(�B��.��/W��%�ŉ�$A&b"�u����6�ÞW+yGl��D���)ǹT1@RVg퉈�ߧ���zRpe��yq`e��v���(���PM�:A�$���T�����4|1JJ�_�"����j�([��5mV��C��fjRf����D7RUo}�E��g�Q�|�};	�eM\�����������a�c��P�I�ػ"Y�a��r7��N$��~BV�PkZ��[&���v��FY�z��y'��T0+&8rQ�A�<�|�ge<߿��<�m�vH�4�߶~bZM:ڳ��K*^�� ^��xT'"�g�ic��c�H=!B]g�)�����->%5��o-��� 2���3���!��:<�M��'l�X�e��wfb����y����\>�~�޺!Ū���d"*-j���~U8�#g�T"�	��V���B�ijX�$#^4B$�	�c���-x�0

@<�4����yb
6OUxGDp���>�cS���*�%S������ l�(5�X�������N����W �"�̜;����ȓ�d	���� 	�J�&� /���v5z���JY�ۻ�U�Lv�s�Lnh��+g��'V�G?D�;�`�0��
]!�������O-�-����t��䥰�Ŏ0'���F�m�Ѧ(���g���Ѻ�% ��zN	*��î�!��L�5��'��k���򾭚a��c#TxH����h���}�g|��W�4��|����.����|�:�:<���l�Iֻj�,J��)s�*�r7p	�|�Z�A�=n��G�`�f��13��-؛3�'�j���t�M� lv'�'���鮒R.l��@�)D�cr��|�as�$`�Y]O��M���r�)����ܡa?HJJ��_1:\b�RI����n��9� �A���|%�7���c9�9��"�V��C=��.JIu^�{�o0ӲXO��N̋���F�� TQ�X1��>%&ҩH5�h�ܭ$ΰ�G�Z�q�ɂS��e
�32�iX:�L��M��룜hEt������غ� �:�Tj�V����D=�S�;)��Q�ه(�͠��8���S�"�
Bp��]�Y�G�ؚSS= l�"tտ���K���5�$V$v�t��B�:}k���inz���'�6D��(F��k�V��������i�m1ǘj&��O���ܨ��7p1� 1Z�Sk���f_�$m96F��1�z�$})�5@��S�`��M6���׀�%+r!�'ܢ�2bSn
9�.{��?��u�2�ޓ%���fH����F��ѹo�Ѓ����4�FRh2�	�ϨT�6rPy���ؐ���?[��c�)c�F���� �{���\Y�v�웢���K��X��ēf���3OVuq{z�]95w�� ��[r�X��rY�[�ca��c�dg��_������Md�j�w�ī1�P�afj4�1�x���F���R	��d��&뼏�u.b<J)W��;*�*�e��V�$,JT����>����r��E�mo�P��y��ġc�)�ΊcĘ��]� ���l�#��(͟cܒksAI]���]��a5gW���|�t�?''������(�+����J��л��@G�ġhM�ٓ�n�{~g�HB 8�<s����{�5�z�[���2�jF����I���lvolr�=��1�*�b�H�%�����j�0�0ۀ���* ׵�y(&]�syE����bO���{2�!�cr�M���)̈́����=7H�2�o��3�V��U��D�X���ȼ0�a��~
"�����|cܷ�#���|fّ�XM��;���ˮ��	6�ꪻԨI�|�4E^���X�y_��
KH*�_�%X,�K��q����G�>�������_�h *���#�>����~�?��Ge��'u����to�t�82X�G����I�������g.ˑWJ�"��]L�${^h�_{�0w�FhuU�6�v�Pf��E���o�@x�����Q�YG��C�6�{�0�1W��s^w�����F�b����=XZM,��?�Cj,������p%\8�h�������o����g�	HK��2,}��Q�Cx�x�åX�e[�6�	�X<_�#ۮ�;��/"1�6a��Q�~9.vॕ�!�'�ڂ;R�:�P�G,�P}1�}ח.K_2��{ ^W��j��3΄�N˚�5Hr��v~�P�>�'�I��B��;��{�A�fH��4�#ӨC&�a`��U�ۍ�����௧V�72��v}� �|t�����"����A�mB����D"i[���	����e����r����сKk��ї,�5����1��LL0�A�Ɖ&WJ��0%U��(?Q/�x��jlw(#/Ӥ�6��d�41=���IH5����;�ə;�_�K�V��X0�P�56�^G���X�}h�;+�~uk�Td&�H��B� t�M3�=��0{_\#����*�r��X����Gn��b�	_�B��բq���g�CGp���aHѲ�7�CpX��O[�y[��y�3��d|�C�i.���&��M�!��bqG9Q�t ��2��?�6C	VK�#�*7���!	�$��OO���-�h��{	�M;+��k�}_iƪ�#<�2�{�&��&����N�h񜋽���+e�§Y�����#U$Q:(C'2�'�<oSm��Su�����f�6bA��4�ǍJ����6_�[�@��� mL������.��[���a¡k�GVkA*L/"+�)��1K���/b���)��ɿ���`�g�������o�!pyyC�/��� �S�
撚>$� 1����Z���A�sg���`o�:�5|�4hTqD��J�Wg����r*����[)�1V�L�����-���)�'�hO����M���d��̟U��&Q���b�6�ǹ��ꠌ+}��nn�qk���޵�I.hq��+C�|���79��_LE�-��\L����f�Ͳָ&�`�zI��n�˿@�_}�%S5���~}�L	b1��C���y�ڇT��^1�YDCt�H� ��Sއ4���V����35ruh�	��B��$C�I�HPh60x�_��)��6�u ǿ��o#>�R�	K�*�~g�]7�[Bf�Ƌ���*�E��5y;q���j�=�O\���d�B��d��?��-��N�U�� ��<�e���
} B=v����7+I:���bP�\ywlYp��+�{�	f+�?��V�,K�{�I��EXK.�c.���0B�.$m�Oc&��0,��	�����9'�Q��>�Q2D,
/�h���ꊹ�o�>����Q���	q�R�u����f��YZܡ��+*0?�qF^,v\c4�-N�bQ�������I&]�������d���!0Yw֢I�d��Ք�����x�$K�~L�@�<Y�A�� �{:���`��O7 ��!{�!�tmA�y�ke�!n�%�,/�	�|	),6�U�;������x������st��.� ���,e�0̭�����=���"Mu˶�-M�zG����<RyX;��==tAr�1b[vYB���u-��+�R�[�H}ʕIJƣ��]�-~���?�<DLш��L��`^Ɵ�!��&��i��r��k贞t�z�C��Z� R
�&�U�s]�m�?��y�J��4,�Q�`=�B���
��\h��M�c�t��$w���ӼD�xȩS8yӖ�(�@��ۻ�`Ғ3暡���NU`��Ij�灇~��!yg��Mc��I��?���fm���/�ռ��9�T@5N��,�׈���h�|'��[orc6h�ޭ�ݬ���m��^3 ��e�������v���m5�s�s�54�WI1�M��)=��҅Ɠ��ɹ�Ѯ�뤢����	%��^7I)����������:��1U��<E�n=F*c�8 ��-�C�0,��l���rN쌈{��P�%Ŵ�V�p�e��Pʶ9�I�&Y�36c�Ҟ:v{� �}�Zt��ݽPc���]�N�H�����(�9��K�W���"E(H����x��5g
}2/� c�I�j$��jt��X��&{v騮E�Y��p�g��>q�Qz1"���B&	A���<��/ڎ��v�[�����kB�<T�>~��q"��N(s�y��qfW]3Ǘ�qC#nb�����ؖ���Ҥ1&l��`��"ɠ���?*ΐJ5Xa֛�6&�;}��t�J9l�����c��q���j����H$��%�׏�"�ع���W��F��2b*{��ȯ6�A���H���7�����i(t���5^"U�( H�슚vG�0��)��ε��vx7����Z�ȉ��d����ԟC�ZU^� ��
6&�9�(m���T�@������>�(�m��_T}U3Q��_KZ�="'	�?B\��Gn��'T��-�-�����8��E��;���[�%slIC3��
�Cp�4���,�z~nzߔ���բa�i/�]/��^k��� &E�/� Zc�������#:2W��%Nd��ͯ�U~h���c �K��>���FL����o�ި���\}����j���/n�դ��'�A;�!�B�X>_��lX�/�j0(N��N�=C{)�d���?
�̯ԗOA�/W���eF^0�v��Yu�]͛Ƣ7I��Bk�z���V�1J=U2����÷Wxnŗ�rz�P~�[�ɳA��S�e��pC�5�K��$�K��-�W�½��	"���|V���;NF{��]����}1�H��ƀp�~�V2ep[x�wO�3>�[����%�8����m�0�hƷ2��N�d�$ח�GcO��{Ɖ����%���=�G��:*�����>�1暏����FFJ�����Y*m��� �{�/	�b�q�LH��W-ʮ�<՘B���Iإ&7��R��Գ��~���g�18���My�a��C��N���t����l�֕�Px��O�Q�%F��L�qL	�U��
ٚ�?���C�Z�	�����2F�)��7��NT~k �v������2����=垟J�sV۵c���g�k��1��WZ��	h�Ƌ
�ރ�{�Ͼ����bt�����B��S�E�?�9�/��Ed�����{�%C�30vf[��*!lXH��kєy>)�fʉ#�O�{�OzG0������B�_0?h��2��/��3��Y�P��\3�E�ښ�)����Θ���8ɅZ$?�|
%���.te	�'��}��=�j�[h�1��=`R�7��T[�ӵZ��4�������|7�f��b�L<N��YL�n��Ò��� ��D(>]o_���ۿ��~9�2�M�"��pN���C�VNx�P�e�%��˞�ၭ%iIc͟L�#�;�ᨁ[-�9�\�n��SI�CVxoM۰m��M���=�ٴ��xPb
��dV�������Þfgj�>�̧v�D�ZT���9�g����`��׷�����&�},ږh�o�:��n��ۧH���ΦxUR��u�{>Iw�8U6���InP���im�	��Bk�i��r�!��΍Yp����\�O�u�C�I���FشpaM��-��x�c+O)�n򼞹�����鷁$�F�>9��'�}	�z/G1�r�B���]9|�+޾,��.�Rt�:v<�Y�5QN��7��(���p�	��e�q��u���./��֝��&J,_� (������ʌ�?����7�:����6�~.��������G�cv(��Us��9����_�w&����b1X��^��b*���`��P�.�'�c3T�C���Y�jՌ��i��v�.y���絽bԡ������>� �>��7ռ����}7� ��������W�q'"-�AD7!��z�/��=da�Q �egT��?_��-��͡��M� ���֨�RGN�5s]��)1���z��d4�(鉭YC	a��U銟h�&�����M� X2b��+�n�>ƃr��T�$
N_�n(��p��RR�,9�UN��w܄� u砺��2�#��K������ǂs�t��,�;�+�1\F�]��E�uv�[�-c"���VA:*y$]P������
��8��6i�;��E�_�҉��TY����ױ��s/��@q�v�~�Y�QK��*�;i!g��]��z���͜�>ʱa9���L�Ƽq�w�#�?wQ�-�ƀH�M��Pd�u��Q-\ɜ-��!D d����伨<�+��pu{я�V0���)Q���� ����p���?
��I���냞�*i��L|��V;(J�]B"�`�щM���p=B)Ip�!VÀ�&��0\�rd������4��'Jޮ'�El�g����.=_0Cp=��g	�2�	8���}�*��G˸lZY��]ϧ�lE�!�{�v��S+*E�]�kTR��� �r�W�o;TUXi�۾������#S
�m�L�=T�-A)K=��k�<ѝ��k7q/H���e�p��Xi��7:;����eC�=@[Ʈ�@�`�r�ؚ�J{0N%�(��;qY\?T�.�!93�֊�^���:���K6'��n�ºf4"��:k(�R�p�l
Y�ϫH�7˜�9k���o;XM}���7̌+���I���+0J�UAp��i7�!s�ۨ�r�pT=��Z����=�D�]�V��0�#D�O���kƫ�����}cN	o�l��r���I�6�������:4�-D)��s�j�
���N��"�ߝ3A���0�T�lM��wԢ��8�y�	���G#�c�4Q��@���� �]�=�:D�p�ˍ��c���E��LP���"���rj�°i�}8�XZag�.B�TA[�.��k����d,5���]��|H�Dp<�l7�rSe��2�Fx���OSfÛX��lCڅi�ޕ͖����t@͐jT�����;���V�b��8b�w��/:X���_0�Y�;�j�g���˸\�pjA�H�)��$��霸��nL��47�x�������3&��F
wy�'x��8�艰��l޸�Nr������ݓT�67&X�0���gjN��@�W�J+*%��X������Қ ���^�S/g�1�G~�;�s��!ش*�44&�Y��"M��"G�H�qw��s�$Q�>�j�|S����Kq�ݾ'�U�J���D�"b�7]/	����iL�e�:���/�4�����9�P��OybO���S�pAZy��'Z�L6�6�F�֭�E��������	�}�7��y�d1
��.�:�R��k7v"�N�Ht�4�Y^��X���fr������2�7��[������5�!����o,P9�,d�	�!V���kj�58-d��_�Y^F�%�_��<I-�~�Q�a�S�~���\�`��$*�(�gUI���ǌVP3{�ݜ�|j�n)�D1_UTF���"��Z�jx��Ɵ���Xnfu�|8=�ؑv�����!�m�8���J�`B�z9[5x剌=�����J�C��;�@�Y8���p�ׁK����A(�v!�kj�w�v4�����kx{  W�]_ڝ ����������G#��5�!&kM���SvG�Ď��"�I�箃/�3Ŷ�&����D�sybW��Y�#�Ua� ��g�n~�9�u%_��(z��Å����l@u�T��z�#RHD��L�T�q����J.�fF�U�^�fƚ����W	f��=����}}[V���ܽ�zJh�a �"�QN�,P3�����aw  O=�}"�,\�� K#�?N:�MRx'���?��~�+�:\2��"�&���\�-j�d����e���pI�U��LQ�X�I�;
����źI8��s�ގD�
�|_��@|:�v`1��%���E�}"��K}az��1b���D�w;����p�^��@�\�����͍�|�s�i�̌w՛��/]�E%����mj3o��Uuy�;�i�#Z��JK�P��~6F�`�1�{�ei�l��$B)v���}�\K�	�,J�=�ǈ�V�"]���`wv��@<��O��QNV��CH�Pv{Bj������Tk�>��$�l�>0��D�4�ް��7����]7���0�'�ٖAN��譚�H�UO�h�璯�#�GIL��^�(���;�)
�m�Qn��1�N�k�K���9w�� � R���#T�G`BB&q��*��ŃN��UQ���5�`�����F����,n�!��5�Q�;��ss�+�b#��W�q��g+a��N�C��r�B�C���̔sMs�'V{C�c�]	l�ո9�w/*���0�ְu\�}���պ>���ț|�D, ���]����X��&$x䗷�V�Ԓ	�PD;B��*N�
��{���Χ�I��Y��AUՓ1�%ph�'4�'���ퟪ5ӏ<]�icͥ{5��2�J#�Fo��;<��\��p2C���6lB��ǖm�Z��ϫ���re1P�M8��s:�\�����1�	��vk��Q3��G�DD���W��p����Y�G��c�x�yŦI���x�w��F�-O	�����!�����3�hWķJi���W���a� ꩚�O���l���ѷ"�"ȓ�A3��%����#�d}Is�~߀ͺ�?UY��pJ�=��?^�:�_y.�cY��m��S���Yk*
�O�l��,w�y��b�����v)7B���7{�nA3R�"j+���a�������1o��=a����*�Œ�nW�-7�j���e��z�M���߿��O���7�Mrc��Bi��D����<F<2�(��~����
HO��Z*V��[���y4�+(v)�k#��סC�������ZK���>�;:�������@���2�� -s�|�L�ѻ���G
�S���5�~֐��7b�%~
{tDV��}X�q69��H�;���VǙ��k�h��32v�f%�Б�$�uS�P̀�<��'�Ӗ@�C��R�H^��+1�������-C�2�?�/�)��(�~�Jq|��I��q�����{�
�
��ݳ�6��A��N�5��Ж������׮eE�n�1��W�o���
؀�!�d���LU�>�3�IA4���:H�^�*�8y��[����AA&�*jуJ�'���62X,풱$��L���'���fqj�"�b����2�����p��C��hon�� җ�<0#(D��g�o{}�C�m�p$�U������ǫ��@��-?�g�̑�?��O��lo&]�H���&