��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��GN&}��>�Gh{2�EeM�~���=	�V��Gt���7�.g��w&��Ț�)�����O:����ߒ�՛�8�x,��[t�t���V�o/%�������e�"��T�U���ʺ����B��Km�fq�TY'�����������yR�'n�[����,'��
t������L�2�)m:q�ⷼ�H���*C0C̊o�5?�F�;��
��� ���o����-x]��4v� ����zVC"`.�� �+	�&Q�T>�>ɼ�-�U���'&9�&[>B/�M���<d'm�D�^K�}֜��nt��2� )�9���ĳ�~D����*�0��DV4��	�<=��P����)�,SK�����9\����J#=��}�rIHyXK&����)N�|�ڝ\VI$Z;��Z�]���D��ek�M���� ��2��Mҍzw�Yp5�Y�%�	������ϻ�U�4�����h�`��ܓ��'��C��U�����$=Q�L�󦣑H\�6��?�ooh{���ʄ�]ʥ���:�H=��P&#�{��i��w%�_P����ɑ��i�mt�Ϊ6z]nk����o��D_&�x�� �}�z�dT��.4�I�8�i��O�A)�yh�1�M��C�&@��0��I#��7UZ~����l��HL���X�I�.hE�4��`��յ��		�1���6#�����c�<E_	��g�s���mM�U������`aZ?M�oH�v��C�
z$(c�-������18�>��C�����F�� mO�7_�7ʚ��/���1 �eAќ���Z�	�G�
�	��i�A�y�bw��~��f@�
*�n�?��k?]��k����I���˼�\ ���o�θǖ��w6���}y]�Sx���m>|�N������A�ߺҚ6�5�!m��B	�8��X���/> z���q�>lC(�����P1\.˫�9���ٕ���7_���+T�X�a I�~�A��T ^���n�a�r�k(��Z�?hR�9��)��'��;��=��2��jg�P���/@${���Zuv.r�o5;��3��`����12	ZcCb�So���M�/Zn	�v�����Tl]Et
��M�eQǢ�%���,(Ruό'(R��|oى��HT"�����</��1t ;��0ׄz\�kĮmēGq"� �ѪI�S}(���#��w�c�$�eZ�s�]J�S}�-7��!A�����Mʴu@^�t���|�	��N�H�$4�� CG�h�a�{5��hq�mOq&Hԓ����]�zD� 79����TN��N��[=J��ڨsQ��A�s�����Nf	����ۼ]}����	3��D� �)�(�Ȝ��H\�*�����EǍӉ�6��o����Z�n������\