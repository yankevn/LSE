��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d�x�%O�ٵMro(�t��),����z�}�ٱFq{y�����f�y�gM��0��ߐ�䉽�<P|]]�ϘO��S�s�u��$[X���ޕ���2b|9+ gC��*��ve�9�	�`��2G2iV@�"���w����Yk�^.S@h�5�;����>���'��4c���5:������NP�Ħ����tV��C�E�����zg x��!߬P2Ѓ5�����*S�@���ɹ��f�I��s	�y�}�3�מ	�$}��B�T ����ܷc�^��9�P!�
V�q�e���������h.����������{:W�m����yq��$c뙬���^4�fh�-���䛼$V���4�&��n��u�h� v�(?��3�l��T
S�����׷��s.aG�bpW�������9��Ih#52��S�;.�#~��r�2�.g���J������)qJ��Q��yɹSj�(�o��U�[HZ&ܿ�:uoܨ����Q��>,-��p����IeA�U#��xh<ky?�S���>�o�«��|�s��Z�<��%
,h4�ظ��\�z"i+�ioM�h�c��X�U�{� ����Sʓi:����� �q|��N�ܮ�-@�W0����oq�u��X��� -ON��*M�xQ�u�B$|ԩN�3=��ΖZAnA��R�mB�ק�����lW�}�$DH��YG�(Ee��(͖:#~̍Fܘa���i�B.(�?�VG���n#�Qd)�m	�ҴK�f&��`]$q�⭹��ZH��p�tZ��"�d����{�A��c�2�IE	Ͻ���_�� w
x�ǝ���+���vd�!e����zFD'�$+7���d��2�"8�;�0"F����:�e�{
h�����薷E��ɍ�umz5�DQ�hb��(���>FLw��F�O�����`��8W��/�s!�R�t��K��<�h�b���*�Y�W�c�3*�����~o��C.n}	�I:T�"Et���:�^��߁�@���NW���74��)/�X��w.I;n�[H�U�M�����r��Ć���fzy����od,����(3.̘m�.b��[608��	���|	����$�]B�Z2�Ux��Q����.��7"�:� ~ͷ*�����5(�T�7���Ǧ���R�-�fպ��: |Ba�)�-�J}�xl�A�4.�:[b�o�jӞ��^1E��t��!Ƥ
X��� �����m�9�����UE����h�_�l�M#	���` �$���0i{y[<h+s�K���-���h��^.G�w��ֈ��ObN���\�D��3-�tOW��lG�m�nJ��Q��5K�ELgߔPM�>�N�qm$	Hf(���>A�(1��gTCz�
ә@,� JVp$����F���]	ޜ�n�`ݻ'i�
�(� ,1�1�-��:>�`C��l�=v ��-k��wV�t���Nw�RQu�*J��t�<�1ʠ!x)�e��{2��E¯����L[�`
�^��I���[�@�:�\:��]i4�@ml�i�gA>?������F�|�����B���X��_���#_1C�����}�������G9����t�:��ܧ�UK��W�U�Z/�  �����'W�^[��'T��kYʵ��ӴY�cuD�	(+w�'�����؀���E�U���E|��"��F�i�}��^�隂����b���
���|A1�u���!�,�G8y������`�5ёg�,[���D=5�Ew���T�d��jC3`�V�z
��&5��5�q�2�׍JN�D]#*CH�f����������g2��J��1�
Od������-O-W�PSU�^i��{2h�����0\^v��t( !�P���YF(���kx�	����|�_�7�L��:�<��Z���k��!^�	���*��}��ŉ�r�X�o�b�������`�8��msY�wadI޶�����s%2K�=^��%%˅���SH�������Iv�����a3�ve�������#Ƙm@f곒���e�`ws��Y���ų�����V[{k�R#����!��W ^��&�?�R*�Mf��<O��SH�J��O��}x�{�tu��G<�%��NS&V�T�����g�m�Z80��� M��Q��� @>H��Caɚ x�7_�)}DI��2�k��n�p���W*�cd��<U�A����y
%f��^x�C��b6*�'!ý[m��6��:�P����bǺ�#�.�9��`�^��Hp~��[L*$��	�|��T����>���ox�OY�wP�/ɟے�	�Dǚ��х�C�$��a��_��)��yU�N���R� 5	(��h�&��E��7�V&�`5��B�8a�G��%l ��`����N��C;��^&1��Y�߮��n
3��[��k.��mw��-pq��,YR:~�}M+lxe���5�fE,Z+�:��<�A[�<�䕨ޖ�J�AZ3���&
�����2��+R�g�n�"UZ�.<��͟,����o~�s\d�H?�W����^G�}�Rj��8@Y2nH��-�X@!�J�qX7�`&��R'�i�;���ۚ�>?�)o�N�Į:Y�rk�V�u)l���\p����$�u���cݢr�_5vS��@�p�E�OJ��l��H�8@�.���R����gQO���\�k28�䰊FZ	;�ܴ��C�K���| hL�)��>עL##� � �2~`5
�����סJ��ݵJ���R_��6��mi�w�Ru*�lD"�G]�@9ݨ-�hﯘ���OV
�A�Kk1fa<�N���"g�8�����K� Է-rF~ф!�����U�/}�Sܒ;�A@�Y�R���}�Ӓv��	� ��C�f��}D#�8 �ƹ������h��@��`z�hu5�+j��[Жu9� ��GG���?,�ؼ}_afV�J�&\"_�W��QM�F��$G���l�
,��V��^�i6����r�$j����;���p�|(��F�v�_���W�����=x3@Y��4E��o��H)"9剕&�r�<�}��/Ӊ��U�/ �繃����l��~��u�н56?��'�k�;�%Ȫ�h�N����ҧWe�y��6��N���Q|���$��:��qU�B��Ǣ	��[��c���H�9e,�>z'�YMI�!OU��Gu�=v��!�����]����Hߓ,����65��\F.WƖ���'����X�(��6���f��������Q=���~��.��/'���W ������*E������b8�/�Rڼ�˙����f�!�6J@�
��4�|lB��Z^-#?[^険:7�_9DS��r�l����owT�r�+VV�1S�o��'-����\���0���M�Y\��U�IX;g�	O~=��*��u��A���Ψ|���N)-g߸�j1-�]��eۿ���hrb�)�"I�[����l���q�i�lZ��P�X����̆7j�r�ք4��E�'�]��t@�5�@PAB��9�!�I�@���9*��]��\[o/���74�L�)Z��Di�l+é�:B&���nWV-F�7��M��x�#���y�n��(^��S7���;�u�gGY�ڬ�,W�5�<��I��5�Ee�_< �����rCjZQu6�Y�`8�s���L��X��t�ͨG�������R����E��wqN�┗h{ �Ǭ�hYW6&�w[�E���#�h�`�)_��bW7�w&P?h��<L,2��@��fx'�!Dћ�GE���{��#��z��98谻�eY���\?�L��*f�z�9x%����n�]�
A"#hqO��$�6�j����E�\~?XS��[�}��
!�<�Đ�Ѱ-8�g^��5�$�_J��MI�������Cdth|��g�}�&RE����E2�R�`�RCtd�Z⟇�M`cNPw�U�=�@��*	���<A����u���a���;
W%XL��z2ٖ<�y����nk��>��� 6�ޮ�3������O������r�J�;ķq�RQ���A�~j���M�p����j��ZFm��S�fUŅP�m�g�o�Zq �s��]K�G҅��)��]�`�X�A�5:�F_R5kǨ!�H��&��	b��Y�0w�C˝(��6��Q>�uiu����A�?*����?Vd�l@T��n��#����9xD�ƷV� {����늇e�ͩ��^��#���'��C�mi,�����`=Q�er��� G�KIy�����_�!m�\d^]�U"�R{�TK���\H+��?�ޕ��G��;�x�1�, ��K�"b]�z>_�6��ƛ��iR�C��_���}Q:���1Źk����-�/;3��l��	qiSoC�<\��)t�xc���T���P�rD�&4{m� � �\J/�Q��h���K����\n\�@u�E�%�ɩ�z��|��7�v��9������9���]��V��=�4}�������R���E�¥�~���G}��y0+��@$1��ι�w�����o�d���U_~i[�H%�;�S��p��t��,���{.�d��'�vjT��e�"��j�p&{�20>��/�D)�����HRR�\UV�~���a#Eȿ�Yk��{�7�Z�5��n���O��v���V%��2�	�^G-O��|i�F��|ȈV�&��|Gq9�-s�By�{5���9m�S~�p�G�'�H�g�E�E��l[��g;�{�e�����`@u��h�mt�)�W,��������6�6N̿�e�8CpΈ-gڿ=O��r!�N�R=� H�Q	��	A=g�3��w�c���*vsPv��C�����F�����2lD�F�/,\8�e8�'����.G��o�2� ��v0���o~P�]?=�W�� :�����CI��d/�],A�e�Ͽk��+��^�p�z�۰�.d��� ���d�K$Nς�)�|����}�K6s�WQ1� �#��� ��W�����]��G\�T-r�}6j��Ģ�Z�3�p4��
i�ݑ
%�=�º�\�����2R<�#\X�j�SU���oO/�d�%���p�$-\�� L����I2�^�|�ğ"P%M͎�|�-��6�\�+�m�l��Ҵ������u�l�9��b�:oM5��n� 1�V��Rmwc3���9��t