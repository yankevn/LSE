��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�.�TfxJ<ȒEb�����X����E}'RN�ݜ?���B(*fP��g�n��(wn���`NO-�v��&ŉ�G��|�n��s+1�z��0�!��|(��� �Q$	�sT��:�+=Y�i�g�z{kҨ����=6(�r�$ɶ�g��Ó&�cta-Յ�`lR��b���m�(:e��<���;w�DX�:8n�65y]O��}�j�R�Ⱥ�a�:z'��8���Z%i]�!�zaK���l�0)�r���p-��H��X�I�}�Z�D�?7�l�$Df~5���n))5��dgv�IǕ����q���6��5�m�=O`I���������c�xt� � �(�]��^�J���v�H�I�9"�"�	\��_b�Š��v��p\�����������p����C��� ���ז��(�?����e�";�6���3I�ڂ�����{�f�ɭ�a{�֯+�] '��ZS�¬rS��  h��ʃ4H�K}}9��('S[2в�_ǵ>|s��N\��J܁X��:2�Pyi^T�o�f��:��[$�nF}���ⲭ�r��Mf9)<iDEI�Szc�ۺ�fըl��-���Ɔb�b�D�"n��@�A�?y ���tk�z&e���C\��
��?�cE�<�R
���E��8��OD��o�%dϞc���<k�ߴҹ��~!HS ��sc�㟊��t9S���nFec�PV���>0p,��M�=�[r}%.���)R�����Ў�*�� ��+�v�q�ٙI���f؛�>{��1x�h�Q��@�{��\��R�!��y�^�ۿU=��I�NC j<��u7�F���K}�����0�A��gvl�En�^S"9w��:˻�{u����]v�YM���k2Rd�X鞊$��/�
�T�5p��~>�`����@��� �F%V.g�SI��L��E��y�2o��}J��\g`Q���zpGO�׊[�6!Ksm�m�Q�+�~t5O�e���x�5ҫ-�4$p��t��p!�g�p�� �
$P��x��v�����Wӑ��C>���xX-v�<XI���������;�_��2#PtU���`)Hd�ܗy�����J��{<�wS^?�,��o��|�	H=���'l>=Y���&Q���G�"x���^�-~Z(��m��Ed�sv/��߅>W84��B� ����O4$8�Ӆ��4�QuY0�/@�\k�ˑH�.���]���5���+NbZ�E?t[a�@+�?[�bպz��Hʑ��C�H�A-�qv��Sx�C����!��}5�=(��p��?c�ú9������d������ޞ@{׏9�(=�C�n3Щ ���A8�L��84��^g0����{V�Kt|N���}3e�L��t"@-�Y��b)s=� EƄ~�F������L�qאD�ps�����ҕA����&���Q��g�K(^��/������+�F���o�Z�N��^����6hv���<��gޭ��,���A�ӛ�}۬�� �����j=*w�����{r����_�*|Y{��©\G]8PG����G��m��n����BG����I�H�!P���l���~�b��K�W�%�")�
%l-8��\�R�$��`H=iK�/G1<�fr$��;��j�ΨE���M���h5�*]�HҀ��8�����E�R!6,\,�%Φ����j�.UzN���;d����Kg���� U�0�\�-�$@�S: 
�n���SM�d�%y��w�}�M�	4yj��4<f�ˇ�
<z���6���P��%�0�E�~�8Dl�d��k���[�2�չ��m�.����W��$��Zz�s�z�*��I�ju*�HlL�"S��-�@~��
���yTF�ԃ��uxΤ��MP��b#�o���q�_b�wN�Ă�G��<�g�MZ�n������+��F](r)��UӰ8��sSf���/p���F�!��n��+s6�;���_3D�y�P�f� }�Ӯ�4����RЭ�ڝ Y�B-f� ��]�wy j5#G[h��Sc����]#�M�p'�0r����]�w���<��8��q�=�%�Z=��R'���Mn���x�b5p1nM�l�q�-8�dg�9��>��� ge��+�WYД��g���DT�GtڕH ��
���S�2�dژ�?�[�����B@������Lo6!8M�B͋W��Z�ΕKI?	{5�;)�.~�y�`fp�M��}��xKOW�c� �S!�Ħ�.�F 1��ӝ�$.�$w��eҐ}��F��-^2�[thKS�pE~���Z���E����O��S�5�yy/Zc�I=�P h~	P{')-s��?��A0�% Q=��}ї��0�#�$$�h�gl��.\�[�Zs��[&#��l�[^/����S϶:ï��_-��
�M��T���[K 	� ��J|�1�׶�C�Od�s�)����+���o,J�6H�D&�v)�A&͏�r��0#��+&���=���^^dn�/Ƙ����y�b/sM�sml��"�$�����9�^�䝔Y��V��������L�e7��R����!H:dc���@"]'D�����\k�r�A�H�v�w0i���I>Cԡ�H�GF��W��`uvX
ݺ�*˙�A���޹���ЂZvE�k����#a�^X�_����	to�K���ǣ3�''�����{��(dC�����s��IXn<��OA
/���:U����nYt2�L#2�)�[g��q~\I��Z��̂58<�U�Cד��KѾF�ϋ��d��[/J�%��'v"��e���N%c4��,�� ������0n[�+n�u��H#�g54Sw�x�\1(g	�Hւ-�A�*q���{Xw���$���x�>c[���ZrS�t�^A�� q�~��]d���>54��3�W�Ϣ�����G[�r3!L�*�WQU*-S�{��ӕ�P��^�z%ފB(S�����VZ�.�az~�,� {�M��i��5ݼ�Q��:�>�o���Ӥ�_@��\�YfT�ZL��-�ߺ�&��(Vv��~,_Y� �NÃi�c��Cq�N�=lq9YԈ5���V�J���J_{@�fC��0u����b�Sףu�r���Qqc��R\k��N]��)�1<�R���gۡ�}鵱�5J��m���B��J�I�u�0�3:ݗ�2*�پ������b�vl�`f8n-�bA�.�4����c5��'퓫�8�l��Րa�Y���r�ɺel=r���
�w1�;=��-r�����E�:�o��E�g����oޜ��~�F%{,*L_�=L�}��^[R�l����|������٩P�[B�F~�#��J(�x�MQr����`q��+o�����"P��\�H;~�H��B��~�^��tt�*-	4��6�J����w���W����w,����!��Xo�&∋L�q��u�m���ϒ�\{�<�G�x�T�6~�����*�v��?w,�$/������! I�$��AN(��s�X0����D���N� {x/�J�e}�g�����*���O�@P&�xa"渗l-��	��+��� �K�D0`�3g�����sS+Yv�L4�^$���Y:�_�հ`��$:��F�hP�?W�@f���^�s~$rL���Ԁb�n��A�*EW��@=lmbk�pKIn��u��_�Y�_>�'�4t�.�	B^N�Z��E�����+#�7�v|�����*���,�޾��w��[��b���!|����KO�#�{vW�Շ����d�7iR�i@&2xn��g������kEptP����HmA��⋩R�J����*ۣ��:Id�-'e���E��	���5��P{2�k	�@л�L�����������W�MeP$�&h�2�q�ٵl������B�_��������S)V�dxeX�R���io��?���N�!�b��F��bW��*�L?�郿m�n.m��iz��7����a2}��D����9Ӽ�8�j) %&�6{�����Ԡ��>��xx;��2�{f��´"(��m�`��`oNf��=w�Q&0�.�L��w�g�}���>����b�x0f�U��kf��\����W���:�hm���wp�Fm�g)q�b��̞#ᖱd�eW�!���>��}}�b�����E����ag/Y7�eWıB��]A�3m$��E��	�:Ǫ�1�3�ǮzP���8���`#sb���T���Ǻ5�����0��(���
�/Nk��OJ�{�rW�e Y�eo�x�;�6S%��c�����%�?���y*g2~Pk�%	�P�25��#��G����II�՝U?��L��q���Oz"���~��=t�8��+TyT|�
����Eh����X*I3_'�h��B�PfR�Qּ�@--U.�_Zh�9Y0���	�Q?n��"���l����Uޛ����*�]q�����޼�ʵ����<���D�5��S/��(qd$V��z�3Z��1�v�$�y��tA:���.����{{fzRwB˻����.#T	����J�2?�=	���S��/#�ܼ�����U:���~s~��Ng��r�ޤ��b�y�$����&�/ �X���
��dp�������s��K���݇(�y�+~T�U���Jӯ)�{5���b��K�����i���(1u,�P �p���Y� �H�M<��3GVг�Z�����%;آ���ibׅD��rqCN3^Z���m
n�+&����B�$�̖x�����5Ҝ�m����ߛ�W+[�i����t�pYX��o;�iwYL�Wcd������S�^�='+���� -��+�� "hd#�X+i�cì�i��K!���L_�O9<��YK͐Fd/ܜ��IݢטJ�jI���A�kf�DH0 ����W�o�CGX�9!W�Q����n#�A�{�4/}�U���*Z�0�R�����vٲ�>�Δ��-�;Ժ�0G��^:N����KM�}����+� 0�V.B�JQ�"��(G��c�(��
����04��/H���$;N;v��#�¬�@,�W)˓'�%(��n�f��2���b��g�_bS�I�l��s�3<Kе��r��}j�up	Ig�y�FZ�,�Ti��(���	ŝ����h�	,a���%'d�&��_QG�rR%�a�J�Q�&Q�{o�����:�,��oA�*A.�����gхI�UA��L\V�$)k!�B��q�y7����F���)�P1/s[5�A�n6�ܔ~t�W)�T|��
jar�3+E|D4�P$�#��&�l��S]Wd�ɤ]O��⌊'� ���Y�iˠX\�B(��ϩ�5�e婼�~#�,�r ���2b:��*����,����['p6�0�GY�&���`��
1@U]����$l.F��M�W��k��������5�7�P
�XM�}8
1�B���M�t�)�x���5䳁P�s��rj[tl�]N�I�!���	~����/��Z�U0"����=o�:�E�g�#q�t��tһ��U&�v9z	��1�BHÕ��mE᧵T5�Ϟq����D�, �;�#(��v	S�D6�����8%��t���N���p�m�5���ȵ�ك*��y���_ܙ�pd� B`{L�~��C��iU��ug��4ox\�����ʃi��oyIO�U�!��}K�UfC�)�)��,�>�ЇM>n���HL])�)BE�W#��aj�N�?�W����z�^���J׎*vv�M�;�^�Fo�Q/)$[����9{~�^��)f�}ϧ9x����]֔݇#S2B
ס����|�����[���J���z��`s��b��d���y`D<=���0#I��zy�僩:�=��7�)��N���3�����'��~��� �ZK�+z���x��~�!�Po\{Z���:s���ζG1��;Z	w�ɱ�!�/��ik!�b\1�,(5�ˤq�y���/iDH����k�U.�B5:-;�$���ω�w
/5���P��-^����bb����ҽf'������3�a�g���p�HB��Fi�o1��Tq�ȅ^J7�q+.Ӫ�����J �.�g��[�#i�;�$j\���L�Qr������D) ^|𤃤杌�ڟ8�*���+[��Le��v�@g�W:�b��e��v���L��}��τ�h�N�9��z-$��6GT����[!�)��mQ:)��(�4���6'��uH��3O�m��o{wa[J�}t�����P�<Lq�St<=q^��]N� 63��������yI�iLk�h7W���t-��A��z�Yz*[����KM�j�p��<�]���0f���Kc�@�*	��� }�MKrx�W1�}��Q\E�7殇�qCLZ�!o����KF�N(�d����D��N3�<!��v�h���[hv�
�>��b������\�>>w9����^�JNƨ�5�����8�b)��V�v;������Gu*��bV�էY�4Q��#��D֣��bRp�Q�2��A�nt���@��RR#�Coʎ�`x��u�̄"��Y���yB;Z� =������&n7γ��s�2��r��2�aG��5��vx�����b�T�{J�5h,!%m[$��>����l�K���� y�|ǐ{���,Łj;�::���׬��k�Q�㗢��k��nX��6��� �R�������N`����@d]x�Lh�V?�	����J����q����;d2��b��O�}���S���ː�ڢ���:{ߴ��
�؆k,(����w�a_d3,5��69Q+�y��/h�U:,UQf
Z�Ls6+o��Q@��w(��:�_�z��	s�U�G�ͻP�p<\��X��EO=_���|T���@.]�C2����
�V2�+�]Q2t���t)Fkb��ϻ�H;%)��⥺S� �5W�vhr��5���~;����,���7�����:�ɱ���Q�
������gƶ�ʤ�ĩ��1��`��
�*�����@���ﳘ��N_�:ʚR"&�2ys��	���Ut"-A����G�(/���U�)�t��}	҂�dM�]��$|-:R��+	ʍ�֯2��d��/ݱ/�/�;��4u�� ���"M=��\��xK=��5@���S+��p?n�{b�+�6=!/[Y��9��r�O
�r)�Dq#�3�T��mYۮ�ROL��O_u��y��5����kt�ŗ�f�������P�2w�kI�����{,=i#s��3v{�"�H*��w���;(�I�\������Y�j�����P6�	2�#�E}��a��]՘�*���G�{�A��[�g�o���!�v
a�"��	;�=�A2�1s�*̇=�(�M)��ķ0NdD�`��׺�*�\Kv��� �Q`�QP.,��[WO�!g�d������I@��ˆ줗��2P|81�('��hYѨ����������cm��>�n��c1�򔞂���/bR�ܟ�֘�@�7���U�����7#TK7::�:��K��&�Q�U�9�^7���@'W�J���gX*\v@�ѧZ)�k�0�_�\��I�34B�AN�㖅��yI�\���F���i�Nd�d��ZgߓX�5[���5�(Xe�#����/����pPܥ�>����/0���%L�Ճ$��4z9�����V�
5s�е�>^S�r���@9�FU];�����߼��Wm4���߃�.5����+t��,̐���.[3��Z��7��[GьE����^��=~���J}!R��kU�9�S�Uk���d0��gU�[�Q#����fU�kD��>�y)�0��`ٌD����,?A���q�9/���׊�,�J�=��L(Ms��z�E����
L��#�Z�P1�6�l�;5�
ˌ��Tgc�7�;��bQr�Eo-����8� ��f�F��5<CzW��7��Qk��������-�\��~�wJG�3WN"��"��]��яkP�	 V�Ci/���e���R.����Uˊ#����$�A�\z
�ɖ���MR�'h�B��6?B�
-mUZ�����𠚞�"��W�X���"IL�	�g.n�S}����^��wJ~�bJ;���z���~�Yp����k��W���ҍ�ԃ���ZP�q�0�S��q�;�?�6X^ƚ��5�/gY�Bա�O���lP������*��kخQ�џ>&ĉ(��U2R���]��}sǭ�ꌇ"�^
,^ 
��߭u�h�hEVtg����ԧ�_���́P�A���:r5���Zάe����>�m��ؾ����f�j�#I�U��TmbI����A�&?�[}8Dl�l��*C�4�Tf�\f�s����.8�#�X��^=�<�����?���?�o���p���42��À�x\�`����y�҅��ˌ��|�� -��������T�b����{�H\�c�Je�A�9��+,t��/W�W�������_l!�z�d�X�����������f��Ϧ�6٪���f�@R��ul�g�#�2��Øq�w���S5�%��O~ltMh�\I�K��z���^zu/�Uȸ�(0|ng�=�NB���ض��{�'$�웉�NHwa	A
뜼k������@^lD���-��G{���:�G݃��������37����c���g-���%\�[�(���r��[N2D��5ج��}��Y�a�7�3>l)�w�����$m��x6jo�I[���K���怋���{"nHkQ�_��oA;WH�����V��6v��1�M��I��bJ�Mcy�|A��G%P
���Ո�ٺ'KN�|��B ~J��JnED��ݫ��>�`��2ɲ��Ͼ��T��
�smR �:��O�����H���e�ڛ��~m0����Z�R/z��U�4�ՑQ�I�<}p�p�����
���D�z���.Z�d�HA��!bo�?�X�J*�sd#������T���L�xۛ%0R9�J�<������Ї�� |@��v���t��rљL��J�+B�/t�FMx�M��L���EΧ/5QKkpL�lh{��_����V~r�"�l�))|8d�@�,�M�(n4wI*u	#K�|z�p����13�$��>ҔC�6����5\��K���1(�=��p�܋����[RGh0�p�W�����.Z���2��F�¿�Q��&W��+��r;�ښM�#��ز�n���)�R�ɷIF���w���Hޢ ���������˯5z�QA�0��3�nV��7Er0���+��YM���.���D�=�X���I��LF`h�5��}L6����n$8}����\#����8��e���= �p�ى")���<�&��M�x���j��@��]$��u8�I��%<~�X� ��Yxgv}|iaE�"Z��ur# �(�e^)6�8��C��{�����`�{�fث}�W��ݼq�g�^�L�z� X�֨j�XZ��A�A��&��Ie�K��A$A�	�ö��O#W�r0LS�`�0��-�ܕ� �h������4G �A�r�RJ���+���y�匇�2yI�;�l=H�+�\�HW�EjP�7S Yk6ϙvU+%�J(EG��8v�Ř9���v��2r��p{���^.��0{b[��g��Uo�1�90`|�r����VeE+�r^寰�[��ȝ[3��ܼ��2�M��J�
$q{��Z���)��c��L����㠛w>��/�ޡ���~�]��᫑�9cN�hϪ�/2�� �=���b>�P�rN�~����?`�c�:4�tiө����I��G�q��b �d����V�R��1�w�++U\��H�q �lg��s�B��	E#"<�{g�Za��'r���6?\B@ө<he��b���M�4�7]V}qΝ�������F;1k����t�h�^#5�5�M�3%P�Ts>�2H~�v7��İ����*��]��f=�>^����N�:��S�'�o
�U��\������%�+��Dh�����b�)o|[28�\ �$���:׭2 �ҝ	�_���Ph��䮧���È���jR�w6o�O�}G�f�a.���l�݃VN�a�r��u��t�}�~��c���?���M�T��0�;hp�4$�X�,�$��_�˵�N�+��5���/��-C�6�դz�I�T)8�?xCŢE�i��k�
�¦^���{��a�N�q��`��][���Y�!�a��^�����"U��A+��4����Ne�#��6�&t��R��$��x�ec�����J��s>��P��(���飐�Ⱥ�Nk�^��
K���,�r�)I�A>�{5*e�+ߡ����vXs�VGi@�_m(�	1b��.W�Ĥ�qk��R��I�	[���9i�'��B��ħ�U�ej[}�󯎋�a�B��LU�q*a3H^
wc�ݴ�?/([����EΦh{S)a(��k'��I��$c�Á�n�(͎�LI-l��� �
���R�Ҷ��P�rr`)�����*���B��䃌o��	y*�2l�ߠ�K� 7�䩡@4i1�/z�7�Fd]�_�{�3y.�0�Ҋ��G��[�A2�8&Z�]n�S���Ex	(
nO_ݚ}��}�=ʇ�\��#� �6aȶ>�#�c�S2/�q5?3�{&�����ʗ>��4lx��x�7����wƔO��h'�6��E{�[���?�6PD�F��#�!c���������I��tr\q#���������5՞^���>g�}}/�V)8P4k:/]� ��dw0��i^(o���vN�C��8e
���W����|���sC�usύjr�	e�]_��
3{�
���z����р��	�%��+�`i��S���u�������3*�ћ0,���G�����?- ,�ID"8�v���*Os�U����O��}��\�=��%�0�v&��^�k4�q�R�6�f>-��8�_f�RY3 �;��^o��T7�:s��H:9��<�3!��"��xL�ӡcY�k��{{l@�BQth��ݡC�y^�Rބ�3U?��P��JXI�(&�f�O�A���P1z8i�!�8��z��(pG�3]i���=������b�%d`]�\˚��bhd�
c��	�ѱ���ơ�Q2�*�s�}�Ԓ�b*K�U�8&�xz���4��=bôG]A�\6y�vWlBEȖ˨'&�^SA��0���+L������fOm�VޣɪS�|��0�h��Lw������V �e,�nzC'�m����ކ���r�Զ��