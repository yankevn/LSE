��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M��	��1چV� -��wk���ŝ1�;B�dḦ��	rt;Cgo���6$f<m��Jb('�`��Sdz$Fd/=[���8Ry��y{^���WmT X!Z���c�����}���1���[�^�VK�v�݌g�-^7�;Jt�B=~�ijT�ADa�sB��V�X�T'��r\M����r���a��xC�ߜ�<�η�L��>�t�M����`�Ea)aa�\%�E�I(�U^���=�XjR�(� �<���3"��QQ0fuH��� �N�s-jh�\�O�nh�:_:�Č_��^�T�)�rz�;�� �=�H��N����^�n�H�~*��T���'�ib��o��&�^`�aPcz�|�dU����lh�#�64�ɘ��˹���)�� ���쁾�*�P�2QY���`��x�
S�eRne�y��>5��l�����`s��{��4:��Q�Y�V�M�dO��J�zR�ww�x�6\QD:���0�5�mo��- S��z�[1�L"Z�E�T>�S���we�R���t#�L�?
#��]��.)ӭ`j��x���U�YlUe�HV��d���uf��e�Ҡ)���0H��Xr��j\k��U���(����%�u���b��A��2�������	bD���j�f�,�F$<�:��twԡ%���Dď� G���+�0;����i�k�ߎ�`��.Y����~X|�|��Q�~#�%�9%��/�چ�쫐7zs�s��EC����p�q���WqXw�P���0�����[��M=���8p�ä�ۅe�B8s��5�j(N�+0���SE�^y^=����� h�pQdA��Z��0K/QP����An�zh���i��=uJ�h�A������^�.,ĩ��ȝ����s<tQ��������$��|��=/s���>&�@�*�`G�Y[<��J�A���+>jQ�Ij��Q�o-e�X�h���	��lxM�Mتdd��
�l� �ǃ���pb�E���ߎr~�&�m���P��:�j�6��$��0ϙ 
b�Z%~)Y���M�}�� j{�8�-�$����Lu��8W3��ehq���͕z��c�u|_;�J@�?,��C�bX�(N�Pe����i53nÈ�8	����-ϊp!�X��ҹ���i�iT����]ppV���:{��,^Ǣ�Y��ǚ��׆�x.�q X~Q�j�����I^���(�w)K�e���ތ��#�����M�*����ۥ�Wdj���,N�G��+r�yᓂ�A����e|\Al_�<K;�+��``A�^*�(SЦ�k��E��]�� R��*��ste����?k��j&�5�����z,^�q`�[Qe��8EY f��y@D��?R���ߛ@�"�����|4G(Thf��F�J"sS�0�<
��0�Q��5���w�{����m*m�?�r�w@���}Z�)����˭��g��mhhk �T�O���I�m���|�8!��X|"�H��N�O0����� ��P����6�2`�e�rԘN�⪵�fY@`�\��D����-�Rx5���)�]���D�ᖺ �t`�9�c�pq�0󼄏X��(n-{�/DK6���98�xHV��!�^�3�X�JP�ߝm�4�(:!�'SK� %};��|��R�u��দH,�b���?�:���4A�=C�7Ԩw4e�J�ڝ�4J���'R���ZJ��?Nâ\�R�;K]��8�g�M��hw�#A~Ģ����g�3À��2~���Y����3q�Dʵ�G7��2	�#{�^��Je �&'��zp�c�f��g�q�ۙ	P���UL�u!�ϼ��Ƅm�	�1��K�S���;�3�{+��^��<�Ѓ^N�.�*M�����$pL������0fڮa���M*_�exM�b���~�� F�H�e�Լ2!��X���\IR���z�SK4I�X��\��㪗���c;e`J�%��ϗZ
xJ�����Eٴ�����[I<QY�N]B�M{�?����Fj_��ȟ��ﶊWS�M��x�>s��Y��0���Zs���l*�Xv� }���Wt��VN��x܂�Q0�"n�9iO���W�n3� �w��8����3