��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*��=z<��t=r��,�3u�:�S�$,���z�U��U@��z�2Mn�������1��Կ)�y����>�͓�$Rb�T�ݩ>,0�J��|\'�������}�fM7�*{]f�/)1�(�S �:Q���4�vS��S���/"��s&�F�;��0���a�M��q���I�M�2~�I����C��	t�AgZbDtcfMg㨎(M���#/(���`��������RF-�+CO'���S�Ө��ߓdM�ٖ,/"�˅�ȏ*����)��+a����k�e\�/�4���ݛ����V7�!ī#�2uC6ͤ�!�H�++�Pxk&��,�1�᱁.�?W��,7�1�4�	`+�i����bv;JGс`F�͏-��,ڔ��\Yx��\�&�����s�(ѭGz��K�4�����kȲ�W�� ƣ���Z�v�����i�	E����P� ��с���°ن�F�G}ԏ���s�/�b$��EwR�f�eC	
�yuأ�`��P7���,C�u�Z�ԭ��mѷ9a�M�Cg�Z#ֆJtHw�L�C�;��p���bƄzy�D@������KDY��䚡�hu7�W0QA�����_���D�8�ݎT���%�@H���P��)�/�\.Ă����d�S����GC�뼢/ڗĮT�L�c�����P}\��8���*x���'��-��Q��7/���������~�7x��zKk��M�H��?�C{���&B�M~�W���"�N0wì��J��c���ݰ��H�W��V�O�?S��ep�=��p��q5��c��=�So��4��j�Q�ο���õ@.�%G���>��Oh��3Q�3މk���k}��w�S���ץ\�3<�b�E{����4�%s|�X�RP9��\��I��~�)��iȱb���X�B��JH�2B���p�ON4Ff���� [V�Z�^�:��@T�'�g�.0ٰB}�pJ��:j	r�9��}�S�ȳ�!���DXpq"����=������R$����-f�/'M�ZjC	�GǠ��3sU΁����'.e?���!y�\����N>".�������US���b�႖��[�0L!�ֶ��nN��g�*\1�^���B�t�s����k <����^�1s(�f�ۂPհ��Fy%�3`f|.�]q�gnޝ��/dF_��0")^�˯b�8����G��teWO���9�h���F�������W����O����-l�9�s�Y$�!ya8�F!rZ�W5�i�A��.���bA�ͤ
�w�/Fyͅ��$�`����]-"�JlI����I��oo�Y�)� �.d�!�6$��_��;g��i;�)��X"�C_O �T��:J��a�8L��X�N#��Ț
����o�wБ���%�s4oۜJ#�f=A,)<�>\������O�sI���=#��`�)��������`�DᏍC�|-;��`}j���7"W��G�f�e�/hd����� �b����lg-wM�D�����F��Б�������n*(k�.C7�!�E�R�B�\W�"(�U!ؐ1�݌L��澟�Рҍ<JH��`��j���$��x�`��:Dpv�έ�ɸ`�C��g���3�.;���E��n�4���_�1g���ٴܐdK�w���k��C�)�/+�8.'+A�|�1i9�K�cS�AMܴCGa�x:�ߧR��6iG�k�_9���_���|c�044]ʺ[V,y}'��4�t|�HDdFF���^_�N���C��##�(�kT�`z��[e�p��!N�r��w��?��b��`��2�Z�R֏��U��ڍ�GeћM2"��1X5L������-? �$�Ièy<T�[Zj8�����cC���0��
��I��	����/Wُ ߍ�{�#e,��p��|���"�o�9Q�6��2�l+�2=s�1q�?Y�����7.�M��
 �r���Q�����B[h�i¡�n�8D��@�� <dNܴ��v���yb%4���Т����A�9��f�.���9M�-�Fx�����L���&2��� (G�7�g����E|��K?.A5[ݱ�{[E�F��c��
7�������UT����ǋ��b�4Ś��	pp� W޻&Lj��8���v��
�'��7�s�]�	��r�2��jĠnl�w~�<nݽ �(�bI����BǴwGT#���z��aw��|$�@a��eq!k��V]e���C��SWΞ:�;˴<��.腛�4g#��ej��V�42J*]u�E�Ֆf���uنz�2q�Y��#��xv�K_'�g�˯��Q�,�|�1�O��$�Ʉ�Ǘ`~�T�4����y���E0,Oē�*�2��W���Ⱦ�W� ��,��t��~"�i����Y�������S��MM��4��uo3���奙P��u��-]�6U����w}h�֩JgO��������J(8�|(�گ���Qi;h8o��������k$�|�G�/c2V?����i[�1���(M�7��l���4��ɯ��l��W������]U���	y!���ďqŖ��{+)�Q������wa�#��1(b��pBcY�u���zN���p~�8�#ؚkO��b:�0X����z�T��^��/H��*I���-V2ۀ=R�����O�1d��ּ`A�4�Gj͇�X
�Ū�m���k a�n(���GbiO����R�Q��s������e��6���ʫ���qKC[�<5���	�Q�+���(��̱Ox>c��/,���y_+YWTH7�2�j{���]}év�g���~/zμ�GQ�Qң�֝��ހS�{����n��'���4
B�v������S�5�L.Q�pXYP��+��l���΃R�gu��)��Z7��X1�*h-�_��U��[q��R;9�G]��iK"��b>3}l�d�Z����W����-)�v��B5�}����
��3�.{����x��y
�O7�Ц�Y��o?�X��3�~{z�))������Rӵ����s��[,M���n̑�rg��D#����wg�:2|��q�b!D�YV���m������t����ʘ���#m�)���<�'/���?~�2rx����U�ʛ���xT �e���!�1R��߈s���-3]�̨�ry�r���C�)8ͻ&��Q�W���.�oh4��f�=
�Z��H}�!�ᕄ`���R�K�{�<%�3��O|ouk�Xhl���4��%��TH�V�M[X;����"��0�������mph�'S �~VY��;�_ܚ;��'a�sgl��Z	������W�?�Z�h�>�߻73�Ż��9"�o�;��h�	��cN*ڽe���!�lf�f�.=�.�{�9�������ڿďJzz��1�&m"@�Xo������*�*䈐�u��vhC�9��S�:��BXXf�W�D ����.��9��'��˃7nh͵}�m�[�:����kW�L�ɣ	
!i\�O��p�=~S�*�֯!І��5�gE��S���	�>U��M��9OM_ ����,�Ky��� Dyy�3=�����/��/��$=vT8�p�|	e��Y��4GQ4|�;}��Y:w�ff^����oM�35�p�a�d4�?�[���ol_�~�\�)~n�������d:3�o���T�2�ŝ�%�[O�z�}�<Y�����	��e|����^P��*���a�$��V�~B�c��ӵ�/�8n��y��fb_)�'|���e4��Z� ��
چW�w�X�-Q�$�"�.XJ��g�l��\����W	�Ĩ}���PÔ�y0���f
>��L�x�K+o���5<p�J�E�xŶ�m��L��~����j6�0�,O�ӹu5�Nv^������5n��m ��Y��?x�-�d�&���g�a�0YYG"#Ua��OA�N�3�	Kkq����.��؍'��~�&뵵�b���1e���1!�ܯ|)������)�����?ZD��C"� ���"�ly������ ��m\I�+ZF9t���TF1m���� >��1\�gQ��ל����;=p%��N�`@��I�c��Z��n��X��r�[ËL��� Q2.���OU;@�Qr���;�X렉�ٜ����w��DA��ٜB")?���NtQ�T� ��Y3�]ec��,��Y0�j&'��r���EeR�G�X8&S�I�D0�}M+&�G���V�s!���9�:[��ohp�t� �/!�-���m���D�ww/W�w���t�d��4��k�]V��E�Q�|#�c�q��Ar�k;KK�h�ݔ�������_���߂��PJz!K�_ՠ����Ĵ��1��$H(�<���g�m[�|�#*�<�~B�b�Z�w������]��)���S��ܵ�i�qk�Y}%��#Xt�s0 �V�P�!"�s�^f����d��
���l��3��麔�����h���)dI�P���y��q2�sO����ȿ- h��[!������Xe�J�ґ���d�;�R�� '�g�E#�eZ�z@�#*������6�<�1�4P�.���_�������-�}��]c4�{5�wu���&{�ʺ�f�{8 Z}��+4�a%��/��t��]��|
�����G)wq�v^�S���~_A�k�KAc������^�L�ed�ă���E��rKO-�b(#7y�nu������[�6uEç���'�z��̜%]��|�l� w"e�E���ӫ�yQ]J��nD�俉%,����a_%>e[(o'M::�f��)J،�k|�Ï�I�Vl1J�+^��j�	S��^mjb��;�~g�i��i��(C���S���twa:�s�e��
�Lpl��Sh�S���Zk���\�p�> 45���¯��IY��J�h�P#4XϠ-������	���k�Զb���y�kJi{�"8 ��1�������ghl:�T�N`p�~F=nRWT�FP�6c,�I3���	�g�  ]����ۥ�qF)+$����+���CI���bXۼ���_�e뒠�Ͱ�1��A��E-����<AbƂ(�Zc:8%���c3�A�T/�\�����f7H����|�$������G�3��� �c�P��F
���m1Gٗ-1m��@�9��ǝ	d���3���n@��e�0Ma'{Xl���j���r ���C��}�7(�4}>6ȗ��kʩ��m!�	/���?]z��o�>���	ܒ0�・� Z�c��ʆ��ͫ"�w���ʗ(��f�����&�ի��舶!�`��5��rV����P�N.��J����z��s�WY� e�^[��&]��yG_K��O"�n(&~ȣ�	D�O� �[��.Q��'[ �����mи|�r������9�Zw�Z��ᆿ/�"�V�O�9���f\�)�q[���6hhm��hHb��-�b�g�� ����3����[ݴS�$L���V)��6'��=ֳ��IS�̆��R���Z	�1����Շ�����Y&�msh����M_��F�QC�sAd��ƀ�����*��j.yɛ��[�/�"�5Mc��Kᗥ���'�����|ab�MŹ�;�(�t]���@���HwW`
�n�����4�;��(d�&ɋs�|�E�h�X��>��FVh��
?�)���*���[�p��i&���6eؽ�׊���=�p�/�mAn�qx��@}���U���r�����)!��=�+�6Ec+ƿ0���*7������K%o�ٙ� ��&M��l	�wƪ^}7���h��I!��2w^'LӽH�p�	�8�y�i
���ϓ�e��D�W^G�n!��b�񷷂�o��Θ����_|/(���A\`0-�� �S�'o1?u�� �&�hk:�0hQ���d�t0r��k��1�:+�~FPH�q� �D����|)сS�=b�w�-P��WN�fY��6���]Ds�\�Ut�
h����^ ���7q�[[��mxZg�Bm�J�@��n��A��3���[�iv�5%���ئ9��T�%�o��&��F�
5%�PH=���4�
3ET�j�*f�``�v`X0	�TU�]7��h%�W���PB�L�d��OF�ߓ'	��h����m퓄u>��>��Ƈ�0�oK�m�?s���}g��EL�'��s� �t���@Bװ㕸9��`��)U���=
���&H�{Ca0�i�x�bH���=���߈K��!��W��a�N���x#�Sm�m�ߘ������h9V���2_F@�2%���!́�����A�Т�Ĩ��谿:���d�O��{⽭������)�ڡ�5��ѼЋm�)�߾��2Փ͐?�!47l�`n7G��G}X�uϨ{�Y��Gg(������R��$
��"1>�6�"������`fH$A�j�}Х���_�h3�l�������8��}�;5�]r����k��@��gT��x����Uj�=/�6,��_(���{&7y�[`ۇ'� �-q_OSɓ���Jr�v�ՆX�Qlaj��O XA9��_6Cvڇp�ȼ�)�|c��X�C�P�+d�a���M��pM�P~ �֖����BۃF\<%�/>Bm3eu��5��5���� ��+���'��(�A� �	H�k�w������5c��ۑWZ�p��N8�d��Wt�}x���\筸7��0	�hܬ4�.%��KkY��;��M���6���#rC�e@~�fFl��o6ڻ<I\^�k�c���(|�3���&�/rFst�4G�<UD�;��"�>�'@�i����l�O���Z.׀5<@�[e2�������;a��WWo~�V�	S ��TP����t�x��Z�ās�i?�+��[���W�$���k��U���N�"��)�7��߸L�< �p�D�R	Fg������P�_��Y��#*Ms�?�g�+/O���~����/��c��I��9��i���u*������G��򑗚jC��'��	\e�{0���Q��sk���U���d���ݨ�r�����%�cކ%�:�&/t���s�����dp���:[ee�M Wgl3��aZ�W8��2�[Bk��[�O�^R^zq�s�_��
v��O0Y�2Ȣ�'�ݑ����s��yw��C��i��"��q��X60-9���`�q��_���fTf��J�$�t���߮_\�z��anV5�Bb��e�zJl	_���5/U)��X�5QPb¶�|��j 8ţ�Hc2%��LR�|p�}� $���|'����{�Ո��WB���lt8Un�*�u���M�X���������TP� zQ�8�[��cp���o!���H'�D���?RXT��!�W.Bl�����w��#���@�;��O�gj���� �f��ք��J�P_�g?M\_��ؓ�F��~�����[���+9���]T�1��4���;w�Y���E���7�FP��0]�f����J�t6Ui����θoU�G�=*4������������`&��E����@WAx���Gy�� �J�����w����������p�-Nk�o^�s�yh����6*�ܸ����q�<�X���3ݫ�SmǤ��)��N\S��(��flʾ�ʐzv�yh��r���Bk3;?����Z���Xw%�U�)�N��Qk�R���_��F�J�"n?��fb�C��PbtM/M���&�2���DXM4����ÒI%ޓǠ] 9�/5m�Ts9<y>��ųb��+�ƫ������m�qc�4R�0��CM6G���Rr��� �.?2;CA6%�q�%pi�s��Q"�K:�s�� (Լ7�<+|�9/���Q���,@�F1o'װ?q��-H4�M`������q���t�[x�t�YkOY�%i��}BF�'u��*\���Y���Ҧ���Ynt��Y;,�q͊����X� �m�v!Hu*����}�Ič�x���gr^��j�yW"�_��%����F��]���h����(ߥ�^���Q��;�BEF��/��6�Q#���N�e��G���ߐ�ԈR|[����4Y��CD`���HV��Gz��'�E� ��8���Y�/�:"������c��cZ��Ά�����şV8���)O}3��rJ�D2n�����B�	`��j߮C�Z��S��b^�{���^�W��9?4��r���Yi�X��c���5`T��i�����|��/��+	X���iE�kwuV5p/����/���s�����l>o��;BN_dR����U�̎�S�T�G��Gkc5f]N�e���2^B�8#�-l}r�:��;��r��ܨ���8���-��&��|�B�9d	�[G��)
��f��l�!��g� �"�G�>��� �3~p�l��!�-IRnH�K��� zM����>�Բ�<-��x��7����G����x�ɰ�ɫcQ��Y8G���}K~|�F��b�$�ebu��LN{�5Gpߙ2�����=Y9�Ͳׁ��kφK�w���]�5ׇ����n�D�i���� i9C���Jt,=�n����b�/����8+g��"T�РS�!Y�)"x�����SAe�/�U�D=|��7TLE8Py��C���PU]�Y�R�k0��2R]�{�rO��r�~�%f:h4�\g��1�����_���̂����y$<ɢ"ܽ��ʻ�ٹз�ͱQ����%(�D��'(��=3�e�ҿȞ�ͪ��]n��������F�"��,3�Tr�/Ȧ�Нe����v����琢=�a�b,U����r;?�0�
��I�)J>
5�Xcg������)�%[��]t/h����
�9QAt9�Ìr�O"�/��х洊<��p(����<���F��B���Vn��/�a�GD[>���ї�1._;?�6�l��k��}	σ��}"�Mb	�3I+C�s7�����:�>�+�v����i�Q������1����h��"	�'�:�p)�����f��!a3�)"���Hڻ7}�{a4M���v6ʟ0��b��-绗�]!�V�4��P5����%���*�� �|�dk���gk�h�$������CN��P$� E�tIM.�? 7b�����Z��?�>켼}yh:T��ے):L�`�:"i�cU�0��5[����Zd�����E��Nkwh��&06�I�P��ѳ{���Z�p���j�����f�@�&��}��aUӥ����[�V�?C�*z��L�#[8tG	���[ �~��C:��)�ۜ�!w������ 2��e|NL k�R��K��Wm��
�������<#��1�->D�VPö�o��5$ђ�\�E��8c{(���@QU����A.2PҰ��Ve�̯�jp���p;�$\N�3M�h`�8�'^w�5Z�lMg<� B[�5�ɡ�^cNz#+������R�T#��2緞N�t��Y h��bӐ��-�6�~|B�x��H�QG�>9"���`cUW�p����$z�aG.��k��� x_Cџ�/K�q��0ZѬ �)�f[W+�TU���Fp�3�^!-}�m��Ă�O�]m��)m�y���N�����S�#Ӫ¨��M��������V���e���@h����e�X���Sd�m�\��� �K��$���.G���*�	�5�`�av S���8)�P�0dS� ��=j_�th|%����RƩ���yi��Џ��[�����!&uvۺY�D2��z���s��I�W�ӝ�Q��M�d('�kD��yɗ��9�R�i'���a`�	S�Y,P~p&[sx�"0u����C��W*x��e�tϿo{�V$�I�M�[�+M��X��ޯ-�Љ�d�6�@��t��^��NhY��߿�P5��+T�g^�xG��:�0eA�O�� ~w_��4$�w.�K��zQ��H���\�I?	!������+S�}��gٝ#m!K�?��࡮���z���w^&*�Zj+�D9j{��l�M�9�r=�.���Bǚ��Q��C�JK���!���u�)�Pk<�InƲ�;R^�ȍR��������AjN�@E�P�џ/�=E��4��.�уn�{�@3V�3|	����U::-U��ٶ#�@U	y;Q��w	+�!H�-��%�L���LroW�,���׼��t\B2R���1�7��*� ��2��9���jNvn5\\�}ދ���9Ad��G�f�=S�$JX�;�����e긠��T`��f����%f\/�B�bi�	a���yc�QՌ�l�!1�du���d�i�P�L���
_�ba`���)��5xsŷ:J����Uư�N�I~����ꡭ� ��GF��{b"��;YSZ����&�l`4�tH�"Up�t��m0��l? �lw��F�Od�����n&0� 
΅��몛��検��ϰ\M��zܾo��T���4n��P&�����q���)Ɋ�F�=.K�׻�ihs��T��^�,z��m�rtؚ�V�
�˹�:tnf���PG�����W��T��E����Vv�8�s6uۤ�(}$N��[���R�"�� �a(Dx�[��:��X�l[s	g�hq�]�%M��%���s����D29�L�v:�C&mk?^*3�T�L���
�b�\����n��O���c����/Q��s�
rHb�W���hO����n���e��V�k�e�����>miv�6�YZ˓��1Q� �
N�9'�*B�(^����x�A.�)>� N:W��QD��_!+!?I11� \����hg���R4z�V'��W:J��5��ߩ�:F��T�`f�G��~gy�Ð��C, z�y8�I'� q"���ׇ�Q�JFjZ]�>m�� ��������p�ә�ߠcp y�����$Z̜�+�=Btkd,������>�4j� ��3���n7uV&W4���-�/�*Q"��++!��/��+=uz�[m ����Ö>֭�M�Զ��|Hn��ū������'D9�+�D>�W��R\�&��0���M�~%�.<��r8����<4G��WV���6b�����t���-�߼������D�݉[{
I	-
VC�2���1$��(+ 8=L�3��ۈ�����B��D쇣 'I�Pf�z�E�)|�I���82����ߘ� D�6��.(J��7���)��mǐ�|��ƒ5�t�����cN� ��4�q{�}�"�?��&��'!P����p��l �3�g��t�	�R�b��R+��A�:2(��İ)�iO��Zt�2|"1V�B�[,�%?��%-fgǵ ����̔�-�Vy�s6BRQ��ۛ�`��'� ��F��A�������)8�u"a\nI`�9QM���Č)��58��e�ѝ7ˊR��l6~���k�t��E2溦L&![�]�]���=HnI��9.�c�F�
��{��?�����~��>�/��Jg�h��W�ϸϼ_�� 81]�}9/�����g���*r��h����UAg<8(�4�����Ы��H_�W��D�����������"��d����b��9Vct�,	�)����6L݁���9{��L)�*�3n�L��e�c�F�Z�y}�����0�1y0�f�"�; ������ar��>�,oӥq�G54r�'tD-����6�'� y�Z��_��ރ�8�I�s��~�	#���!vǛ�Ɗ���/:��1.k�d���x,\�`��86�WO�'V
ҋ9�h8�A|ˊ
�+�K��1ŀ��~��������7�^��ҋ���*cϗ�b��Ԓ�Y����C9�x鞊}�Ћ�{�P
@�m��m�J|���߻Q��7Њ-��Z��3��q_U_�(��!�H����q����xޫƶmﰤɀFynr%�+�v�[ �E.��2
����M��=5e��K�Q�1LV䱷��$BB��>�k-�(Ę�.���$ľiώ7Ѥ��"lk��,�z&�L���B����̀��pU��[�n;����̠귍��m=v��qGi���}<�-a�����H��X���h��c57.�Gw\)�v��Yb��|���f�p��V�i�xʗ���O�a�+_�J�_�B3I R\��5xM�y�Qh���o�0�zL�S1�J��k�	�=�3�
���	�����ڤ�ج�,�U���I��se�
~E%P>!����X��aD�dD�e���x�79eǓ��6O)��h������cA�_O�x��(7�����߷M�T6@5��h8�V�?�_xZf읺^o�r�q-�,�dD������ҺN� �ĴQ-��s������}Y�1��L�:Bb�7�"�y�k\T�@}�Ln�'�]2 ��pYoP ��x*�����Y��׷��G�����r}�Q	~�K	�:�Ţ>�q�>�{ݠ!G�1E��-o~�&|���ik䎏�.�̝YZ�jՠ���s��3��#�����Y^��%�a4�W5�0�-2��>�3E��;Ëk����8�
�fA�T�.�׼\������UP��]<⺦����J&2���놹d�Řl�d>얄{�xgE�"
D�2�h����	8�,H &厥���ť0����܁CP�
�o �0������0;��H�`,M�C�~�/u�W��s�\�pYN;\�� ��x6�h�j����r�No�{��h�Ŝe_1)ʻ=)��y��3B�ZaTbX%9l�;O����4:p�F��ڣ�#�K�jGԩ�]U��@q����΍o<��	O���_G��$���&=;� �,O)�/S��U�wg��1�͈Y�4�({T��������Տ� 46Nu�@b*6��#m�1ӆ���d�]���LqӪ��k��A|�����6�å���?]xj�%�-`�&��
��3,���x��MI;�#S/1���[֝�tK�D�T:�a�a�lc�`V�]�0K�c@����C��3nLeZ�'V��;��b��-m~;���_�q\�B�G�|�B��ςl% ]��EPm��qX&�B�t0#�@l�����*u���] ĺ��G%Irp���	�DKQ"Io���dg$��N1eli�
�#KW��n�-�������l��ǅL�W�9L�T�JB$�$�EXn!���(��®�F�PL������G�\��cf��d�ً]?쀀.n=�aF��FQ�}�L(�Ύ�h�thj��e��͹�}� �G��s�i_j!a�j��y|��Is�E��V���^����kH;p2%X�N���TA-�
��r����b��18��iSd��z:UKMXM�����.�#����aWp�5ra?�j�]f�8�u)M?#{����%��j">���c�߶}���v�kuP+cp5��ٔ�EBD�I�Z?�)c6�5%�n
��$F!4�n��TEW?��L\F�_����wֆ)�<D�,��xb1\�O�2�duv�7�6�Kn}��� L����°���螑T'bo��0�Z��EکDO�ň��	�x� 1r6>u󙓠8��9��*�ɟ�u/��d"�����u5Nt\k?)�l�'��L�WK�V�O[�}_��L3aU{1I�( �8�x��g��Q����R�J�����mΖG�7sJ�������:a��(����o�ʷ����\B�GR���OݛOv�j�c��F��A��-�wU�:�qR2C���I�f�k �V?�#9����� ������s�
�y���9G���'J*Wq���/��A��=�e�W�.D���j��X��ȧ	�L��9*7V�c5=_���^
J� %ΚH��)N=hd$��5*�-���l�`?�.!k�r��A<*�L���b�Sn#�b�̡�e� 8�����!����5��	%�}OC[�u�����(�u��x�䈦k���`��mo|*�O�}��E��ס[�w\��M�1��0�3C���kC���<&X�`� �@��p�C39�k�BO"��OE�+2[CGQ�U55牘�����r��.� �$Գ.k���~�H��l;	i1;+��}GפZ�ܗL��=�f^Vd�,���>#g,м��Qi19��R�b=�@,��˫]���3��C���Ns�w����I��VE�ΐF�}���ui������xD�)�6�VQ�������e.�V��=��G�|ʂ��]w�ׇ�޻2�U����k���ǯ�n��iO(c���]�����o:�(Rb������R�Y��H��tu���:a����2�F+��^dI��
 "�9>���@7�� 0�Yۣ 7/98�"��t4oOV�Q,Z����)�:q0�����8�����e��s���}"1�/�o.��]��?��)B���F�!�X�[�q z*��8��cyk )�{4ۈ�����r���Ы�M�^��e�l�I�dL��<B�c.�*��}�@к�:���g��kO�݇�9!jH�f	�Rޞx�q����TG���d<'8��n�������Z�f�wt����]��Zm��� ����e�NB��˝&��G?���v� ���Ep�.~'���K�`�I%@V�M����4,7jx��r��T��׻�O�w;��*ŕ��z:�N������( . �-�m_�&0�MU&�K�D�O�6��w9���p��sA��z�]�'��WY������.}���Q�3NV��|i�p��v�(놤��͘�� oBھ�.!P,�/U�F9��6�{@���)<�_]o�Yҳ����F��(ՉÑHu����y�wU$&���JH��6^�i z���Ҁ�F�i��л�r���1�+B�Y�l�����E����}�cu�\���+�ۑ/U����p������Ӛ8݄	�uÉ�𼆫�����F�}��b4.����O�>^x"gq);N@˨�LT]O@�������f��!�n
�cN�{��t�i��]��U4r*��R'�N�D;HaX�~xYXV�gո�t�������e�r��ܞ��q��c�9QK�l��Qd�9��f,�NA��˳`H[�-��D[�!Y�����1L
P���l�`acDN��СZ;,�R��� 7r8�]Qȸ�~�2ug*Di�e�ր[�.���d�E�)r;�I�q��洙t�g�b�2�៽�r>�Ew�GBX�L�ڪ �~��w8��36D�o@Vt[���������|��eX�_X8Ƽ���@�����@]���G|�L�C"�28_(�!��ӳq���5��+�����9[m��%��b�[0�@���h�'t_=˓ �$�E온�G���2��glesR+�����jShF~�s���`yl9�;ER+[^��u�h�^jR�"���Y>�e�:8���YWb"�\�^�T�(��+1~ŝx �+o*���v�+�Ǔ���+��	8۫���om�T$�� P{�c�����C�N��'�V�4�s$v�YCDpp�h�x��R(�y�<c��N�*�[ �o�iXAf��ܠ�/�9(;��Pg�!bdj�J�T���v�=�n�M��[^���J�IftkW[�1N���q�Cc�>��0��D-^�3���,��t�\�5 ��������4N0�N;?*��J]�+4�̴��k�DJ#�
��!��,�e@|s'R���>вJ��X�2���0��_]���G�~��"<��5�:M�^�Z��������7ញ$xV������EC��c��b�S|!v#�L�/���&����z",�||j!u� ���c���+������#V�)oQmD��B�	Uc��ݎ���b�J���'�\s���w���B�$9�dQ�[,]��0H�U� �a����}��R�[���AqU���LU���hdr,�44�s�4X#��&�9b�T����b=.��4�r߅\��Y0Ԁo1qx.'����k���{�
mJE�B����G*1.�Ycp�[�Y�PH`���]z�V��(|�m/�?��\�.����٣]*C��Z�si,���w[��gR���;W�oe�[�M�<��@���Q[:i�)��m�l�� ~�����TKGҝҎ�uּ ��Wq�W�_�D�����}&tB�gC����אꬿw�&��u���x����"C��o���7c��U�f����� ����$s]j�`!T��2C*27PZtѝ(G���s�-Kp��4&����~]tf��j*I"�8j￫�pm�\�$KUu}UYԢ*�@1�\��R��<u-�5ӬA�����y�.-tA��!`_|����0B8��H���� �@x3�����m�J����/��#(:�n(��PNO�xM��|r�&���"�C���p$���r>�����#f��㉓��}K�Wv����qg���C��j5F��
�C��Tx���A��>���Ⰰw���w���\�7�(�<����BD��ta���}v�����G�����~�ꁘA&��3�O��\y�m6��Z�D���3��O�p��ټZ��n��,V�}��Ǽc%5�:���+��n��+,3��U��D��ăYZ�߇;�r��� ��[3S�5	j޷�B��=QU������rA�Y��|�j*61����6x�]�B�<��q7�sJH%J*^x-�1R9��WQ,1:eK�z�	G�1�BthC���d�ڠmHH���a%�)���?����o�԰�ُ�_)��$�'�ߑ,��V��'y[�Q�uLU��Bm嗶�\QnB~�d������Rk�խ5|��#!�j�Z><Pw:�Hw�l���iW�6/H��QF�9L]1� ����L~�ѐ��~��/���@^X��!�`��͒N��W}�va?�-e:�L!�\�~�m�.vѻ�we�Za+�))�	ޮ�	��Ba-^a��$N��#�[_���	kn��&���~1qO�>�va�S7�c^s�2��R&�F?� LDt7��9���Et܃�o�Щ?�nd9����h. ���	�J�C^s���Wֈ^@h ������oї����}�r��M�K;�Bƞ����LhЧ=��D�U��A̤��I�%՗7�B!q (�Ù�8��/¹�'v�"W]rc2�6��*����ay�W7��/��t�y7��������]��ۆY��4<����^���+�];�WTކ9��:N!�6g����L�]ٕ�h>r�uD�/�l���-�U�n��i���)�K��A#����Ӂ��V�#_]���%M��������~>�P�� ��-����}v�b�r�]�M�G��_Lݞ����D|Yz�[�����j��_*6���fa���P_ 'ӸZ�[Wh�'��*�4�K7�Ub�v@����kw���S��.�	�$:�
���xDzb\��h��^.�L;�@��yi��`�l -"r��ES�Ah�xg[�!e�%�i/�;�}�)8�>Mǉ��	�5J�j˖����W�10��#`�CI��ʢzl�%PcS��	O������5�C������������Q6��4������R��|��ڮ[�|�?�[��qX�-�v��I!�fԤ�B�~9�ٱ1G�?
3*�9�F�X�������]�������Kz8F��3w�	c(�A������k"H�Yӏ$�H�lw�U]��#Ԑ�6f��L�/�B%(Ȫ��l�YS�_�!��^÷�pC4[J�@QCA��3c��k�T�Z�[M��pR7
�ff�!!"�
����WC�J�p�x0lq��J���>��5.	�S1	�m��o�p��n�G@($׉�Jc1�ZR����羛�"������Q�'��!K/I�c��L197��a���4���R)�����=�@��N��w�U ��8� K���l�֙}��675h��8W��&�֖�b�;�;��I,����7/!���h�VJ�{�i��1�/��ևs���΍��<����$N>�ps�5�p�Ϣ��ܿCX�}���f���
 �����{.�(�%lȸ���u��՗4�dP��q�7�Mf�<GӚ1���%
�k��p��8�?Q���v5U5���}W�t��s�L��H�.�5@ yM�'5�޳,��5_yQ�d˹�E�v{/"�UM���ـ����  ��,�гv���ڟ��+��S
G�Z�A2]9�7h�������S��>w�Ւo}����*�e_���M��KfÔ�/|��p���ii�������Z@x~�A�&ǃZ��D�P�_���@Ć'Z8�nntf�mΦ-&�ϡ��I$��n5��UF����� ��f>ݛ>R�����7�؝Ǥ�Ky���\�*�!P8"A~����)�[vd���'��A�2�T�S�GR�twټ`ũ��RВQ�����{=حk��?���I��O�&�8��"�#b��P퓹��3o���a��,ELT+�#|�����Π�������X�����6��i�c��}j_��ﮢ�D��P⫕.��$�>��Z�n����j6�"��Є6zޯP;ߗ�9��ג��䳲�}a�B9?�??��iI@@�dT+H<�V�s��q�=�D�� eE 2X���f���ՏR+=�.�	[�Q��BZ5���@$8'�����<O>yr��juuǆR�Mt��)��L#Z��/%0��J��څR�X��Ǽ��AX�����)j�k?�����Qe�F���x�W1�� �-?ZDZ�T҅�4��_�6w��@7�c��ܗ7���Cb��q2&�T߼��0�-~�Lm4��-zm���hF��tĴ�3��b'�Ψ���n�*��Ml|�6�@��I�\��>2��J��`��+�8=:�N�;\s�}��Yb�"g�묕Í�mv/� �A�OG62�狌N���y���'��_��7���\��hV<������r��Y���{��w�Px]JO�|�"�#ՂOi���r��w4�������K���?N�*��D%_p �xF��@��W��x�*մ�1��7dl��ǚsW:�Ԥ~ņO�9�ў�alHy#]��y���������U�H�1U�m~u+�E��Fؿ�$T��7��G�q��!v�h9�2���N����G���(lr�]�̆q��]�2*��QI�Ka}��c l�߰���S��[Pj4��Dnӈ�D�9x���XYg>���
O��I�*��s-=�	���7UR��9�jv�ƑnJ㏹�Bʎ^���7V�������s<�rv*G3�)�h�)��֙�~���X}�~�܊�צ :!�P���`�VW�#I�|�Oܐ���$��l�.oH��@�	��~攎v�Wy��c�}"1��ʇ�E��$! ID�-��̼8o"�0��7�F��0��Jw6u{7��z�}���$6d+>c�@a�¨�\n�d�.AՒS�}�R޼ C�f�.����v���ev���1<)���7����$��ր=|Wx#Y��}�W���AJ]�iK#���l�� @�I `���u�<��^����u�̗A��@��	��\��Yr��Pa��k��I�;�oߢ_�Q}!����,�m��C�Z:��� ?��EFn��*�<4�L�RK�x����}9~��i��4p@��$�^s�c�j'���0?���>�>���s��>�����y3��î���(�������I�m���T��s�.L�3�s{,:2�C�*&&�a(�����H�L7��%�q�Viv�_��d�ؘ�x��%ɥtB��s*�z��5��'7 ����\zǦͳ׏���Ӵ����IN� y禳���%'V7ԧ�iH�y��,�
ُ�ךh��)To�2�nk@@���d��͎8�������Te�����a��ѵ,4�Jf'zv)A��Yx��_s
'�;*�>+Th0�{��1��0�6y嫟����1ƌ����(#� �MQ����?��8�mG���A1��tF��/tr���>���795��$�I{�7�����Ʋ�Z�g5j:�f���y�.`-�h�$C~��j�$Ky*,�&8��)Um�_�ۂ]*P���.�ꏰEXJV2�ʠ�¨�'�\�&.�g��Y^0_�����mjHs;|16�$���	�ƗŎ��x�	v�n�dRgH���V}^���6��D�T(��*��m>�D��O�4ܭ������f��TKp@�冭��h���#C2�1S�Ǭ@$�����z���~r��j�`�)�p��h}��w�5E���h�\�<+���i������v|��H�K�!1L���yn�>�^8j���"N�
I������k4�����ʢWDU�X�R�Qj8���s-3�}����[�l��2ʡ�^�Ѡ�M�5���v��u����el�I6�)cb�L��Z�='@Р�aʒa,�Q5��94{8��{r�&�$\x�Ps]�E���R��򰒾�͋���GRA�5�����������?��"��B3qA�#�^.�s�U�Q.�0H�?_�ƻ�`x�Ţ�g��:}[� t�9�'��{���?5���7���w�zE�\�l�`-m�$��o��H�}�<��'�ҪOֆH�2ߺ�����醬��E��W��!��P�Vç���E�C�C�5R�G�Vn!;��O�4F&����cwPR�i �&"v)�˵�T�u2�81%h�U8?�v��-|�������M$'��:8n�ly&��+�hIu&��J0+�Ro�KD }F�V�{~7f�p���J&�^�T䰎l_��
;�!�E�o|+vV8�_ڎgz4�r{�.s����<g<Lk����w�w2ͤU��mb��l�-�]|�m$ej#kchg04]�#�.	EK|���}�Y���q�'U�����a2�l?��D�9�צ��Ț
��ӏ�k���[K�ǁ�__@��K�d=��/�=�-LD��rs�����Z�W�Q��N�U����U�sl#^:���g��Sh-k��%B��n
H[�w������'�+�}5oȋBjJ�U��a]�
�[�b�Q��#�R2�ܙ�p�5�vG&f��{��vV�z�K���Gl�R����v�Tv�뉌�KzRrc"��+�k��ő+���rҿ�p�?���__"E2��'��a̡&��wb2[l���P�M݃�B`�9�jõ64C����S]<�>�/�逗���{;φ��g5��+"/��(»pa�?_�>a��T��?sK����3p���`!wc�~�����,�3ČW�'y�/0%�A<E�Mf;ځF{SEzF!$����|�����<"��q^/�q�R������+/�s����I�r��l;�����!���Z��� ���;0�w��u-��蒶�M������v��?��1"A�+q<:bvN�`�&Nݡ��2ܭs\��{8 �����~�Z�j4����1�ON� E����x� I�D�uV,ГQ� ƯOA���'� �`�I �0+G�/�����F׎!`�gS����B>�4��=Q)�΀�9 ǟ�א"�t�L��E�3e�N<V��(TvDs��Vˤ�ɴ��O�y��𨜻W���S��\�:���:T�J��y$U�K�Ԩj<@j=O��VT�K�������?L��h�'s($��hz�#�Ew��KJVFA­�7���ҝ�u@b���GӔ���R���ؾ��nYI�2i�~n�y$�څҏLۋ�r�Q��ֲ�� ��%H֝@�Hn{�^K��N�o�A�� ���l/��R�l�׈Ѫ����]��z�Yd�g����m��;��	��ˇ�{}�6�������ٹ)M��x��|{š�?����/���`��Jop�u/%���1�	��wt�,+��U��+��q��\��Y]�˭G��Lw�@;f:3(>R�����'�J��X�8L�}��>JAV!�35�ڻa����v���
V�V-r����(9Xgv �/��9�=�s�&��O�d��h6�����c5i�<�(��Q�@��_�]0�??H#Y�Q�YڴH�	I�h�34�G%|��p�iP$�+�i�