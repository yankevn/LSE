��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&����p��µ-��f,>���{�Q���X���V�E$�%�����%Z��2��<L��f 8}� ���m�E�� ߑ�8�a,�D��FxEu/��/|^[��%�s����J�jJ���e_�i�A-P�YC0��r�wI���uHi����x�X&��t��[��L�W�v�h�RUb�r"��78,r���,��5;n�Sv�VA�! �b
6�|�JS�G5A�7Ӧ�Z*.-��\���#��ê��CM��8���U|L���(Ɔ���8V�����^7��d�Dk�T��L�Pm���v���P�]�I	bf��s?v�'��>�@��0�W([j���έ'�H���"كC}��9N����H'�	ϟe+/i� Z�@�k�V${K����*�����n�7v�:�7����ܒ}�|ʹ��ڙ���Z���t�u�4�h����9��8 �֎�ol_3)���|����܄����p2�ZK�)�u��	>���t����-O�Q]a/S�������\��_<b�гGn�ѻ{��y*-���_���c�vH�}t�Y�\]6��yZ���
q���7����<R%;�H��Noo��&�j`��z{-����_�6.����W�md����G�b��y�\��ˉΈAk[�x�UNa�� �F.��cрM�U*�,//~��J��8���.��jJ���%��y��]�7�+9Q[Yݕ��<ѱ��������\zw��só�@�ě�MĹ����d�}�sB@e+�U��JJ�Jlr��>�I��8Pp~Ƒh2%dֹܽ����7a��|��2% s+���j��{)$��h�;y58��[��6�ITJퟳ1��+�)�QϮ�;BR�a{|x��W��Q��@{BR%B�iU4�߫:��w��U)����M�%5�@���OE�-ǿ�8-��/�=8w&�h����Ѯ�ޖYG��ͨ��%�XBz���r��z��)r��ո9yྫ����R��rŜ��yU	�Tc(i#yۥg4]o�IZXĂ�,	� � �x �.#�Se?[(�P���p�J�yh�Ě��7A]<�H��;�6��;I�t�8��i�w�����C��Y��$�]laQB~~
v��u�=~�)��M=$[�ݦe�h}Hp��zX[I7%tk/�%a��t��@CLz�"Va���G�c�`��l"��u�Y~P(�:�.�J�5���0ې���d�;v�#Wk�/�(�P�e\�J�j����"�2��7��7#��ds�+�f[�/�r��Y�����q�Mv�][~k��]:)Q�r�� �У�H>@�4�3>j���Mp�԰�v�ꊷ�y��M��J�/}i��<�G'���v��#�x��M�nFv]ǜs�FG�;WCr��?�q��W���nm1�f��[�}.�M�w���D̡�4XhF-q��ֻ�,�$�Ŧ��L�%��`{�Bmޣ=;���Ej�2�����SZ��I|��aw>%m�R�hH�@;g�����;ݽ����t��)�{�n).�7��>b^˓�N��`Â��͟/R���?yk"�z�*���t}���� �)2�l���+�<%�$uG�u����&`��c���k�Rً��G���̧Cr��h����g�]�V�mRDI ��e���oJgy����}џ�u���>�閵�!��
0Lk@�&�1<����h���>�l�=��"x��[:��>�FQ��B7d�
���5�*�qMP,:)��Av����E�V�.`�:���X���V�;72�a�iPHs�Jy:
�jˊ���T��1 ��Ս���&�g�I�Xި�21�YU�̊ZMr�°cZ_)T��s���n�`P!��?���E�:�Q_`��0a��Ȁ~���&	����y�G��g������ꇫQ�0g'��!� �K����|.���ۼ�}d�ߜX��s,����R��t��`��iU��7���H�}D���O al���*����ϰ:m�F�+�]��_"p#�<�����U��x׷,���<v��	��h��B��?���Q��	]p�3t�"�l��@Z�9ϫ�x���}|�i�����Q�M�
5X�\y��׹��ϝBj���\��W-�ހO��Y�=Q�D1w{�_ͼW!��q���ꊔMB/[&tO�����_T����mW�>wP��KW�)��K�f'�1���a��:	-�S�	�i�����9Uc!��-1�V�Z�����,�K�Α->�Xhl�
\��xY��=Qo3Z�Y��7��]]Q"�ye��KJ���d��9̊�}���|����Sx2J3�q]
��ݺ}�-@}�>T}}�����J�n}���&��+R�A�R7���d���sm��Ԉ0�0�������S/���b��
�<��GU�o&�V>zK����}��g>����`1K�z�����`^�	Վ�՝0D�[���2d���Hhhh<�@W��@3a] ��P��b�N�F�����[&��Ŀz<��N�a&z��Hɳf67k�C6�]wn^��6[�|ӓ�_�P}H�-^;G�k�lg��N�
f�Lvq8���U�+��Ǆ�a�(^403B���pET�mS86�"M˻Z����` 	IE;�FJ�eRiFj��d���C8���Y��S�	�A�Vx�ﶜ�L*D�����e���Y�����"?,�*L>�bhd��ˎ��C!�L�?~�aFl�ޢ9~[w��d�����27u�[�vGYzэ�SJ��i��*��]�/XdM+fSn��ᾉ�;�m�j�Ù�G�GI��.n!��ko,^Bk|�8Fft���"d|��ÆL"ѳ~��o�3��4gҔ�QW|�C���/�&tܕR�ƍ����Ꟈ�!��^cK��F�$68�����l9~��������[q{�4�?f���j�Q������tq�j��{��=��v
z/~!4dqFx���BKEa�eX�%�b�_��m�m~^���˞�O��K�����dW���5J g�)xal�"�{��38
c�pt�V�����Ze��)�q�ۑ$����?-�#��\��v�5Zs�`c
t���2����N% /�rxbø0�׫@���P�z�udB�i�}Q���Ǵ���3�`�p�i�L6��B`�O�n9�+׬Gy�����#*֍��o�oL �3�mӬ�!2��+�'ֽ��+x�$� ts	Qϩ��%��Qw�&�l�M���qw��"K	3ڣٶ�_�i��$v��J�UX��w�����/Ő�{<|^��}���Ά>�N�^��鉴��؎H��R��dX��7><&���<�@��T�i���E[k���RD
 eRyA�C������?��ٿ�A�2z�0!SȷUb�W�]ʍЪ��p�����3g	�������
�▇;٠�"��%u�����/w͸��Mc�Z "6��0�,�Rz�M�7��u��^����#g�De�*���k�m�C�\B�_ɱ�*���;�.���\��^�����C��*�h�P��X�7�%0̀ͬ��:�eE;`��l�#��*�iC�Sm�9PSK���OAW���b�)hq�sh8��H`r� Y�i���)��h�)�1F�֬��l��s�.�~����-к��GR3B ��=�]��*��IK6I�"]���賈?)rq���s�����O(ӛ��C�Cq��#�h3��]���pf8�J�^i�� 
qeG:�Q��^?Q�����{C�B�4�m6)�IYS�d���e_���D�𥤥U�N�e�C)�Z��A� �W���%J>����9*���%X��������7��h��?�B�U�+O�i�<�P@>�����m��kC_�&TcF�sh�Oz�Yq$��<�pp��q�{ޣ�������D����XEG�?�r�@-��eA���Ұ5�xD�}����u�_#(�w,1���k
S�j�NK���&�O"�� �)%{�	Ư˟!�p�I[��I�ZV�z������A Ix�á����4���@��ʚ���������ŏ'%MT���Bʜa?������Jnd�ǻ������쁤4�/zu ��r��{5#�T֙H1;�i��>��4�N��7Oy���m�?F»E�T�%#I�����<ǋP�$�z2����D�f7�^y�GJ{��u�8�3jk���� k6x����/_F7�`q�O<)��������#l���X�D����v8yy�m��R��ߐ'�0/�_}<���9���V7��c�s��X��+�F��4Қ� ���i6ÿ�\��rG50E�^�ȝ-:l#�b���!/��g�7�e�����W�XjZJ�d�����j��n	 ��%v�o�Ҍ�!̡*�0���s�Q]�aaU��eP��4h�� h�{��)t/�#Ȍ�.r d�/Sy� &s, ~�#���>d=:a2�2K��D�_'v���]YݞCS����:�^f�W�X@�kԜ*m�#ш� �vE<Q���S�C�T�wd]����b�}�F������ Y�'Nu%{�!�JV[$���y]����(��@�=��K�ݛ��0a)��]������}��4M�iF���m�2!F�a�E����YaB�ѲB�N^&y��͕�E���������6��#�,p��^���{WuT:k�b�;�b����p��N%Q�3OA^jR٥���B�+"Ϗ[��a�i�k���嘡�_���a�����U<4���z���L����!=�����g����)����,�MZ겡�a�'�]�߯��l��߮4�'�@���x�>�ׁw�v�$]_�-~��8p��p�\M�Q{�љ�M���<�؆���l��G;����S�S)�O�a���5�iU�`���n^V/��;�qv_�͆�x}�<�%�1h�*S'k����5��ԍ�I�~������T�Uk�.�[޾sQ�8��,<K('�>�>b��L�Ғ�%曚-��np�MC��G�	�WY�T�d��<��PZ3\b] #�c���f��a�%w6栐9�S�B�!��$�5��on�lj�R*X����{�$�:'�)�����}��n��4t��*�VN~|��L��M��=��;�7H��@tL�R��H��B ���+�^����UǶ��3L,:�8��	��u@�V�ar��X(WR+y]�B���j�f|1بl�S��VO��E~����ФI�*�����J�C˸U�y�gBJ�-�H��7��M�p�0���5�[�f>6��ͭ�7h��1���̚�F:�*�8i!I�+��G��d?� t㤔$=H;������](��q�9��͸�(��ulW�m%J�mt[I��^��~8�=��i��pN�c0u@�����b�ع(<��P���|�VS���O� ���AoBG_=����A���n�"�@V��������N�����]��mU�j�r7�?�q�n��&��߶�S�(�KQa�tQp`/et��;l�}K��B�d>M0`I�ۧ�D�!S"�ju�o����NC��ꈷ��c�|��5߄��*I!����֍j�G�X�"S�����U`l;�U��-M���V��j��Z��-�]^�]<���j>�K2N�铈��p�'�":�D��[Bb���l�$�P]Ɵٻz���5yj��hRgG�$�ѭ+wV5�o	x�欲�C:�(�ϑ�BF��4����i�H��r���ë�H�p���Tog+ΉP��9��ִ�yj+n#O���_ЅY��Q����ϳMc��XbZ��@�?�Oq�냔�����5��!k�0�����EG��TuV�B�� _�D��B\U"ZW�n��q���d��ۚ4��d���;��9�o���� @�J�#��'�2:��ٹ:��<�n�e9��Ҟ�gXOg��KrK�:��&��֜<y��6o�o�����d3��S!�m�k�|�&�6�w������(�|H��1�W�v	��)���T�#�	$	��V��A�#�����0GOG�����R(��c�ڱ�.l G�g�,�ՍV��L����N��u��MM}�bm�?vNܱ�U���ms\[:Qd�����䯪T�>MAO����Q�s֞��gp!��C���̣�Om��T���؏����+烚i��)Èxm�f��C��[��+7�d��P�X7JcTt�RY�~�6��p86N���.F]t��I�Ǻ7�żS��r�:�#i���F���\<*r%:Bq���QzEzrF0�Mhb���ӗ��aa���*�[Q��ܒv	>��؄o|���4D��P�τHU��9x�����|!�N�AV!�|���@�a[/pi�:����f�| f{aǃXkd����="�D:*��0�Y�o��X��
��Z���9�]��Cߞ�}<�?��-X��i�^��`r��k� ���߸[��)���9斮����Fg�|\��◠��!%�;�e��u_�*$:�@���Ȱ��yF|��G�/`C��=�b������������w�!��+S��gg�;c*�Q_�mmځ�t�o�a	��F�d��o�U�6t�=g
h�>�OX��-�"��������;��=n������5��]�|ǳ���%�S��4F���(�ԫ�	<ꃤ�]А��n�H�7����O�����Va�3��\2]7qe/��o�Ƣ2}���v�J�0,���@q��ywaZߣr2�\cB< �a��?s`֣3�,���%�qa���;��d�����/�ɸ�*jW��cU5���� ��V�3~�%���3=I�{6�R�:�=~4�-S��6eo�4�ͭڅ�4Oo��%ٯs�Êi�z�s�3��{Ԧ\O{C���<?T>�N��8��v`ܾ'�O]����Y�ťiD�('��N�!��� g2��<�K ��G��TnY�UM8 ��pc(����=U��JߔR�{IZ��nY1�O� WRixUƓr�1F������b���gkgd��U?��٦t�#֎^}.h%�Q���NT��qG�����BF���>����U�/��5�gW�z�)Y�Qr�r�$+�&���_:DbF��Vɘ�`�*��vv���AY�����V�I ���O�j�IIjڻ���PБ=�C�|m�>�r2���I�0O�thz-��;j�
�u�s��x��� ou"e��(���vl���>R\je���C7��^^�Oj)��̰	�{�׳1�>��#g`&�\�B��g0@5�K�]�{#�eY�i`��lc�dR�"ĉ*�&�j�{3&
��#��������07��%���`�!z�D��G��� ��mT^�.�#8#��'��!%��M=bщ]z�z���o��g~�٘)3(Ȉ�x��W���p���dW� Q��X���+Id55�fsS�XF�e�i�M�f�c�q�/���bP�~�!��sl�\�#�<���-|L]Go8`C'�6�E\f��=�@��o�2�4��G%_�U����6�g@�!��ktp!c���6�hnPK��� P|?�S���WW�0F�8���u��J�}�!,�t����S����!��g��?u*���t;��_t%�c.��h��
x"�壿݉q]�B��A[�����M����PZü"߾}�ԯe�"xs��U�.��L�9&1r�������(�2*p�-AZ���k��d��[1�pEE.b�.9e`GG ٭�ݐi��X�ᄿ��m��������ΐ���di�����eZ�#*����ٕ2�CF2L�6}Ү���?�����������F��1�nA�1�t��'5�Z�C�X�2ށ��J�\��Ј�4�G��#�G6�NѼm"�&r�t���Z4"�S��5��&.(J�Y�B�c�'��͎S�G��9���r���s������9���GQ!����Q�G7��60}vv���Q` Z���ʵL�Z�v8������nz���l���Ǫf�D�}Ȳ�v.��s���(9/N�x��D���=�W�&᣾�؁h��pCQ�G�l�}"<^��Lo��?����u�k�-yh��³$����[b�ݖ5W}������3!_VA`1�&�-*b���b��2���W��]��~�;G��t�h��I�Q�?߁����h�U
��5�O#�� ���/��ঢ়?ӵ��r�.�|����"�~���shv�{�T�=�ճ��a�lC�#uZ5	ota�3}b��	]����f������L���y
�{� ������'�ѹ��	�^�n���ͯ�
����P��%��Ӽ���wa�pI|�=_��ԲK/G�v��u�b&b%:�t����LKc��)�����lR3�e�鿡�~�鬾sCm�Y� ���C2G�ղ+�2:��fa�z��u�V�I�ߙg���Cj�>��R�+�ְz:U�^�iҝH^B�{Ω�Q(�Y#n�^%|l��4���}�̯��ۧ�%�U���
�>	�톳d8$>��0tۨ#7m�Qm1O���̛��UD�3Ho�zE�K�M$y�Z2�^���{����'ֻ�W�(�Vb�s�V@��'��H@hq�(1��(���nE�e��F�#����$��d[�q8�9옧4����L�Mڦ��G �k2'����#gˑaC��?�=�/`i���+���&���,v�ӽ����=�BÓ�ֱ'�雪���M��7|���p�ͤ+S���(r@l���QV"�_��Y��(�g�vK˯	�?@yo9��z���F�O��99k�_�|$N�Y�v@����k��-��R�,��WN[u�8��P6��¿���@�z��s���{IF'-�7� �3�Y�=>B����5�mԻ���Ư(e�X{� �X��c���q����Je��ŞZ�xl�"���^�v
�A�������4u��vNo͍�`�EW�˥��l��~|�ǘ:�:{#���.�ངL+K����G��#��װ�y�2�:��h���;"6�E���j5�HwQ�TV$�f���^��<��hW{�����g��v�Bxٲ2����A;��H�9���ğE�;��#l�B���*_~�lǸ*ײB�3�W�S)X�5�
Y?"��4I�/���;�� _�z�4�~��4Y~($A\�j��~�i��de�x�_�:S�LHS���y5�֮�UFd��d�ǆ[�qMh�fZe��QT
3��������F!;�M5�l��
����'�Dx��f�`M��x�8��zA���_a"%f`��vݺ¾D���'b:�C*����c�E���k�"6@3����\����>���Xy�$�I��U�b���;���Q�(�n;�#q���g�����f��Q�v�T��
A�0]�����������UdT^�J��Ғ��_��X�e��G
���ǿ��i)��b����!9��}��-�V�vNG,N�"�	�C~E� ��%0�Z3�B��g�������(�9�腽�,���cd	�nI��'���Vs��[�SsRcnޙ��:^�>�����Y��e>o��,��|î�ω��a��e>�@��ψ�l��v�Ǡ6�u��\V0(�4;��Z����u���Y��眚�f6�z��%������vͱb���DE�9d��f���Ǝ�2XHh1�p�h���׳�f3V����M\ݺ�Z�L��"�"�:�����I[�kkB�^L�n��]�K��e�^7��ޤ���s����a��z��Jɰ�+�ഈxP� W~O�H�Jq�0�݃d���#"Fu*�1v��������)N�Z>R��h�B��&l�.�շHQ����t��$�:�FL�v���c���twVp]��\�y�;��|���t�ֿ�t���[z59�6�����L:fJ9ݹ�u?/���;{�\c'C<�w�O�]���J+��CY?�B�L
dh��Խ���!U�L�r7���Ȇ�L��|2��Kd�G�_s �Gx3s�X:^����:Z�+�SM�ؐ�P��D��N��i���i���*�*>a'X�y�W��Z���ؾ�oS����ط��o�]����#��o�@kx�CM�3{�s����H�Z����}K٣���	qXU vάK($ѥΡ�^"9*����ܢ�m�0�yM1�����4����AM.Z\u��w�+�)���^'?�tTAG��g��a�*"����<���,���˗=!�m2��/�7FJb�PP�GI�F�%(StO�*B��:;�g$�1b���FF������feN�Щ�%U�6����*���b�j�E�+7(N�r��Cϕv�

���I�-��֏Z�B�!��?�6�� �mHP~�(k�vt�hꚟn2\���n6�}�p`hn�0E���/����/�����;���F�X#qr[@gs�=DlDF|�cg�;�L���}��R�!%xսa�X�2_�gIs�xc3X~���#|����m�����Zs%��ö�}tg>�`T�Ԭ��A�3���S���2���	(��/|�9�z�Y7"G����62�К)�,fLS�u� ���A�(����P�T5>]������/�|ٴ���wO�Ya8�r�4�P��Q��)nc5gӇK�:Ix��y�+߀�Up������F֟�(7����so֬ �����B o��#�i��|nW�}'�2�(~us��~*֍�A��[_χ[̎��[@:������g�q��J�"�ObU�K��w���A#.l�M��a!�������L'=�����[�5p�i ���wl~7lb��RrC�`�5w¶�����y� r|ej_��?$�`�W�(ZlT�\Q����t2=N�W��O0�x��E�(KW��u���9�yQ���&M�D�CH@\zM��lו�ǒPMe �t��k��>4�)!z'֔��}��a�]�?i'����{`����N��;U�~	����7&�(���f�Nm`S���T�!΅n_c�t�SQ�˟�H�H���nَg#@�D�P��"H��\�q������on������"Sz.H���'<. f�)�@��b(���qO7��q~�f�qm�zd�9��:���h?�L{i���!ɦ����"��b��r�i�`+u0���O�S��|��"y?Tt;,=���Z͹����!�@�I�ª�T~��r�c��K 	')H^��dl���Y��c+�D4�ʳd������"�If(Av�u(#�^���@V�:���r���n���p����e�jk����B��2���PRC�W����b�	D|l/Y�}�/�_&	�;13څ���Bܹ,T�.��Ѹ�wA��{��mK��N+����K�|����\��'v�㺃k�~��Z_;��WxC�Z���ݬ�jOʚ��( �o���P_>�U�yTQ�K������g��8KG2]1��WyJ���lxg��@]Ո��rl&r��g�bM��RoFO�&��F�����+10����}�o�������w���I�;#Y��*y
��_.g!F��7��l�W��j�se�=�0��� &� `E�x��5�ξ��WDi<m�N; 5Js����0��8�b����=�5{F��W�䧘��Q�`����݊
{ኺ��)����LC ��4!I����*~�DFi��yy�mPZSJ ~$My-I��i�W�����!M�!�[��{�����9AX�m��?�(�{�^�Zɻ �M���@�;�>Ǖd3�|��������V�H��&Ъ�u
?2,7���(�c�~�[wI��q(�6�N@6�`;g?��7��h\-X�6�ؔݹ�nu�J�/��W,��RǄ�}�����Τ�\5sp�2�0ڝ����	ߴYn��������)�ڡ�zD,T�$6į�ن���{�h�1�5-RR��0�y���s7lw��t<�p�liH>/*Ut��r؇
�بb��9�n�:���~�j0� (Gs�tf�i-&Y��"H�}z��.�d����3i�Ǎ���C�84鞖�>��I���:IpHCi��fU�������l�����`�'(�To>�[��q��[qS@�&U��* j�y
k\�O���TU�	O��S{7O�?���r��O�[�L����� �*JƟ�0�{c4@�9f�B���FUa)���&96��3��'69q��;3��U{uE(�(U>��.U��.��Ѻ�O�Y���������{�-!=lB���Γ.b�ɸ���$A���X+�4�ox�?Nn��D��Θ�7Ɩ��ake��J��qC�@��w���!�~���s�=���=ϧ:��k����q/��9����`c�B�K�韉	Hc�Ӹ�l=����2�@��1rM	�|s2�;Q"&
xP@ݾl�v(�Z��5���~8�����i��?c�r�lY(��Y>CƠ,Ĩ���ZMXzGҺ-¼	��"�R"��*�E�x��j��2�J�yC�N���vp�9n������%v"�Gϸ��l��b���*��!3*�Qߠ{��"�����G����fR�\;Ȥ�~�}x�E��Y�T�sy�W�+���4c�j����ٹ8�#�an�3�Oy�����º͈��Y�����"8q�����I@�=ٸ[ �Q9�M����*t �ۭ
�ǒ8���_�\}>K�+����%��""��?��1s�=�o,�O�7]�e�B{e%pae�%\t�A���`آL��h @�NHx; ��]>
界s-b:4~K`��#D����/ݗ)��k����~�?���^��o�8� �j���<��ȅy��L|mh���
��� �������A���.�S,�6-V�X��m��j�W?���5��r��g1��� G8 2( �!����3�Ё��h������� ��!� >���9y���G`%�~�tsǠ���"�[N�nU߹�0���<�ʪspe�㑷�>��%�+S�s�,Z=�e»ۅ��Hc jHj}�����M�g�A�T���Z���̽\�,��������!���M���DW�%:�	�~Z{
E}=�ZS���0��"���!����=I(���ŝ��~#�Һg���/���+��{�ܳ�F�Ť�$Al��6�U玬�_�n�/��~�ލ���/v�\��Xܙ�8	�3� 7k��;��DhǴ*�,m���� ���'�P���t<�T�������oܦ{�Z��tdcձ���8Q�)�ȕ�K�W:;\�^B�������Wy�����96���mO�+w.��;�z�g�&���¹U��_Uj*��y�Rv�V����ʻIcFW%c4�N����]���y�矬LvB��2��k�P��.�������n����H�6J(�ҿ�������&s��D��<��/��/p#
I�����|F��C����Jyp)�#��ʓ>|n�H�k�_P�4�����7/�4���*�9�k�(�s^!@U7����:Q�P���p���Ձ�N���7'e>#��T}�����5VM6;UJv6m�D �'4�aF�xN��
��ÒB��#���F��e,��<*�y��%{,L��d{n3GA�rQ�ɺɠ�A �����``�z����b��Y��~�& �*�\�:��!()�����c��^�8�^���Y��넦|��"�����Cy�u�u���"��98�)��!yY#x�\Ց�h�����8� �~�E�[y�Է�'��]�����`ZZ�_�ԏ��/ߢO�o�`�|G�1��?ٯ����활��^��4�S�}g�ж�Re﷠o��$4��.}���"R$5 ��Yˣ�!A'�+����sk�H�Z�xa�~��EB�l��-��˺3����y]�)}?�;�\]��V��7��P��F�>) x|�=
�'l��l�ms;o��H��wJ�CL6��4�����ʶ.�/�:*��gϤ�ZX�F���ǧ��/5U ��A��Ɛ�eH��Y&.L��8����)��#� ��,3\�1}�����Y2�+�k�d��jCf��sꖮ�If���ހ�7���]������Z�1
����ș���g$tN-���`��lI�"���D�7��y�r�iO�$�y���z���GbvXv8a"6M��g��:}�{�v9am�4g������T%"vu_c&��} �(7�'rq��p0�����	*v��"�P��$mH�)p�➉���a��� ղ��(&�q��b���Qࢄ'�"{O�E��	t���1�(`)�D��)}�3�T�-ǳ�\V����k`�F�s�u��x#�O�v�����d4�i���0w��j�o#�0 9H���(}H��4e�B�Ol	��+��5��S't��͓�� D����;��o���B����jw��Ye�XU�Y�r�~�B<ƞ�}}���)����O����gb�?�T�C<YX�j���F,9-R��}'ߕs��%��W���}��n\+�[�\�� �^S�˒M�/9
K����OC��+��U�l-z�\�,�f�o�4����ΘO	T���&�c6<��uӮY��<�̷m��G�?\ܙܻ�f)���èKj�nS�Ҭ�!-�g&���Wˣ5.uۧ��0��������w��˭�ҟ�U�^rZi�S������1z��ܖ����=q~"l�ȡ|��kX�c1�L�m�h�Hd�0���S�HZi�uMپl��� �զ��-�ƈ>��A
��fР����)�h򓙖�s���x�0撓����Kx#�b�*���l�T���8|�k3I��-i*��oFyBE�GF,[���5�x������
�&/|��o�S�,:R�y+����6Bk�֙e� �SA�����ֺ��8Q��o8�Җ:K[�K�W�����]�KGmi
놿'��f2k'b���ߟ6�Ǿ6-���?�(�Si���ޭ�ƒ�oX�^V7A���<�<���Kj�lA�r��%]ʧ�SI��?�!%��y�amQ���l��sfIg�q,��7��TՐV/���v��g�ō���&�u��H��(��1z�P��\�+���Ҭ�z��9��;kLy��I/��j�����t���oh���O���!`������8���4)�;�u��0�Sd9)�k*o͚�z�z瞫���}"������oJS�z�����7��F�Wȳ�#-�Ǳ�H'�A�T�#	�0�PZ�������|�D���s�1�e3�z���YJ�������W��]m�oy�d1���!�SL7��7.3�sk�*�Ͳ����8 
qhQ[�J���3] �H�{�i�n�l��hݺ��H��t<��Qf♸��./�Z]��X!����4�'�;�������S��Tk*Ki���f86�dn580<��S-�2ò6�