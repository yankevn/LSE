��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��?�I�J��x�H����Ŋ��>��g��{�oB�*�d�L�9�̮[�A���Oڛi�ޓ�,Y\�e'!�
��ae
ޡ��u��
;EP�|�xʨ�@���z��3^�w��>!V��P[,tƓ�{���x��\��/e�X�{rD�+�����a0��S;�zD�V�)��oԡ����[�����!�	���c��d2�3� �SJ�2��Q�z8_�`�K8:��ZV=Wq�D����O:7��m��X�f�����C����i�)n�`���7e8�_re�*+�H��d�M�\�??���ȴGN����fn�&�Wp�p�X�B��% 5�i���T�{�Ajɻ�W[dI=��Oc�buB�W
uq�wC��	�8o�.,���ɇ���#h)�~��Li?������ ��"Con�����r2��A]�{�0r��[{8��R�Dd�U���a�Z�d��K�>�DI�y#B�-�/Q���de��j�۳��*n�]	}���E��>�9������[�}��� �����c�~�
��(��S �Ӊ���fazQ�L�6�{�����Z����?;PV�-���!�X�M��@�!�g8�w�@h��Q0����ɦ䞨m��:of�QP��PC���CJ�!�	�ɇ����	~Nܞ��;q�l�pL�=;R!�ҾW!��+CЖ��9yR&��74}�[���l�s9s��ʆ Йm�#S������#]�M���Z�ﮆ1����7�}
�r(9Xy]����=������6%�\����!���-J%Ut��'��ܶ��&:}����@[#c�fR�������8	�;�Q�	ht�X$l
=8�7�.�86~1ԥ��-���O
�K���u{�D��c��I�Nv���\�Sŧ �^}%YA�C��\Ήʛg�3��MW��l��pZJ�����2������&Ш@ݴ�U��V��d �궅�Hξ�ӌ����	d���p]"d���0�x"�9;^ޯ�$2�	��^ΪE�*��7��ܢ�����"�#�l�������2�y�{�5j�ʏ�щ˓��oW���$����;|�i�T����W����I]{��w�����	��x��P�\sGP��*$h೦
qs׳8A.��e���-rؤ8
�e]��DG �G�bn�p<��f����D�z�r
^�tRw!X��Mz�u;�?����m�2��t��4-6ڽ�Pi����# wm"�[��#9���w�� ��� ��2�svB�� � #k�d���I@��	V,w�|����V�B@�샖)�!D���
�XǠ�A���r�e��>�t*F�er���Ύ�6�S� �o������oTX�˃l��`�Yx�-����=� ,��+�lH�{��V����"��6�g/w��˄1��{ݔ)�) ���B�3Վw~�q�|RnT%^���x��з~k�j}���b%�;E'� �3k�}5wݒ�)����T�Z����������ۻ���>�����O�+wu�JQ��N�߾��b7Y|�q�r�|8��
���5����� Kf�_���3*@��d�"N>�9���t4��j��
������@E{I\yM�e�6~y�)��*9�$]�������¦���3��p���Z:�G�9�N����E����S?L��{�Z�x;<,�I�������U�l��^��&)����EU�|#�\'�F�Å��e>��l(c���j�,Y}
�8�ZAk��4>H�c�*�(뙴 	%��~7a�k�����ʐ�ޘ!�e�[�5�����~M`xS�ӭs�h;fa����ݘ��5	�6�� �1%��g�^�:�<(q<"o%��=�ã�O 㗆"
1��+D
���o�W��Cw6Щ�̮/g��Oyw߁k7ia�-�#KX�����#��I�3]�T��s)�9�=��8�p̫E\)%�u�p����~�&���p{���%��.u�>v���WvB"��"Fyc"Z9�D\>��]	ޚy���&o�F�l�e�ce+<�I�JL�C�{J��k
��8mݡSS*U����C��&B�݇J����8K1yO�{�=��}��R2�A�WO���
�/H�x��a¥�VU�x�ЌJ�/���+�8i2���u:wQ'l1��bǺ�dA$�ò��<�:�vqkz�cV� h�;N���t ����#f�{U���ڳ�,^͂$���Kr��"n�=o��V#�[˻i2��4wI<0R�mܳ�k&iG�`��E��e���A�+���
[{Cs�^�ޥQY)� ��牱S�}i<�рζ 36hH��I>�������p:lݍ��/�4g~}�
$�r��Chp.t��D�6�������`|-@������=J���ɑ#BTr،9�mW��:sM��.�(�
yT�<�;誫��S��~ic/��+��S�l��ֺ�;1r )]b���.��}MN�ا0 ���|�����C�Ϻ�T�sҘ���VJ��t��|1WY�(so�Pt��k*��h�G+�f$�P�k���䦱n�8H(Mvs�:�O�>�ܹ��x�=��l��Ӿ�Ξ0������t� sj�%�����I���S0rȴGS�uro⎞�̄估b(F��ֺ�b�bwm�$0U�84X�����7�n���5t��X��Og�I���L3
֢K̈)�е�:�N�t/03�d�5$�����<��<��W��a��FF���o"�?0�`=�Ƽ����~=D��f���5o�����N�R��<� s��Yb&G��, �����6�z��,}��:�*z�܅�z��tA�����][��K�%7ooR���!efZ�#���p�(��Q?� 㜩 5�|�5���?d�\��wj��<��_&�zC
��=��(�$����8J��7��}�D�E�nV~�m��B�`��T�
�4Òb��� �n��D�B�;o��3�g��+�}h�\B���(�������(���Wdզ�g�7��ζ������ҿQź�{���.[t����tV�]�~�Z��^�h8��^E�v3�N���BWƚT��H�~�<��`�B�pW�Q�Vi�U�)QF�t3�`o�H
i��fr���3\�Ŗ�7��Ck���,M~��
'J�/ו�?t��KFͽY���͂K�J��e�E�}���q�xKL�᫦�	�j�j0i �H�:"t�
'��c�Qh��%�b6���A���2�y�B4��������]�z��:�A*�y�$6~�<�=V��r��|p�ۄ��z4��E͑_�صn��R��Հq��nX��+{��/@�@j(�od���ɹ��4j5{��h}�������4(f��S.:d���-�[���meT�ꭚ��v��8c�S��ib~B�X]����xr3Wu����Ƣ��7��~F[᳕������%�(�%K5��i
~�8���'�;�e�
�4��uFެJ%<
��mK����e%";�P�Tآ�=u[����OZ�XT�x��/���ꪳ쐞�`���]@n�&���<(���Df�t�����U֕�b��4]U��l������vq�E�C�K�WFeT�{t/���%�%Ǯ5@���;�q�C2��!�O^�=:E���T���`��A�)��Y�$�^wJ�'�_��UsN�Ɣ3�Guk�5îC�{#�=�����g�z�9��~���uX�����KsN�X���=��e� ��H:���Ee����Dz�2��q6�&��5R'�v��P�r<�8�������N���A���B��o����.���z������И@�������1DU��ȿ��F���l;��D�ҏ|��Rw����udp/:�!8������=��  ��C?�� �Stm6���	r��O2���qG�Ǎf
���lF�����Z��Q�y��p�%�{%��ͫ��
76ե��c�)Ųr͟>����j���r���ǋ��ߡ�"u���MRCQ�$�D���3��A�O��MR�)�Fv�U-�@w9H=c��+��,d�����F�z�w�y������oD��yۧ���J�p��:��ɔh�)r�I��=��qLk.�1��_�\�:��ȶ�q��x
K�����\�V�F>^�8�w�~	��T+�`xm�Y���󭯒@�<�y�]�Uuz�B�ۇa��?[����X�s�Gŏ�IW��|��I&ϼ�8֙��f&9+��0:?��S�n�6�!�G��~�E�:z�kj���E�$x�e�X4�/���~鳭�O%_j��*�:����s�廿h�=>�m���:UÈc�:�Ej�d՞	иd�4I#�F��XL˅*|��|��4��%8��*Ս��*G�����\<�0)3P>%_d�gr }��,��u����~+�;�Ѱ�����O9�`��}��]��ܤ:��V�]%��/�D��)�� /@����t��&T<n{�����)� �XH�4�f}�P�0��Xk9H��5����5�8� ݄w���8�����<�������FɮgL��N�g�jB�`�b�%[�	{�uHw���G\QaÉ�<~iY�ƟS�8�6�� ��!�u�(Qʩ1{�M��Pސq��j�����
�n_�1�1�#�E��~C_�(P�tll湥�jZ;�8�d@,���{Wֱ5�oN��=�չH�"��z�o����f�?ק��r�E����Y�����d�6�} k�QYdPw����'���[� ��N(�1��8���V�Dǌv�G��q�����zL�j�R�Ixc�������70rʘ��e����; �ޑ���z����M��L`�.>or61uJ%/k4��!��1�{�Ǻ����hw���#������6c_%�$��棤�K�4���}�xp�9<�o{�a53�Ρ�(<��ۤ0��z/x���Զp7�]�0�U<e��L0�Bֺ<�0c�T g�F�M����ӷh�Н�8WC�tɤzY�d���'�}����&�,�?wE3�豹�����-A�5��0f�"�qg�aY8ǎކ�?�2�E=�ޏo�����[=�s*	�'��Y���u�CU��b|87Rq�x� B�x��I�?7�`S�1q�m9y5�ap$ˏ��zT�7X�)kdB�1�Ƈ�z����a[� u����Ot��E޶�y�i�C0HFHqpF����>~J�Č�*��M�&}���jJ7w|c1��~�,hK&�LGY�q�x]A�uq��a��'3z4���<^����X`!$��T���SZk!-�����L��_.@e*�n/L<&�Z�ȧM���Hܿ�O��}� �cs-`N�� :/+�:˽�e
��4�ձ2�
�v����,��mN�9�2��>�!��u��'�.��
�������G���A���|9
���b�ޡ�*�q]�ܺ�����=�h�1V�k3@�<1�ٸ�p�e���t{\ d���q&Qڞ�
��y�u0(�XF`�/�X�2p��X��X���9g]�D4���cg�Ө~���������4W��x��3�п@J$��>�[��N�0����ͧ�݆>D纁WYEDJ �iV��M�N]�j�҉AS����w��hE0��)z!�kd��z��h����YUd���h��he&������1���2�����c�� 18)���Z
�^� �gp訪�j�r�7�ٳ�X�&��2+�ix��|��y8]�-��E'O���[�+��
�=P�HT�hA�����J�H���B�J��d�M���p]�]�2]>��2F�̽���-�nE�B5fE�$�`�����O�����i��Q�5bb�c\>�GoB"D� �+L_e���+�_ڃ�J�SH��e/}��ݵ�PT�د���-6��<��=�#1��
W�u+k�Kʞ�/�X�����q�����饂�l��b���a�6T��@̦O�֧[�~t�w���(��O90����Y������S⅕�/�Q��	ޮG�T��#���I�<��+�����G�� �B��xf%:��6���2C�U����K(�'#��(O_F%�l�w-�׹7I>�@�'���{rC�Tn#���M�-o�۫��o��U�<=�9��$(�������3jh~��q���з}:j��G��t����bo���&�E�P)��j�:�^��\TN9ǣ�;O1@�TP��K�rM�����X8_�#!����OU��x�(mPom��g!u�c�� ��Zx��c�KE��ya��Q^�	���&�S4:t�s$�-E����A�=��(�I��q(Z��l&��^�V�858}7~!~��]��R���4j�b���6�)��U<���+��.�Ox&��srXvh�l���_
���Q��.�G�u��6o2�G���Y�����Y���4���3-4�93�DM����|��A�� q6gw�Z�Y"Wrb
�	T5wj��ԃ�_	7sȞlװn�AdO�z F�g��O���r��H  ���Xw�CbV#ݜ��)*=�� �>6�k,;ϗZA���oH��y|D�曫Lh�t@�/Qcv����z�e͟���^��	��*uI:��{�-�w��3��B���@�'��i�t@������{�ɹ�@�?Q�n9����m��A3�5.�TR�'=kZ�V���1ۈ���j��~k0�����8	غJ�RS#�l�f��h�Z�����.I�$/���͟�L )�i*�)x/��T)��U��$"rA��t3��3�z�A�`�C��0��\��g�F��"�r^d��Q�#G�2�xh����@����*��ٶ�͑�?d��I����c�m*װ=��DJ�|ث?OW��L�ae�2��|r��8kg��-��!���	ml�v�c*$=��ϸ���gIR��N��d��t=o��V�T�A�x�r�`Ѵ�sTs�#4A����`�˄���"��ʹޏ}�EV_퇈A2��J��/d��b�/�-׿�^���m{�M��j���h�
t�J1�Y��jT��ɍ|�_�_U���rU'���tP.S�a�תՍ+���i�^O���<�7�Y�����y5M��?���	���Ŝ om���%
U���N�n���1Xӝ�g\�N�^��ujQ��{(�!z�{��Њ�O/��142I���[,����z
��2Z�½�f��QL��> �������+١�@'KDm>7k���y����@�i�����b��	��s3�L3�%eXj(a\~A7�Q���Kx�����}@%-#,Vm7MT�������Ӌ����,.��Nwz��O'a��ğ��l�����n� H�,^�`���aY�<���5��k��~��U���;y�l���h�ŀ��@B���Pҕ���na��Z��r�NS\D}�GAZ)���Ci�j��$4V�^��r2&M����W/T�勅dJ���b�V󨎛�*�n��{g !t�6��fk�����;��$�Ɛ��Î��S)�8�^�C�p��U@�y�.���F%��h�Eg�@���Fǖ��s��d���T\l�х�\l�1D�UO�����<�[w�pO��`���/FA>�2��Uψ�#6i �[��T�c�
��s�����!�F$ߦ%d����ѽP�W�<�(+/e���W��qc幩��mE� mL^����`~N^8�C2�]�Fq����uy%;L�S��ċ2�Z�`q�� 䶬��9.R�5\kK�ޫ�Z:����Ƣ�v����m����Ṭ@9I͈	s> y^Vh�֫4�������k�h��/p���S(�
%1h�s���k����,�;�Xl�A�X�`�L�5��#�`�8\��4��̩�0�Ҽ�*!6{k��Q�(^9o��Օ��&J�9�7���ψͺ�{=���WW�������юS K�=0Ѧ���*��-/��9̖-��n�!i��]� ����L��2�X�rX\"�5L��8�\���Du_���aM����ϋJ!sX���n<o��P��w����i�r�چ��7���v�l�&��
�C(�i-�@�<���p�"�(e��4|d5��c�``ÃЍ��9���u%M�͓Z����5��䢩�Z)����5C�c��[.6�!�D�N�qC��3egnY!��s���u N��><VKؚ��sG���䉁B`.�49ίDi��܊������՚��
�����Q��][`~�o|�_{����'�n����A�y�&��dzo�6���z��O�L����Л_��]I�01>�b	����7��2n�3Mh�qWB��gh����Kdp(�G��0U��_i��������6q�[k���Z�V=�	W/�
+=�2���# :lO�Ǭ~�ޢjHx:i����*r�=��I��f˘����z٠}�*5�6�Ϻ���m��7v�@Դ�
'u*�;rrH|x+��$M�E����x4�sh�%F���&�U��B�%�P��y�b��� f	 ��׎��p8��� ��-�(�5m�諾����t�^���T ��h���F%dk0ykTؐ�#Π_�_W�T�����׹�����ӄ<
p���0T/�G���㹫ƃ�/;�z���� ˝g���<�?=���r�����N����^�KX�5��1t���O����(_�=�}F�l������|7|�͈k/{�H�q�L�x��HR�y���s�����vQVϊ�N���I���k
� �U~�;�ɼ�?�j�PC+`&��~Yd�Z��dݖ��Rʐ_ͪ�:A�C�j~��V�sϽ�rdW` �0�	cw��<��q�DXp�4�~v_$t���W�}���I 7��V�L����2;x�c�0��K+�;�j��
�#�^E�:��L�������^<8���h��o�w=]	�LI����5�'W%�Qֽ<��"�dYd��,.�
�4��M���K(�qZOJS�w�m��;����zo��W3�򐏾�ڽ����a�@O_Pbgiq_2�z��#O�*�u��yh0 �h�PS����tt\"%���#�:������J����6�N_w���1�
B��dH�%���FM���$���=�ҳL���uǰ��7�hk�lˈ�#M��Q ��K��1<���2����������ӹ����K��kr�C�tW��*g`��?)c��ъt7��y����^qd!��^��=�%�?���,t�V���ٹ�����Ӌ��`Cj,�������*4|N��=	��� ����z�X!�C���8���ݫ�`^^�|���oq�h%�>�Q|�E����c���Bm����~�gv��:�}���(F��ƌqu���ҵ@���ʽ��K�e��i��M��
)�(�EUBMG�V�ú}Õ�}�M7�F�D3<%s`��v����Ek��c �{���#ʝڠ��̴���;�8M���tY@�]���j9?�4J��Q�=�I�T�0�����#{CG�I�V�,t��E�,@��;m~��H��(��GU��|eS-V���e˼<Af����7 1�F�u{��}�"xM���c0���{���t<MЂ:Q��;ٞn@�."�v;�n�����1�)L��4��8LD����A^�U{��!Q��U哧���>v�%�]���6�z#;v9�� o�*���R��W�)��d:1������I�R.��`�ǩ�D����9翇6:�
�r,��,ä9cۡZ%��-鶘�:�ڊy�о��g�w���N��v�?<�F��ڿ���ݯ�~|x�U��>�̚yt�S���MF���Y�`|,p��"����hYkcA�p[��r�؂�ӔFqy��*�J��]��<��:��O� cY@�t{�����QW\kw�,�R���Y�h���kn�7����V���6q�R�D=X}�P�쵑s��ɶ��ƙ���Qz���B�-���k�|�V%�	,��!�+u.Ӛ�E�Ӄ{�T���K��Z��= _7��&h��w%`���~�W���L-��h�&���������z3�Q3����}�4���x�V�NJÿY�Q/�Ԩb��쉚r�,�����֍�;��䚢��� V��K��5�/�����3/h2+�A���G��@cTP��L-8�8���g��}�
q�F�k"A��b
KB�u��܇g����s��n�Yf�9z����='�k��!�L���$��S
(b[>jSq�rg�P�l95�W���`"��`��H K��/��V���s<aj��>��a1��^7ç@j~v<��a�`�X�T�GFr�@|%-�����r3��{Q%,Ӏx5|��O�<��ZΕ��|zx��/,��a��2�/{0�W��^�m�`� �ؙMW��\�d��V�N��@��������
����$��yvt[�@�7N}2й��1��s&����D�����2qr�2��⼄��+��T͵F�W�xx���\�'��$�bIVE����	���E���S�B�4�]:�9����S5���J��t��Y䪽�ڿǷ�.��\*<�ܤ�e����ѧRmsm��B�����.��^�D��N`n�ɻ�d��,'f]obZ�e���=O�1>�Ľ�:�SJ����������I�~�Mh�t��޶99h����l���&�

�S��ɠ'���<NX���}�:�VFV,(y����FC"��� �BD�t����M�5�&
ZM�{@�N3����N�d��� �`$5Ξ��N�� �t����3�߯��v@�﫻��*�c�N��/����m����&�σ�����~_���>���`���ǤL���rzhi;�| c�%�Ʃ�c�ğ�rb�"��]�&#!��W��C�
'A�Z<�;�<
}@$B���Д�>'�suh�1���$��}�L�yY���5���J�(�[���H}L�O�<1�Ҭ��2`=����Lq�/vF���ֻ��pUò�]C6;}&���K��D��J��#u���>�,�͆.���C�̐�6�!��^9����l�DG���Hݨ�`����#!�fq���3�A�cP�&�E�4O �E�kxV�}V���.��gU	P�HFRn�)L܅|��a�w�������j%U0ݫ<��I��/�`�i%�i�_��Wt��y�C7���<�ٵ��m*��N���'��I�мT�K}�y���|%~����F@�	|˧Bv�ʖTR��0_���+5��i����q�THiE� �V{�Zs�]�)3�T��#�m�������G˽UѽM��ԫ'tq�I7onqU��[ƕA�d��hR��te�5��9���7���D���RC���;��a��踹>Ɗ&ʌ2X��T�˿�n�6B��`����@aҏ����̉�X1��<���#��?����H�$ط�9��uA�]�+�_��&�|��aŁ�HD=��b7���q/hZH:=�p
s�n,�D�_�� ܙ鑣,���ߛ]h��? |9�7;����y
3J8m�m����Y��[M�E�?���IO0�~� �
�.i�������ˆ� ����d����3�}3*�|�;���h`
e�4h�l'��-�tG����m��cW�cQq���I�ZD���&���G�֐os{?W� E��Y�ac;m%� 2љ8�w;�?~
tltԾ���x�i!����c�ojN����*4��ykƧ� !E�5��L��=iH&iyE��;�݆ʂ�t��G����ɝ˟�ս��U���7R��&�|��6i;*;B+	��[p��(�0�]�08^�+e6���Ѣ�̤�Go�d���Z�h?"����і-���N��}�>�f
�2ϰ��1�掞�+���q['��.nq�A���H�c�����?pk�m̄ƫR~)N��QT�RG�G��f��E�v����wnhemәͷ��L҆VM�Z9�_#�����r3˂J��մ��~�-Vc����3�[�[P,���:�7_�`��A�C7b�M��4���Å4��[ �ȁ�~��1G3^c6�1��!���<�~��(k��,�me���E׃�d�Q��j�8Ɲăݙ����w���١�R��*��d\�wB4,!�,��*�������V��/i�Ց����j��¢���-g���[\�@����F)�ʲ��G8�$�D�`���n�V�[a��RP�����j־�2�@V�}��d�d3T��]��/�7�9��G������d;�O��qL7�κE����M�o�S�!A�"�"��SKpU���Xu��'D�6ݍ/͓���l�i���"�]��b��Y,�EJ[��?�dg�O'�ԇ�=����5�!A[�+�	�8�Jէ�� �����@į���+1�JWb�t߯M�% ]R��t�ʳ�"�����vހ@�	�O9JK��g|v�����Đt::���a!���vo�LM����A�!�^8m��#���g0�O<R�n��_�8
*ww� �Ô� w�}Q�ъ�m`8o�1E�5ދ�$ĕ�.��#��=��Z�+Q�?�ջ�d�^����x�ӟ]>��q�����B�$���pO���A(��準K��l���Mc��3��<å�T�2�j%�&����EX6� �pI�?�����.f���G�w�e�z��^�e��p��1G:�L3���	A�M������`]u�7%환����,N����f���C%$��̘Uz�4��Ӿn��d^vPy��4�mzlJ�:��F)�	1{��u��c��G�K��ה#b�#$���3����C��Pd~�����;{���!�u^� ˟>xl�����e��'P��
x��s06��,��7�Z�pt��K�M??ڊ�qQ�����|��ل��O�
֊�PIt�M.s�B!f^,�v�Q���-�*�����G����D��n�/�hz�t�*u�{Ey���d�p�<pg^Kd!����E) Tt��n��`�.�+��;�S���3�Wd�����lц�$���'ئ�!�b���W�;�	���VG|ܻۖ���%�!:�03������5>�TU��ō����
�D	Qr�?����w��F,P� D��Q�d��\�EQ�EIkH��4��R���i++%�Y��S�C�����3X�-�Yf��V��c\�+�����L���v&D�Ʌ���q��"����;�m�"ЉYvQ��$������a8񧇲2�"\�%��PY�/Æݮ�r۝��ZZ�v/5XȰO��+hz������r�Ȥ���$:e5�7l�����DQ���+W`�mU)|���xa<}Z�P�|~������߬P[�g��/����xv�`�ѾH	��t�`g�`�j��\�< 8��asq'�D�c���FaC����+�n��!
�M�&��Ϛ?VB��^�!E�YXje
|�ij�:_��Ы��c�:�Id_hWS�R@ʌ��`���슏1mI��h�}7��'+)����E$õa�X��`q��Q�N�	"�/�j��ӂ��.Ab�Ǚ�r�;<�!�Xk�������f#�x�S;�bTA3�S!�J��T�R�wVWp&��#)PB�Br�C�����`Rxǆx�<�� �"���/�r>�7V��^c��uu��%zw�<"5J̐��P1��@U��ǉ����������@��8Ze޺�z�~r;e�*|_��J���5w��FT��X ;V2�K�r�G��,+1�z.�N�F萀(������h��Hh6��f��q�3A�L�G���k����jn6�y=�U�����K�>B�cҜ���(�<��T�"��煤J6��t-�~��U0�xbg��C��Ќ	󨔹��Ғj�g�ܛX� 1���ʳU�Ɓ�����&X]��X����� ���䭸�C�x����p��ŕ�/���cMm��܁���Jq���sKf����DV�P��S��I&��c�QB�x��ȍ�����]��U��d��K��ac��<+i�v⹈}�j���b��.e?3�?�	T���T���ԯֽ�������sQm��\5Q*>i� ��0$�\Յ�V�8�2���	k=c��]����n둈��b4�4HҤ�ƪ��f�E��� �m�Lf��E���e|?�)5,8$�K�k�h�W�}�j>�AT~P��hUYj<��]�w��Ì�Z��B*!w���Zp�Gm�N�"�t:Q��V�Opu���E�1�Y�e�Qgs]�V	'��"�2uåȑ+��r�z��	}Ly���������C-��Ts�[ZW(Qz�"����g9S#m��`D��/\3@ŢƯ~�ۿ�d������}����n.�-�5sѭ�N�ԖmJ�����M�EV�Gb�s�����gjg4�y�/T�;�6���>��f�Ns�Q���c^ ���zCł.,T�fd�s�\t��Anv1=�C���B�AT��Ԭ1jI�c��MV��;nÜ2��+�[kY�ߔg֘��@��j�1L�ε��K��r�F��^�c���:"eb{:�[e��vΎ�&�6r~��T(�ŝ]�C̦r��Aڭ.ҁ�-�f3����O^E�&2�*_��{�mO؍��#r�4`�+=-Ź���V��ΈǙm���e\!y��s�����0�u�=:.w��I�֭�-�E�͵��7p�0�{�ȹ�!P�Vu��頉�Hn��{D#h�ٟ�v|�(���
����NJ9��R!���yP����i76,���p4%�}�&��/�g����o�v%����p�a�$�U��Q���c�؋�����^��ϞM��JQ3Os�\U�漲���i2�$}�}l;��%V���_)�cPU|�˨�h����P��ܳI�1��jcoye.��VC��3���B0��R�;y>�W��s�*�e�y9e�c_ Jz�o ���ߚN�/�rf�)
��q$���z�7a��6�7���`F7�Tkd��HԦ�l�Xb�'��>v+&9���$�(k��#>.�o�3��;� ��C����%��y��,�i*Dt_K�#����'�կ;4�q���Tx�~T�Ivt���x���S�N��o�Ԯ���m�~>^h.&ϕV���7�Bь�* gЂ�|��0j5gΗ���8�JJ_�f��>�}oq�-��9��=?�/k���7���fQO������� �ǐ���[4Np�l����7��@T6��Q���V9IVg��T2���M��-��0þ�"�o�,�O�r���1����p���u�e ]�� L��� ��_q��)��|t2��͕���Ε]��bd~�ɽ�Yl�F!��	b�#6�e�M��v9�5fy����b��'�iP5��^�0���V���e�_~��3�zWF=lM�_����W�M?�lr�(�ŜƲ���j]�붶C�6�ޟ�kgl�<}�N��H���;OAxU�(����� n8�?B�ǀ�[��O����49��aSm���lt������~&�6�S�;E�S揟䴝��R�滓R�g�{�\�)4���A{��"�_�+�C
ۣ]�H�����
1�nd�W�3�5�����20L�����\V���|Ĵ�Z�l���B������&½��(D/� �!AC����7���-�H7R���3Pvi�BU��{�iN�]%���[��"��!�m�f 8���|�șme 8��3%�0>'2�w�+^�4\QE%�M� ��'$�tyz�D<�:���������e��-vS ��0��[�(�yw�E`0��[�^���g��֪��ѯR��y�D=���'ɸ��k��x��뵘l��<Hnq������3d��t�v��(Μ�jD�	|��ĵM�0X�uM�b���:�w�%�ku�L�aO���$����X�T�)�a�{+�����o�x���P�tަ�$;����;�Ѿ�>Q��mX+:=�by�K�U؈Zް��#��iѮ��|��1�B{�Ip���7�x`��	!w�3 2%.�aap�FO�G��5���e��,��?�8c��x�M #*��^�3��,�t��3a�7�z���oS��x�l��qE/+�MXahB�^�h�]<�6���$21Z��	Ƀ*���!�m�]ؠ�)����&�������{��ɛ��T����	��Z�������mcI���dG�%B�|@z��� �mM8�2��A���6�-�W�_���@�|7�q��d~�W�~�9S��]����t�K��~�8���t�Ր�N8)��������{(1 �2���E�䥕�7�M�1� �,����o��C�I��+�T��/4U�+2����`M=м��K����K����m%�ҝZ��������%=�w�M���B�f��O��yz�l� #���ѥ���A|+�Nۇ lk7a��nr�[��j��O�%��^��ߒ*+���}�l1��R9�m�?��)��Y�]t��a|�Ȏ��{�b�s�d򌨅}mh��q`X�I����
i��"8��^��s�����M�o�I�-�Lq�¿�����Թs��{�1�^��T?��df	:�.P@��i��-Y����v�d�X|�������+X�M;� ��-���{Ax����f:`�@��<m��k��<�G���`��+����շ4m(�{�V��x��B���zoI=/�D�_���N���?���^gA�OL��y��/Ɩ$�y�.��,_�;Tk]ͫL�GDd%�+B�X�P�1�ϕh�t�,0���g�\w�r�>�&o+48/��Vݥ6�'M�|��#O�8A��E��|��j� ��.�dY{�C~�[�N2AD��+
0��b���`3S����ɛ;� ��di|��(����jC牌*'<B]�\�8�9�QZw߲z�VB�M��$���U���H�m|��`�b$CA6���ָU;���Xң���������4إ�*5�~��� �H�2j���:�\��P#V��+����o9#�-�������Gߴ�_����~�4����ţ�x3EՒ�)�l��ĝ����p��	;!ҷs��H}F���{�ղڤml�tLe0��F��d�/Rͷ��(m�'^ё.x��#���^3uU����42�Rm:�˒�����/�Kg���� P}�ȋ��im���/Kso��q� �?_=�}�A�Z�8��ְW�#��e����^�Mޒ}ꌲJg쮙]#h��vu\��e@��Ku���ڍ��9�����g�0�Ox��#�L��$l�
����@S����=G=��Ec5��4��0Ҧ���2ϔ�M旒�3���9�`�q��bb3!�g��<V�J�| s�"�h+���
�b�@K�=r�ܹ(�Z5���U�p�Z޽��r��wSE?O��&}�u���]�Rif��Yq��I�äRZK#g�I�
u_���z��l�t5��)g��c|��<��'�)^O��%#�Xn�=?;���E�z�cL��L�CR5QR��"-��[���(�h���1���!��/�@��m3�n�T_��P<�9nԍ�7OB��t��Y�X��SLɀU��TV�aXJhk�(=�-���z1�wo��Z���/��Ѿ/_��F_B�cWin5+)�8�۰*r�Z�OW
�!>����@���E��ýa�H,С.��7�鉴�z
�/�`<2���E���3����CP�9��Q*S�>�%��4�%��(~M��QG��_��r��Ϫ���;eܤi .�,�����#���C���S�:�xq(��[��WwF�g���L?%���&?� �w(e�q #j�x淊�C�_��S���=p�&��$m�u����$���F���Jt��f��c�:�ֲ����?aV��<ܭL�}�iGM��e��%�u�=y�vtĚ/�i�����L$	�y�0� �������ǒ�?���b�����p�Xx���kOf�Sp�}����	\����D=��0+iq��y�HJ�x����I+KV�X<��a��2C��ƫW�o��
��&�V	�:W����:�7��3�uVД����-�RXw!ch���(�+�=� ��^%��|�SQ-1��ܵD�MtDq5�Q*��I�q�Dt�7�hHpm{�F�(S@� j�� �f�CyR�'���Ъá�٢��z�����'T�LzߜP.�4�0�U��SD����Wna��2�&Yn��� ��+î��zG(p������І�2�6/L6f���n���5���U:'2@�`>��gz��$��C|�x�T`�>R�. ^�V\��=?k�>q���2��l䈪N0���$e�����h�̙��y�5���r�BM�W���D�����6>�/�S�"�TpV��$}�S��Q ��Ѣ� �U�+k�����Ik�H+�L�C��R�nֵ��k��S!�(���f�忲��-�߶�S����3�a�=��B���!	��q�h*�R�="���Z��J^�U�"����T�H��H��/CUb��j�K%�IlZ���=��h�i��s���p�e��@��&-v�v=�#-cx"CN[���K�o��VV
+HO���^d��f��L.R�Ǣ��sf�`LXN����5V�.���E�s���r����f�
,2$0�Ol�|��$VYJ��. ґ������J���|�#���h�&i)���0�y��B��	�T��� Ј�i"��$%_Fp�jo �RCx�I(ŋ�T�R���ƺw�!2��^��p�!l�V�I:�������l��*���Lt�<�)�.l��/�&⋒������6D������A�{�֍G���M1+�$�z<6խ��$��ű����&el}��[�d����ZE�~+�3���'����B��3�
�ʴ�ٽC&a-���j�����H�6i�j÷���Rֳ�K�kD@��ؗ�'��c�*�(��2 ����s`rG����i����YH�]��-���̸���
�.���1l���}�+��D�8� b�Oh�1�δ�����Pa�B�v|�i߁�7,�OJ��P%�2Ү�c)����y�!�������"����V�^��"�tyv<+���;���^�����|k�+��|��M}��!������IZ?,����Q�L�>��;I�+�u8Z�u�.�21���_v�)1;me�q���/P���$N�n*��@���[�u��Ԋy�����M�=���e���.sr+���`��7{��V:7&�Y��z%�æ��N��������PA�۱���/�@D�Uu�@�}�X���E�5��]�Q�����A�EW]�!3 �5*\�l�)e���O��=���>.展w���a�n��T����4Xym�����:G���=R�\�Ҷ�8���q�,�s������N�8�N���WZ��Ѻ�E���w�+�=�65db:\��H��Gv��5��bI wf��ckG�^IYY���~�~�i���Hw�D�7օo ��߀~�T������(;/ <�z�0FҒp9d�K ��,�� ъ)Q���� 	N�-PC�i�/�W���Vɿ�*G��T6F�J"������\�j^�I��b�Op
SJ��LP.���sރ.O�e6�Hc��}�[�	���kr�����'��$7�fO=�����4/�$b:>�'�3�����3TWz�^�o�m�=>�8E���s}�'��~�|���Y�E~���t2�=���M�F���-d�}�ˡj�Q������r?I؇�w5��4E�S�.+*����B�.a�x?hR��s��$�G��=�{�u��$:��jՁ��A����M��d(>��sbX��;
>�S©�x�s�M�.��gG*7�̬'D�����A�/�(lq1:Y+l�����VH�1A-־�������w�%��g�ECN�EaBlp
w�L�s|���wB�s	T?��7i��_"`��>wq]�ʣ�+���[`96��\ ��kM�5�䕝D�F���Ì�&#؂���b���g�u���vdZ�]�k�#��2����zuۻEK���dy�!���̺ϑԭ��@��rW?M���^Eh�>�Cu��0�*�xJ?ac���^��@Ly����Sӽ��9M/�e��A�j�����#��D+2��<����:��%o�V�@���t��w;��1\���m_��+��J7��I��W<���^��C��Qѭ�������0���نǿ��9a�4Hu�$��U�C��>��S3�T!���a��V#���q�i�,[�7��$ݼ7���|��$b���a����b�Z���q�e�w	R|����t~a��O��uK��e�g�#�J+��F}emڣ}_��_O]������p/�z�(y��
N	%c�`���9��	�?K1�p��攆�
������x_���6�\�7@����I���RF�8:uU���zG�;�7cJ|b�����a��xҒe9�/Ɖ�:��_�$�$��)̢��w�֘��M�`�r���uL�!����u?�lN�2,ϩ����?�t�>$a�]2(�|s���e����_�x���uW��z\G�x����5��SoMg�6�7;����Tq~�m`�U4�GV�v�0�kT��Kt�I1����zP��[C��&��)>�Jc���4{8��7�j!}C>#��l�\[E�x4?7t󿝟���I�֖>��~K`r�<���I�v���ܳ�4���.�K	��"ŭ)�S{6r��X��1�Ț80��&�{����p�q�~o�U����@	��"�꬏�s�Y ��(f�m���,�N�;�;>�as�v�UC�^��l'�P&Wu�i[\�*ס���~n.O��)��kz�+���r��y����.B�c"pu-���#�p4���1!���Lj�o6^�j���G]��j�R��oDwl�,�_������e~	"�;�YuG�!gE	�q��)����0H�K&�8���]��*Na��3�f�c���"��Ad�i�>��E�&�gNroH��GLUB4�L���m�m��
D��,����u7�����4�g��2\��j�Ӑ�Du^+3T}�ij�M0"���[(���!����ڃH���Q��~!����B*�7+lw�^�`e��J�;A�Qv�Ǝ�3r��Cq����ĸZ�om�O�
�֪�;�c+��I,�E���s4O~�O���N2�~=r�����.*a�1����Dt����y>;qq#��g��EV��F�8�QW��䭘ﹽF|[��Dm���;��./74E���X��3�K ��	8H����*/'�SzI���c$#߄Vz�Vj��q��N�?�Bת���Ǜ

b�\���]D�$o'�tu�Z#���	�g�/UW�=�~��]+o�k���b��>�K��_& �K"�GdD�p�#Ȕ����G�ވ�a~+��O���k�:V+��p"�.��SY��Q� ��\5�{(���)�����3_痲/�������#`"�M�Ci��s˟���������c��Ϲ�'7ru0�O���=�x��V#��d�Vے9��4�.������H�R��g�ԩ��k�q�k6R��]k�g�wC(���pY�Uv��8-���)eH���Wɓ���'s�zv:����D|����sUy�.ط��~�v��B �LP��I7�_��[w*�����?LG�C���n?��vւyv�;��Д�^t���V2�0�n=�G�l7�<�?�B��|[Eq#�$�� ��5�|�
�2:�9D�"��x�?��I���?���nf�^õ�5��
�v��+V��H�Hj���%�(Z$0�uꐁx\����%��1S3Ѿ�u�$WE����4UbO�_<��>T�g=NTE��3�]uN��,�7��v�p�JL}ْ?�֐cq=(\ǉ�Q���>�*�|�2q��P�g/�sd\��x	�\��-_0�*����n'�ڔ�ۊZ8�IR:q�QN���>i����S\�LS�_+�����*���3��L��������
U ��GP/�i��6��v���v��y	(P�ȕ�3��� {5d���0F�0�����@δ�OA	�!��ѕ��=+�}�jwX�JP�)Ƶ����l�\G�d-+����i�"S��<��Z;뼋h��xy]�� ��o�_�� D^����JocJL�crq��]@�g�i2 �:ŗ�UQO��ډ��4��Q�Z�W���Yi��(%_���\][�M�u�L� XZe|h1;L��E�?p��Z��b/i��t��Y����-T򿱫y	�o����Խ���o�p�.�0NHʷ讌,�&bGXE�����	Xf��р��ӆ��r��%��Vhw?����a1g.a�� /#�	�	�»�`��C"`�[UZ4��?)�-*�!��kŤr�ݡ�q��	���NF�#ՀaР��W��e<�o��6^&qI����7E{#��P}��)T{?�,�E��_�[,Y��Ѭp>c�\ +@���k��8Y�9+U*b�ȬAь6�W�P�7��K/��y"��3�H�TF��d��X���+_�8�r� �{�ߧ�\�[�prWI�z�^����L$"7�M(�7�r`YA����a6�*����V|�$*�D������b�A;	��e�ky�>Jz���$dw�k�j��%1�J^qp�0��4���Iw���{y|�"�65/dcn����L��G0X�0�t�Ći�6
nku���R�����BK��iV�F���X�<�'K7��
Eյ���c	?�o��ޫjx��2�~�bP��H������/�[�}8g�1�>���ą����vB�;�����sO��6(��7/S�A*���[��+yE��e�߁�)�舿�7tGU��l4�y��(�48�	�7j}P|S�5?��fj���U���醤������b��8hсy�v-�����!���9��8D����%�8��}�Nt��Pt�Z�c8��]h�?R,���� 'f��T�0����A_1�Ⱦ�Vf���J�
�<�Θ�o�0+��Lu��E�
�|32+١V+&�}/*��;&(�l�[�f�MT����2���c��1�6:��(�ل��a2�s;U�-�զ��vB���q�{N@Yk�0Z��S�&�@���B���k.�+�)S�^�Q�[�Wωo*��ӟ�4j�"¨.���w��p���`n�>+�5P���^7D���?�����fA?�h-_/@?u4�	�M�͇Q��s̼�*w��7��B�^���b�z�O��]B{_\�T^�OIHK�!�}K�ŗe���3�#�ӹ�ZwC�V�a)�'@!��v�K��"U�7'�J���� 7���6���L#��wxK��(�٣ὺ$�@T��*�Zݻ��A���7��eD��JF��KL�Ξ�X���g��Yz11��G��������fE����2J�Z��R����֑������1?�@��� ��f�3e�̼����4z���/v�h;J7R[j�7\�$̒��j���P��c�C���xw/ k��Q \|�����A���X����_�nl?N{j�c�f=V<f˄m��6V���C���|�k����6��`�* ���6�q��z��$�!��D��*�c���G��=n�I��8yT
�B�(�r�z|��U���O��F�T���Os��L\L�b��Ah�A`�omث=���2["}��#(�L���^�i}�<>Z#��┼�����藹����ձ�d��֘��`��O�+aVMH��t�@ɵ��ܦ:}��8�7&�%�=[���\: �3P<K�R���ۺ�|nx�Ѐ�6�_Z�ư6������Z��E�������$�MkKs#�?z# `���<�*n�%�؉a��J��&����Io�~(/��?~ȯ�h�k�úr9�n�o=?�����}��ڊ�' �#�@N�M��7�,{"z����b%tȢ�����5g�w{�ێ+���B��b=,@�g���rܪ|9�y�D�Z�sϤ��6vN�<�g���JyT"E�Ťj]^���"r��Չ,/>�	i��d��yQs��8���M�T�ZW�x]����� vX��h��z�HM�m+w���
D5���g�1i��'���a��+	#�M��p�-8�W�W�B�0p��)d�w_�I��s/e@���p�R�5���,h�� s�cl��]�5��\���)���Xx]č}w�a�U~��9x�U�����ͱN�
X�/�
\h�`%�w��?�`���SW>.��ܾ�#ɛ��[t�}W6��LJ2�eu�`
q�!��	�lg=�
p'w�� ���l(���U?�7�yl��+e�8r�M�(���}C��a�M�`<���>�R��`t�%�[Y����l^����ϫb~��n��� Ǉ6���~��Q�"��;9�u��2��}d!��!�AĝE�MZ�iK �+D�������ze^6{H:P�W����tc�-U���o|h�Y~s��8r�jv#��'BfD��1��=<~Ř琪?	;�,n�?�N�[7#�b�]�w�5���(*`~*y�$Q�f�`�:���K���d����ՔZ�,@6TY�'dH�e�X��V���[G-:���M�-BTS	O]�6�Z$2�i쨫�5�� ݆L���3������c�����|�c���9[�DI�^V�	vOC<���^ȉ��Lz�a-�4�� ��7F�M#Z�˪i�6�͖�j����-KbZ�4�>�g5��/���
���������40���h��8NcNՃ�4�.B��}�A׃�uVn4v粨J��z�P�*�B����g:a��@�ٮ�k��.yl�.b������6����Z���!��EA f�цW��,I���	��x?��l�1��H�Џws߯�����kڟX�pt���W��C��{�}����)C��ǝe�����2��ZX�G��� ���jմs�Pl(�'�.�k�L�keÏ6�^�vh��ؖi�5�����QQv�p�A���%���о1W.��ǈr�p/�F��/�v�`���($ڂ�	����(ws�&��I�.j�c��p%K�����6ᴿS�?�O�b]�������� ok0f�K�Kb��ֽ[��6�	BMK��M-��x)Xn���I�����T�Kt�2�����0r~�C�Kc`]G�<����e�~.�r�&��H@�z; F9����$���o<��X8@&�u*p�ԯ2ճM)d;93]�k�O�H���aF��iu��bkP��S0�)GeČ͟��zˢ)�7�}�����e(��AL��HF���x�^�K�\�Pe~��H)��=������݌�A)���$�a��@�pk�#���. #֓r��(>D��[��5Y��c�Y���'��եEo�����тc�@	o/��i=��ӡ�\�3�Y����Ը�{��qO����8<��.s3`W�^*FP�o*)��p,�7a�>U8�@�:=� ����9�6�fB�f2���틍Ѩ?\��d����4�r
l@�R�Q	���*��!��&�F�ǹP��z#s����P*�����13C��Q�q}�ݾ�+u�l��a�[�q�i�����^!��` [��g<%�ZN�
�󹜢����v��@��F����+�� _�}���31�d�5�$|���,��س-k��׳0A�c����M���a��J�ݗ���8y�:���f��=� uc��,!k:��~aQ��Tُ��b_�r;�i.�2�|,�F;f�����ݑ�Ǔ�|�T�,�j�������v�hڇ YDt"�=�s�W���A�f�s���l�C��î)�K@��Kl�1i0�n=@��f�)GbD�AT����#P|S
��	��[D��NV�Ӿ��
�z��rZ���uK�D$I�2
p#���Qn�!����w�e�B�����R�O\����=@	�����Ҝ�-�2\��
ӊ��Z�̶�M�A�=a鞢�U�(`�c�n�����w�7���C�_?�4�-����Ԁ�WiT�Ꞻ�С]�7�ŻI�f�6����n�$�]&e��Tsv���xm�4/V����t���2���5�Jg[ɔ��)����������	���!_v�Traz�qx4r�7�T9S6.2J6vi�7�yL���7	����X��ع[ڨ=����B��N�LӜ���d�W�o'J�8��-Ǆ�K��!Ƞ��ZlA�PV����`I���ʒ�HQ�{k#��YYl�a"�Y�t$��bk�f�m��"tإ�
��8c	XA�#6#ɂU��.�!g���K�A�xC@�|L;�Ϡ^�'���hw�b�5�>mm�h�=B>U<�Ӧ	�u�ȞHn����H0XJ1�ț
T��g�� �a�k���<��	��!M�mqp&���&{Yh��_�^���[Ty ���+sQg~�9�4�o�P�v�
�VH��h����N��2��8@�l��[�1ǘ{��c2�t�ҭ �~y�rه��盀�ᛎ'�1]T�K��V��wY�\ilz�{/0|Ud0meNj�!�Urڟ�m��j���g��u�}�q���(Z���K�M�D_r�P�z���MX��a��xg��+3���;�lr1��ܔ��-�+7y�a�r<P#$�rJ����m�d��e�T�ZqY���M�eB��yܒm�n��ྻ:	 5��m���*� r&�zqx�%u�<�]Zoh=��9�����.�ɳ@��hO���\*���0a�1悿�;�Lt}oKC���x���W6w7��y-U���{<AMC��l&�3̿�4���n��d]i
�A��\9X;�J��4:r��F�o��(�]�V���D�&^	/a�%V��U��	�`_C4�ABțؕds���Rw�ҽ��C�|��7P:T����3��2=�;F���a��(��IЛTN�c%�ԯyp���E{VŮt��ۧ�ŷd�m��q�p�T��@lT��S���TO`��+�,���'���j�a��T8(�O`��T�U��"ka���4�^<�-�>TS�X&�x��dR%n���c���T/�o_�L7��L�6�'�i��ѝܐM��ڞ����S���3�S��(�&�wͩՒ4�d��q�Q��3�.��'1|��7��>�㞝�(Ʌ9�ZN0��*BSX�vIÞ][��y��R)5��<��>�1�$*����i^�`_�O0�NNb�L��0�w�|�Y�fB�e��=��q�J��o40�]�d>-��I��s���_�Y���,����}��+��%%*�/y3�zM���Y�o8�I�?:���?���>f�Fx���Un���\[�_��f��*�fe
�= �g��{K��pLΞP��i�}��� �쉋�'�c=_�z'������� 
Ft���g��:�S���g���dĖ&��|�ZI��9r�Nz[*�
�nm�ݹ����QEj����R��+Ԁ�G�Y���S�����O����m�SӃ�*�[sAԊ��jq$� ��yh��#��!��f�;�Џ�%
� -�� �������`Y ܝ���=:c?��>)�F%&�Ř�Һ��]�E��|��;���)�b�.�/�	�m	�I����s6p@B6���MW�GJ
�>fY(K?Ԋ��hq�&�/��o������Ǉ�\�J����u��p�{�p����xڴeO�3"j��+P�7ߚ+�
񖦜������9�����m]�8�b,��r����TX�	�W�#*��Ӑ
���fS�+)� ��I�pW�4��
�p��ꕁ=#�9q(�鎳ٗ�[ڙ�L�EL���?����s;�T}�R�#��H���9��S�d���](T@���7 OL���������ś61x��nwY�u�֪ק1hN"��ڰcu0X�\��3�ͤS��ۧ����c� �zq#��Y�l�ȘE|�nQ��G=B���,�7@0��y��S��MI�g�ܓ@L��`xh� �Ge��[��o���Ǫ�8H����������υӖ@��ܤm�v9[�����w��'��O��/"��������G�.�g�?.�C���T[�È���4��i @B��;�C�
�4ɻ�0����,/�0]�=eJs�=?2������W������S���-x(���LM�Q���#��q ֑�G���_���pj�,�l-�?�8��2V��(��ۼ��I���6���]$ �ϴ���c�=��j�D"Ӣ�ױ���T/��QZH>��י]�V�?��.QE��%���!���`U��:���@�V?�������.�7n<�_cD�#�J�f�H��c�g]�,��9��#��n�{.��9HK1��n�ѷ��݄��D�W㤥��d�'�nQ�����:	�0E^jq�A�V]%�YL%�{u�"���d�sLC�JU4Zٖ�}����R��܁#Q�{��Ф���p���_�N��<���i� ��0��h�;O�$�Ğχ�y�MՍ��g�g�ŕYTK�^�j�t�:qd�{J�P!�j5��+d-�1���*���t��"d�8����)Ѷ.Va�5���4W)�����B�f���-l"�Xׅ��?c�CG� Dr5��\i��aHCT�r_1B,�I�)��D����)�����y�H���\L��К�;�Ӥ>>���x�@R�6�X�a�à7��EX�A���7��_D�ॻ	C1���Fl�iO�%W,s�:$���ڬ���>6�[sV加/��qr5�0iL�/u:�n<k6ckT�}s�����$�s�|Q��x{Ǽ
�[j`$E�&�^���Y"1H3�c9�� @<��h���r�(/pB��;H�q��E��>�
��r�?��4XE��CC�I�����Tg��P
 �gZ�:ei}1�Krv���!`c& �ǰ�F��\�ޠ�q���p�$Ĵa�]�ԹL��(W�r�.Do�zZȅ�#2����q�h��~o<s6I��@����=>s$UA�y�&7�L�r�������.� ~NF�ܯ���,<����D���*�d5��Mf*dm�L6a%�L����� ��л�.'����:tH�`>>u�c���5��]��ELG=훋V�i�8
ޙ⮰��yx����Ka^X ~;���%*&���>��x>v;��2u��x�ft�0�}�xY+O\�J�u���&����NFvr�>��{	n֔����؈����=��.�N6�R��q��׎�܋xØ�1�d ���f�*�qB��M�ٳ�U�hCߛ$�D�D�Z#;�E�E�hqN+�e�-qcD�If�m���ЯBjh[N1u����f�\��тKR��C����s��;B����Q�4��{�X�������]�q5G�oI<����s���H��s�k�Ѣp���$�3������@�"��b���/�v�yѹ�g��J���39YWA���-hnL�P��kq�<n�6�*������BF���'��}v���7\&Re6x�qJ*>�2�!�o�`cE�Jȥ��>���Y��R�fs8D�x-������SZj]�W����y�vմ�^̈́"�I�����D�+��S�ʄa���������!"����_>��97��O.�Ubw:q �xU/��O�5���)�9�)M��09��$h��Fa���z��Ԕ��Q��n�K���l*�C�k�e4�Δҥ������&�-AP�:
���j��1��p{�������vf{4���[�k7�(�UQ��e�I�
	.;���P�
�K���mznD#>�օ�5	ی�m����m_�C�ͅ�p/�1U. �˂��>l�G������jD��[$��;���P�u��5�^�}�N�F��5��������I������l� 8��U~BRU�⮂�&JE�^��lt#��?�@L1
L]Æ#J��C�~lTY�iM���P.�tR|���}x{��t����'�t�|�#�Fu���9�?�����ln˓��^�Hb�ź�y�k�M�\���:�z|Î�׮GT7�t��r*�����s��5&��R�u�q�rYsm�#�`/��;A�/,��n�`�P��
� +�wb���/��0��N	�f�
�1!(�F�w�̑4{��{��E���$�4h�?ai ��P�YT7O�NH�<����INu;� ?���%a�H�f�C����B.�5ws�9\,J���lڰ�PIˊ>;*N�YY�ж��g�'��-.��k�S_�����P����#��ޞ�^?���/H�HZ2�S��'�,�' �ۻ�9�w�P�71;��ƶS�z�-~s����3�ƒ��\�U膯��Z=�U����M�my1(r5��a=",�D�]���u��!�/ѡ�J�;@��o��0���`/��)��YEg�6���`�;��}S�G#�z^$��@��9 vo (V�`ZK�c;38m:jq�j�8��1�V��&:��=��!OP�����e�j������0��������ږ��M%���H�����-)a`dO�����<���za�*qа��'�=�:��˟�Xq��R������^�*uO�|��wV9*�H��$�R�8ZD�-�������z3�%�|=IY|J����['��n��PS��q�g�)x����_;���<��;QG�(Lќ�� ��s�r���)��x,��^�a�|Q�'�^�y�|��0�L��h���>k�h�ЀW�q����G��Q��s�ː����;���O�����lE��]n`���n�,�Ըr9S����E��S8n�1���.a�\������<H�a�FB��HɈ��%w��|F�ƥu�]���x>�S'��%�V���nx�]��*[����o*!�|'�y_"6$��\Ԯ\����Lņ���}]���%~C���Ûc�p��/U���C�$}?������]�~V��<�`�뾂�g�m�F�{�#%v۱OS@�7���\����P;���;xC�D�zK`�jQ���,��_�:�ݠ��)K^lt5OՖB��3�΀A�!�%I+� &r��Ί��̩5�����y�H�0|	��m�<�T�"pK,�g��W�%#�3���ȽIP�����j3I4�{�W^#+����̠}��\�03ƻ�i�ˁ�/Lº����wÀ� {sRnד�ʯ�O���<G~����m��[d����ʥj��6F�.���7̈́�����L;�ȓ�~�
̀���,�j6��,�n�1�~z�!�Z�
:^�}�宐ED�c��<��UD�(6I\�j���*�}�'�:�M,B��Icm^������v�E@�P4���&hj����G��SZ��o���]Km�닜�Tw p���0���5\"���A?&�EP��R��,�zY=����У��lM���$��O���5�%�0�I�<�3ݣ[XI�W�H��-�Hsѫ�����ʲ7�}�V���g=]@���fY����^�n4��1v1�4���z�2��yl��1VO�n6x�WIN}�2!�7��$z5�D�x�=��c΀4,�vP��i�����`{(�I%��d����߽f�Hl��W��&�︹Z�H0�a�)�x�1�J�:5b����#�B�?O������!�������\�@�d�$�\��^�O�������ak������歞j;S`�kȦ�j=�S�I�|�mdʎ���<Dx ���)kZl@r��",���Z�������I~��7E�X�R��G��.J��-�Hȉ�_Zu 3K�!�c��<�C��/�B�}h�ܸB��Μ1%�kamSR�¨����)�"%�O�|%��bV���7a��{�"�'���Hq��X�n�}�H��ͪ��o����X�m:�!�,L]��VP�J}Q�˯#_:u��
M�h��n�
��R2��ڡ�w �Nt�#��:� �I����^>��Vh���0���ꢜ��u
/Zo��l�ܗ���zff��Z�6�
��J,%�H����3>UR	q�\��7�`��x�89!m���7�����6���MOLC��Јu]�S����c�Fvw}eI.p@Q��n�|��᪾;��}�n[Ƙ���7rh��U��=�m�����H�sr�'Zp�����ؖ&U�no$�ܻ���xZ�Ĭ�Ԗac���b��f,�!GŪ}�p����}�B����%N3��#��|~���X`JB���e5�	u��đ���DE�	�E�32�wR���v[�4//���|&�&d�<��AP-��Kb��~լ>�ES��'���QתsIHhD(NtL�2j/`���w��\��*^i��܄X1