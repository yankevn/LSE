��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~3�1:}��Ap*���C]bt�Jb����rg`h O6uf��`�4��0�\��z'�Y\��rC��T�f�X,x�.�	4�j�/�4;�:���_�� �Ĝ�A�F�\8/��ޜ�eK��ր'� ���|N�C%�S\K��x-�כ���fV��"$Y�ځ�����+����C������Uѱ�Y�I>�C���pw��جE���4F]م�r�l5��{��տ+T�"?V;Xw�<ޟɷ��� }C�&��ڇ���Dw�%�����x�]�o�f���iN�"R�%��o�Mdu�P�:�|T��Ε�!��(�����M�_|JL����Z��W����� B��`E!A�/;9.�����Z`��.|��Ɇ}���KC�j�4��J�})8�կ��'F�c���}w�����"Bnz:�y���eP-٥?Q`$ύ���	��A]��(�p�|uʿ��V�B�d��wM 
����z��Z���NS���T������yc�����kU&���d�0�ߡ�-��E��K+���PaHSUߦ&�$���_zA��G[���,��>�c����lϡ{�����y7��M��m%��U��C����������?�(2��bȑ�ǃ�/)��=�'�υd#�!=�Z�o:~�[�@A@�ܟiq��_�w�$�|G�e�R{d�W$��&�m�]c��%�]m[�]��͔2�U�$N~'[��s�è��c�잃=�Q%��&U�6��冭9�'IX<	�P|�TH�	{$S�bLpձ�jOJ�{�G0FU�b$+�@^!#���~)N��4�{��K2�y��o4v 6+G�����0+O���֖�L����T���t�xtvĮa a�/Q0!����VpN�4	��FF�2O�e�Z���E
�29ج�n�[H�	��[�أ�h;�qúe�xfO&�{�x�\���ȵ�C����p ���(�����w�a��A!��<Q��RCf�s�o��w��b$m.�1M�f��@�Θ�ǖq�@���i���%K {�g��ͼ�󈐧	ap�a�.����E�V��L���/N��ew� �ܬ��V��}���K�^��o��,>﫬x�إ1�|e_+:i���C�K�XI�y��>���'�Dcдd�7e6kk׋18�D �	�%�f%��&lCl���������8�kR��z$3�l;��f���9[
�z�JЋ[��A�Z�s�3��G�e� /�a�8�Q��IY�!��1C[��[ɯqE�{S�0&8�;W&�%(�bs��h���o�����9����q�+�63[X��}�fHǠm�J���je�=n���d��ZݥxE�a��W���RΈ�}�#�E�4�ЀY��|U���R���LQ��A4C�nq����~�2�s���9I0&�f��7t�!E�1�
��HV�K%	_Y�wo��Ĭ͈z�A�����m�����	��z�"���
�{��B�<������~~�D�;�Q�(O�@��$����ev�)�jH�KHX1�%6hJE�:����K�;a���v^���|���ǨT)a;V���.{�q���QXpP�݆
H~�����J R�xbR:Re7�g!�v����������<���|��*N��N�X`2qا����<�(�Q�z��sJ��8��,�������m�H�q��h�s[��8�z���2ǚ ac)ln��U�.5+�Z^���(`=��`�D-�J��0¬rQO��D6\�{���edd��U��S�v3�yW2����y�J
�rC8@��D�Nz��{]oZ!�9��� oTx�~m�0�\�@bʃi��k�[�l~/4��9��I�!� ��bx����
�!�=[���Q�);::�s���j��-9��L��<f�f�V����`ݮ��=���M�+�:�mi�9CE#R��h��w6h�U%��[_�5��|S�m���%���a����΃���L��ü�?����gf�xlչ��z��=�N_.�I�];��e��3K��U�������d�%���فk��j�jHA���R0~gH���G1[Lh���hN��Ao��ɑ��wxI�?��'H�W�T��k��̦�<��G�Ci��)=-�F+f[�2�[F�Եg\��y��a�W�
���Yl�a����
��xޜ��qU���Ij�a��lB.b�:��|qF@����%+�Ff�5���Nm�4��Q��҉(�3,jϫ)'�L�7݇���훷1����7Ըq�YE�.�3xR�q�+֥�6.:.�i[�P�HO!W��0ב��y���W#�/�P�S-p��WD�s>�Bgo$��E5_���m��;JN]b���6$�rI����\�V:���r�.���v*A��mRV��%7+h"#V{��n��(9=Z(���;DN�*A��M�&���^��΢\ğ頋y�Fd/޴�/]�.+���� ��fƲ��ۓ�˽aϗ���C˱H����].R�[�ԩ�8��)�0�)�'�-㟉��"��Y������)�Rl$�������Dgk���(�v���(����G�]:|���uF�vG (�5OUQUO�Ł,J���B�/�*�-;0R}�-����f����i%a�&/"��'(���^���=���{,���)�|�<e��!@#z�}1����A��Þ�l�q���p�o?[,	����t@	��(!`..�|�Xɘ��HlT����R(;��+�*_F��QLX(��
�E$��CA4�^��9Sq/7�b�k$}bJsH�N ������mt~�5����Ԫ����تD�!�Q؂؊t��Q �<�� T�F���q��9�]D���:u�[�=�[|Bʰ����K��[��=:�M@�� jM��\�ĸ���70s�V>����Kzۈ�;��})�D���)���v�J�A-I(�����3���;7
�4��m�!�ځѪ@-���V'�aH���jG6:�,l������Vzi�>��߹�W���;e�8rnb#JH��D�10�[�P��|��������wQ�/n¡�S+��k�l��	�J�?��=�E��ҁO�o�;@���p��kOO㗀y�M1rv��v��u�=vj�����e�Hq�R	I���8��+�$���Sƶ1���Jj��	�-�q��KR��lsg�����;�5� �Տa�Ho�]@���T�:�%[�̇J/���3R5�beev��(�O3����#���9�������w�S�q4(�)RW�Υ#����n�鎟@��/��j�~��/U��w6�~�aȁ��DU4�>�9q]5{+T�3A����AQăQ)͢�q�y�=���i����`=�^]+df���p�R`w,uk����+4�r�w��fP9��Z�������b�(�C�s��Z��6.A�>�g� �b7���R���S0^��T�a/d�g��+s�}��E;�S3)ϩ�	��AK��w}�����Iư�f���+��7��⡉�;k��hU��P��������7��O����@Jjiw�c����['ZL��Vo|<�b����	WQz6��3 _μk���u��Ԥ�Qn�z^�$�k�u�P�:Y�NY5k`ː����}��[�,u*�W�P�<�6:���s�ǻ�r���"������lk����O�9jݏ�tA2���q.�_O��bn�e�O#�䇰�[����O���Y�ա7g�D�Xi���q��8km�ɹO�#��	�0�g���G�YŢ�aS3����5S:Ҹ��r�aP��e1ף�ay�	�l��9�IQ�)3i8�$�8�U~�G�P���m�����ݭ>Z�ί��\����!�O���y-CK����;^����6tn��=C  #���Se�a����`���V���US��f�3<av�al�U�Jw��h�!^�����W�Ǫx��k�u�g��H:F�q޻�����mdbtN���np��3�xT�5�>�|l��s�s?OZ,+��K�N��f��lH��uNf�v�_�	x���jy����@�����]v ��������w�x���²T�����z��
�/��~Ř�:!����	Ub�I?�]��h�^ꎽ����nI��T�>��H����V��r�
D+rTk}�ˏד%>��d�D�[KV��kx��V��kZ��^pjX	)J�Al���Ɔ!�p5��P��G��{�2�E9~�H��V�7@�Q�J'��/a��#��e�_-}��!�����b�,��3�}�u8�~	�����h�@~X^��;�j��	s�]�J:"��>4j,]���yd�sX>9<ΊR���n��j�2\�߈�?�_���W:�P��5Ǚ���:?�2�b	� zo��Ԙ�5�cq�Ґ�69S��FT8ˈ��5|�$&X�׬�k�oe�����ۚ��@��H���Դ�1���u�a1���q`L`lTj��K+|vwb	��o�.&\d�-��BF���\}�4	oK�3�ٚ7�~��sz[��0�H��p.\���Gmq����/�>��(������M���/7Mk3n,�L���%�\?��`�KW�.(�8#\�����J��f�d�|�AY��D�y9���2����7�6^�b9��+T�䠫���uh<�|�=˻ �/d��vߍv�K�7@�A��i��W�_f4�H���lk���V�oE�Q��J�o�<{@t!��^<�wr��<��X�.���p"q��T��3����� Ҝ�Y�{b�R,������@S�܀���y4�K�{����ϺĲ�h՛�X�[�$�4�i
���:p�)TӬ��H�����:"��<Dn���0�i��5��o�/�7�=�5�n��r�-�>�Ko1J����ӊu���:䊳��+�`G]�.L��Dc������\�S�ևg�j��k�ڧ�mE%�=�d�˹���њ�w���8{���V�mgY^��L*�9���
�4��+�Ks��k)�?=П>�;V�1t �\X/�!{�`�Q��
"f������	$�/΍�˺̉� �?�;�s�ϰ�Rs���:%���Ћ�F����8��_�%J�h-7�΂��W~xw�[�c��[.��C'0:c�����۩��!7��'��y���B##s�ſ���(һ��.BL�`@Ą�s]�^=K+C>+p�.�\���-��Zz�bN2�	g�Wĭs �(���T����L,����������/ׁA�^t�VY�\w�Q^˗���m��<eI�`	r�P�y��@]f�.}�Vw��@�{�"xs�'C����wZ/�d�.Ӣ��
����r��2����D�Ǘd���ۃ�	t���Q(�"tіCR������qRȸ�^/>��o龊F�;zps��k��V+�{��I��:%\�*�e�~���FB���"D2H�š^���t۲�Y�u�S��=V:��Q"~��f$*�iKG�9�4�B��e3����yAl�-�V�&ׁ�d@ЪR9���<�	A����;��3Ufgy��F���1�9��])*�̖�?*lÝ���T-5�/�O3����ݸ�Vw)vF��0i2Ǩ�bt�?8�7��Q�ژ� ���@ �i�U��[�� W��9B^�S���3��$��ǺnF����@z�Rǎ�+��C������W���L�윝��!�QEX����KSnR�	�*��`��]��s]�����\~��!jE��u
���A�xB��콁�ulV��o�>W�T^|���
Õ!��F=����;�CKӳʊ�k�a;�rA?G��=eV:�}Ki����U��D'��ᛝu͹��_�@�𻆂Z���:Q�$�1���{�\�})�ڃ9�'��|��܁��5ߛ:>7_1�7 #�
A<��;'Lb���_Ҁ�������j��D�ZI�3N5�~�]������$7F�z���Nǀ� H�Im�ka@�v��L7���2�I.���u��l��^�(%��)�K��{J\��;M7h�IG�O�����Mi�a�3������F����ky�*�kyBP��Y=��?�M��ܴǷ��DT\���k���r��酷U�N�����)�4S��Z]�Ҕ��z��!d:ekD�|���<_p�����%�ڴ��9�w��_om�Oj�I�6Ն��6�ο����SF�C�C�`���[퓄�3rH������i�Ē�*S7a}f�ڷ5�x3D���W٦��.�_I����\�\��n�e�.�h���(����[MK��*�V<��n��<�a��
r��I���ש�!7��u�m�sΞ�?�Ŝ�bn$Ў~>��&�u��Sf�̀INu�<{ٲݡN��y��ލ�|c��Cj^�~4�rq��1Pp���	FkT����+g�G�����ǾÉ_ު�!t<vB.l5�;���p�H9��t�����F�n�}٩���=�o⻎x���Ө&�nO{5�Pk�n��p��{㐟�����R�:�u��@�q%����;�*�~���|D[���fJ�=�����.}�1U�Y"�E�w������[iut�C�2���I�S�4%�T�4{j��lZб��ӃZ���C�z�>03�\Z.� �CX��
GI'�����	� �/�7~�#ɺ�<8h��U_ݽq,����ҝ�	Y���I$pH�JZ���N����{#iۍ�4X�ɫ�kL��tP&S��h�17�/h_c�-��u��ƣR�Oo#�^����S[ ھ�Tq���x�|A��k��\Ken=�6���؂#)wƆ�)2��$+��x�����Gv�@O�������;u3�����ɴ���
�:���9���v�#�<(!�ʯ��<w_+��<�0϶07:<���
sq�g�}}�����l��jL��9�V���W����(!���&F�GBz'шA�0@�S��wj�J�M�ן7ơ����M��x𝐪�_��ᘷ�l-���:�7��i����v�_<���a���e&b�>�7�*CY���E��� �7��	��Bi�����*Ȧ,5<�C<%��xs7��	��kVg��X%p�x4	�{õT�,���HOk��5 �bm>? .�$'����h�X�CX��F�DÉ>X�z���l�0��6�xi0/Kuz^7G�)��c�ּۆ~�;�-��΄�o���.g[���j��'�0�|���a�󺢋e��׹c6x�	��&θHߪ��J`�I�a�8j��7�e���Bs<s��ޓ�T�<I8Z����L�NM���^�M�W<�
���R�#�~m��y����;����	�.�w���BH(�F��-<�C�	D�GI��
�D�Iגk]�'4��.{�,��i��I�I|�&��n)+�-�\A�/욛E�BC�Ɂ�Û�u�F�N����g"0��Ŧ��� �&}P�|o"[4`f�� T��f�v��1��,b�����r7�+}���:$V�u��P��\v����t��3]͗+��xw��=`�r���I��UgC������ê�b*\
U+�v�Bj��z�c���4(���/9dc��Gl#d&:tN 5�4�'�j���>}8�R��}�`j~�g�(y©��b�?l��vENE�e��Ɓ��p:58Y����C8dC8�A�mR���lTm����:T>E:p���J�qu.��u�R�q�M���l�O�Kz��FW}P6Ԋl�wWD�PE(!X$��[�Dy�-@�^_�[��#��ٴ���Ӓ��"(�C��S~�	�H�n��B����ǃ@��$C��U9��O욚��X�=��Z��ĕ�?_讀�/��|����n��ޞ�0�ZtxÚẹ���=bč��ԧ��K�S��v�K�����Y�������S�2�_�w��f�~w��B�?��`���}�;�;� @�U�ԅ!���L��q�sZ]�Y�󘈾�z9�A���D�n��o�.v'�_@s��ͲJT����|��7��H�(EȲ�A��$#�����qnσ|�-�|��d�8X1�2�3�h�u�����0�Ol2
�<��
>��������� C(��'�9�2(�b�@`�� ��e�T�������_�}
����W�T7��i�1�!~�������j���랮h�*�v�}(f���G>�J�s-����Ǟ�ք�������C����$4�%<�Δz�R n8�o�y�,��z�o�L�6�O|���&�"�8��:.�x����=�q���3�����L��E5��ƾQ@5�Όw���%�pυw��2�����F��*>ł���Wٗ�����>�4��*FI�)>9ws�*��6��舴�I���l���2`k�~�)�|a���MN]!����-�N<S�%r-l����B&zgR�I5PH���=�k߫vL�%��W[s��'��-]Ɖ��M��'�r���r�j�p��͗�;e���� S�2H,��|�fN��Ve�p���RNb!��r'2m8���!d�R�c?�e6�r�~l-�����5�e����w^�R�˔���G��]�n�gM�M:#jd��B%�����]�Ⓔ�Q�*��Zڣ��AV�}�r��V���/:u�ejƻP0!m��dO]��Pu���r�"�R��{*0��|�4$\����+"̧c���,3�� .b��/�J2<��B8�_l������۵w����>*�kxF��(.Fw/{��f��2������5E/C3I�(��Ή��H���m����ut��4��O�Ya�bd��4_d�Z11�ǌģo�t�/DqB��׷��`T3��<�!IK�����q�M�ij-d�w;g����aD�����q}��"���$}]�S	��6/w!�b��<_z���8+~d�p���
����!��(
�"?���Ɖ�� �%���D��|Ϟ�h�
��7':�U�Ov�������nc���oIy0)��
��4ND��?S�";�p� �����Ǵ=r�S�0�Gx� Q3�k@[֋"$��N�(e@��h�xLw�/����7��[��Su@�N|�[��0L��`}$�i�8�c�]S+K��u_dwim���q��ѐiM����NG�92C"n給�<�		�U��.��o�L�������i��K���ʏ���:i��Cs�9�?M�Z��m�4����L���T�߂��ʙ�,M8A3�x���L.�=T:5����0��t��	Ӗ�P��+����U>��T�;�5��B>D��/�L�^LM�w��/32�e��"@�czϒEM�\K�I\�hevf�5	ƶ�C ��
�� �X7)��YT˰b]� *����d�{�V�|��ء���k ����ة�1Ȋ���,h-@.���7�s���<��k@�2�r��`����f�O0�4C�ؤ��}�q �s[�2���$/�a���!Lf�����0�o���q��a!��t~���VR�_(�f�3�Ƅ�,3���Ѷ�{o�4n��k %�=��J��M<�?�[�n���sL�������\E[=%�`��"��JM$͚�>���t3��q�:y2���.=����8u�W�W���c���X�Ɗ�L3a#�ɻ���5���)��k�n�Es\ϑ�gr	9��R���g��VMG��DGғ�I��u>�N��5ѽ�;�����`=S��'�ف�����@ckm��m�QO��k�����!F���+��+
���tM��/F�@�k�gť�cW�	��w\�t�{X��E�E�]�X)Gs���w�WXE��G�=#��QY���Ηp�m�D���Y�6T��̃�j�W�����.�z���S�y�`[D�>ԕ8�����i̘���g�&��^k� /�׶��\��
�/�{g��JK�02�n�?v��wԽbȬ�SĠ��\^@Ӫ��GK�g|�<˖i96��8f��+:m�� �
�E��N~�Sn�Ŝ{̅l�A����c�k՘�#����J�J�/������8�U`t�TVf�ꝺt�0S��^�@(PU�&n���ٻa�A�M�B�_M�E��8 ��E�,6Į
��ޑ�2�DL�{Nx&{(��������_jZ�ٗ}8�#��H�oL��:�a9p9T���@�Q�Q���8��VRE*ǚ�H���&5�ֳ�-��v1�������>u:�����³E��:Ž��K�h��VV�s&0	hԮ[RL�NպC�GvX��0JU`N�*�6H�1O����N��l!���aP�%�P�A�h�#�A(����VZ	�UY�
��o���^����Wh����eE���M���\H�P�ڵ��dSG殇'{��٧����!N�k]Ǽ<£8�h]TL��_�w�rҷ	�@�� ���Ҵ!�p�P��؞AhQb�׫�Ӝ��E�<�Hٝ��{�@O�|��I��{`$�i�3J����%�
�X�W,�A���u}����o\��(p��^�����g���!�c�!nRJ@W�s=3A������E�X"�f]Q[�Z�{Ƙ���Q���M��Ni��8�t���8K3:ײ:�J����M�d���RP�i5h�[�Ɗ.���?0;UIp��~��Pk���X��s����n�>����Up�ɵh�W��9#[��@U$
��5���ɫ���	5�ݑmu1�؉��a5/Z��8��)HH�Q��܃F��`�A�����9�	�� !�vc~���Oٰ��T�_�.%ע��/�d;�$�a���_�T_���tNF�Ewf ��ΐ���OߟcZ�@� �^��`!��Ä"�:vZ`�8I0��+(�"{��{��c��oO�V�ga��L@�@��Nw��)L|���$Y&�vi�8�9�
Xoy�Ə�#��NAPBߐ }�o|�,R~����L��k6,�2.�qC��H�65GJ�;�4 ��V�s���=N����u��Jl�EJ�pB���F�Ů�}G��6����8�*��I~|6x����1^�e!�d�{=�.Y��F�!6i���ǉB�+
�%\���NÎz�Z���K{Xz2�O���b�d,	���ѩ�Q�!�s�{�|ᜑ��Y�O��i������ژċ{�1�*;���j���_j��7!�D��P�VI[4�*�2X0�9������82�:Śf�܄��E�"Q�S���r,uZ��N�4�
t�������ĺ�F��� �C0�4���kp���5��ņ�¡�|�SraR�$ÿ�
=u��Mϧ�+�4��Nu˙+�o�V��j?�ay��*�[���ݰ�I����dxG�lDo��X�2����N��|z���� ���d��Y"��$����4qB	�k���Of	D�0ǀl�)�	�$��Mn$����V:&�j(�n� [.��v�ļ��.^θE՟�P\��(��.4|��j�|s�v!����Fݺ���N��j3���n��@s伹�zuq�H ��p��b����$�#��Y��5���Z-��E	
^�=���۹ P�%����**j��С����тɌR?󕍸�	c�`��y���6ҭ�1U�8�%�*��{E�JI1�M6Ɩ�,�?�@�8�5�6g�%����+]�m�;�K�������S�"V�6�Ӌ��`cc�xw�Jpt�ٽ��}j�܊2��2mG�������/n^�r�5~Y��q�O$�s樯�r��x
8A`~��y6q��l�:�J���k-ME,��r�����3Cn��
͆��5@�)鵵@�	Pw�g�Qܲ����y���Qv�.�%r�7'��(U&NE�V��C��s}��������J���	eh�ݫZL�ğ���瘿����%�F�fw�W�)ٔ��
O�&��W��;�<����)�P�d�5�nO��/ИQ^���-�0�GI����$��;>�#�D�'��c=���T�Vf����\L�I���޸��k/V�����9�=3��@we��~��=F#ۣ�^u���Υ��C%��V��u�k�Py)��/�MP���V.��'��,V�>4��ԯkܱ��~�x�,!L�N�F%��* ͊���W�I+ĸ�y��)��ۮD�Brh)�c4�[::��Z���g�_���>Q����ٝ�p^���Ŷ�y���S�����Cc%��s���`��0�'G�S�c*Vb�(,��V���QB�N�^tm�c�0�Zm��7��_�N�����^7ݰ�CRb�SlǾ�}������4[8�3 �7Wb8��e�}y���`����\�l��i4qs����!�f���V�Μo|�3�J;�D���b�ݭm�.�d�^>\ldm�$���-�;������ƙ�!0��L������%Ҡ�1f��� Z8��"�E�{m�'4Ֆ��D��b��D'o#l��|v�H��_>u,�n���� �'��1rErOz-BC1�59o�9��O�*��Ԡ+v�T��H�J���b���z:R�
�.��w����9�g��[��h̴c�w���o<�W�`�9�Kc�z�ʱ����$�ݿ8#�l`䊛Z�l~Z�q,0�P 9y��<)�Et4f*]�=�A�
��v舫�+���j<���3v� �ھw��<;���Y�!)g	�ε1�~��e.u�;x֎iR�����*���D���@>{z-@�J�' ~N�`i��;qѸ�s���L{��v�[�S �a�}���p򴥨�>*��~^(��S�l�G;��u