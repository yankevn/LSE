��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘ��$���V�M����q�$Drfl�����2�bP�	��j�YG���-sl��0JL�r�f�I���[��Co��4���8�
�/�dT}9��8�5b�(�Zv�P��Vx�ޜ<dO8���<gT�.�w5o&s�f�Q3��h�A�p�tb�V7�	�8�u
�}�)�Y��XW���y~�����a<T��m��~H���/�B|�1E`��'�m=\���3��\�	�q�������
<��]��P��Y�d��L��k��_�m0-���zB)�ލ~��Y��%�޾���ߨxu͎-�ndO/��P��h�K�R+��sA���ay��d�b �c����򶤴(�RL�a}7
U ������`w�B���;�=����\�y�哃�ܺt�70l(�.�����]���`��&�f�ua��:����\ 1�~��&��ym6֎I�	̰n�7&�&�u���TS�z_�h���@ץ'O��ٴ<�E��p�c��4J�b)�*~���{z(�0�~[��V�tY��7Ąt�0Γ���*胞\�T�����51��%�e�I��@3� L��L *ƬA�@���\�P4Utf8�� \�S&�h�5�z͉�y8�"�F�R��A#�,H�0���~b?���8X����fbE��{��� \0��>l�q��EG2�x#���gBa�,��Єt���X�W�m�F��I>#�5�
d���f>��1�Ѕ��H����`���X��~�d[F�2����mv�������Woq%ǊX'�g��ic��U�/���k�#��e���$m	�G���9H)�M]�(u�c��ǃ�X�U���5'��H�^} R4tI��)A
��s��f*n' �\E*PF��t���e�0���P���La�ø]�U^�l>�_�	��QF��lR�H�1ٮ���zi�ȭ\��TOX�=X2^�IN}''}���4��:eYX�y���s�6H��K��_'��
�y�h~`�,U�䩝s}1r�����-ޢ�كb�*��I�N�lb��h�ˀ/�\���1��Bh/��<EX�9Ь�TuG
���3��r�b��(M�}	<�������.JG2?��uZ'z��	2Bte��+N AE��:�t�'<�Q���Q����]8X��+�~��L;E�^��c�7$de#"�A{2s�v�����d�U}R�!o�1�b�'���<�M�e�՜�����DY��t ;\B�����'<sO[{P;�d��g���7{��p@�~Z�"袡D����V����⾬d�9�3.�[������j�����20������"����z2||	�s�hjy#��qѢ�O��BXL��&"^��PiU\��(��j�+���
�=-�J�,h��ϱp�|��E��Dn��J����Z`V��U��6�3j��F�L����*:��p���&s�/~(u���_W½I;��C���허�O`��Ts}�{�ja����)��i�!��a��*Pߣ�,����y%����©�M���n�w��a��M٘���5#�J����6�$���@py�_r�aJq�$����!B%h�\�鴹��+2�Q�������x�{��=&�],+C>uҁt�ֱr�y(�a��gS}�;	Ji�/�ZkQf�Ys�AF���9�ᙼcIw��p�����ڿ�-C�V����,��j�m���(
���U01�<Zy�S@�S���r|�X]���p^�7�Z�8i��yM���ף��15&��̋q��^�����g>������� �
1Y������>'�
�t;��R��۠x�ep�\�d 7),ě�k'R�-
��{�O0��?��@��
����CJ�(m��S=�� �`���� (��	���'�!V���<m��^N'���Y����"�;D)5��Xi�'��Jj(�Vk��dpr',�e�w+����hb�zl2ni-�و頓i��1�Ѵ����r3Ͼ�@m&TTb�����쓊'Z�X'X5 ?+ao�H�j!Q�xy���uy�gW����y��&�q�F��)�o��D�*~8����ecB �p'�k��x��v��N�<$�`˗Q��b�r;�X(�<���C h1�wh��-@;<=u�yx.'�l.�Ib�!!�*�a�e/T��C$U��yM�Ь�.D[VL����U�J��衝,t<4��̍��,��6 -���-��q �kf��<���o�<�ky>��h�lr6�!�h��\1x�,��Tl?	RY��>��>�����j���z��Z��+����J�/�w/��C��|��f�F�~�H"ܤ��
Җ�׾���^҆u�JD`��f�x`�G�#(qB�k;+�2�~�,�K�{����L�׋,�L(�m�~C�ۈ��kլxS��֋*�]@+��E���ʩV����|"�U?SV���������_�����rz�'�W"�\��'C�3���&�d��:��	�Ev�@b�H!J��@o�eh�ˌ<*ow��jRN���~��v������a�<�fi��5