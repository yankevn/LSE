��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��-P�${Ga�E�n*q$iB��j�ŶAl�NO�p$x��'"R�y��ㆇu��+{� ��/=��663*
�A�3de��L�Wܲ1Ԍ�%)���
$s��M�^;naj��6���G\VW�-�f�ѺD]a�@�K�z=7��lBEO��,K�����V��c�4ێ�rj��.��������HO�#����(���C��C	��2�hl���y)!�P0]��(����y�/�%�8��@1ks���2��ZU�)5����е�cU)4�f��{�E-�S�
���y�M' ��NU	�)\6�nHة�����a|F��>��GOS�9�	U� �,f�|�Ҙ,��Ч�~���^�5��O�vZ[+w�I5���WZ�y�PJ���t˱$�	8d7���2��0m�Áw��b�4�T����&���­�)�"	+Q$h��?��B���2Gat��^ ��jj�Cd�c຾O�	���`����5��/��L%�j�fb�qF���鐍�4�7&�lf(�}���������],�9"�P��fk/���1��U�#���:ć}��O�1=�'}|�<b;��XKy���\�P�
g#Ш
XK���
L6��(J��4�S�S\�L����2	r�g
�S��\k�QY��
Y�c���hۺnD�����ߝ-E%�{����V�����5�6�<2�[��ar�a8��_V�`�swG��?L �@���Ճ����yΐ,|���hu�
nխ9,�۟�*��u=����[,���s��n�P,Q��8v�P�p��rx��$>�$�<̑�7��R'^Hu�F\2L�Ԕ0z;��!��!�l�Ֆ��t��0�M�,K v�*c������V�^�D���|�yд��"���:��[i�;\=�	�ݭ� 8�Th�%»�]`�N[�u����B��!����̹�9��v�����[����-��I��&��:�W>ޯ�N�W�@��a/�lV"��������PR�/�8-w�h���F���W�������,<��t���,	��3D9-���)��ya�!�^N��Q�0��LZ��+q�sP��f�?Y��B�"�D�@�?�d��C�D��[\�T
|1C%%�������:;5w�iE�e ���(ɚV.�|�0ۅ�-͐�T/o����:�s���͉��?�9�<s�4d(6&[ ��I���÷L�i��j>��VU�<_��^��t�l��b���� �� �z g �k��<#�e�P+1�u�ی��x���]+�-����7��@�~_�pL���A�������h`�_�TJ/���u���ͩ!��5��D\J�� ����N�B8��q/��/�w�2ݺ���w���J~��g�k�q}�ݽ|�ag�o#��L�hV�ҁ��mOٍk����NMfz+���)Z�K >��[�A����xn�JW�m�/��������̰�{�j�i�cASNi�����z�#WFM���:U"����^�i~�����?�W��o|��Mi�	�/J��kQo��ϬNSQt���������ASm�YH�u�7�r��j"-�Lע��$u�����)��DAb_]lyw ��J��T-�QM�~�-��{�b0Z�Wr�!#̅�Ű�ԛ29�:S[�2�&C�z)�l���ģ��C�"J#dPb��r�Gmk{�b�l�XE�2j@���;,�pH�&��¿} Ū�p�񘾧w�e���|�ks̢��)�'@<�e��{LG�����(:���!��>�upϩ����ՠ;	�*������'^Hl)3��Ɖ�Ug ��V�ӵ9Ua�¬12��ȪS׭�rTܺ������ VD�� o�(w�aK�U&��F�r��I�b�̷"�U؛�Z�E�r�_���Y�S�D�)�Z�rL���&K�y�CԘ4����I��d��q�p�y����A�2��\O����/��=��^B��������>�E��P�����;���)�-��X�&!��!ψw��˽�h��*����#vX��	"b��
�m�C0�>Z%�ok�ӂ����:�S�������0O�i�v����~HX�.��2��r^n�����RН�A������;��[*�:������VRF�S��4gz�Ξ����Z36%͑�3�S�p�q��`��χ&�4�����2E���'21�!Q3���T��"0�?%�]���	�����t��A�qA����g�ڼ�v{)��LX�� EU�ce�`�Y��=�4��s���� �Jj��%!����y L��rU�{|�zހ���dF�4_hmjM�������̠�ywZ�}�TH�ѣ��`r~.%S����;����%��R5��5J�N��f\\�0w��5#<�m����2~h��EBx[�b�1�<��Sת+	�:0oz0(���*lN�X��_-� �4&���4Q
a�ϔhL�Nq��'�O78̞��H�" כ.�d�"����a��X�Yq܂��� '[W�[�D��Ά>K`k��W�E����	�N���M<b`EL5����}/`z�,���K���<n����p��ć����1�u�	0���9RU�d�����t�����Q����Ψ����)S(�xw��4^/s:�g1\?���:��I�wI�����tceD(k��۵ƿ$��wੁ޼��L�)CCD)�\�$й;� �?���0*�#�V<��w�slB��Bv@��!�`�EX�����<������Q�]�}6w�h���]��x h��oȈ?�@Hח��k��%����d���섐a��Q/p�[���n�G�wV�IQ�q1���mn��0�+csF5�������1܂(��Z���%��|}�����A���#�L;��7�����M�w�@�e�ޚzD����e�9��N�¹,�����o��_�#�E�&f��>Vd蠈ڮ!�a�bl�nw5��7��`�T���`[sq�]"�U��6�FN�����XY�����=����=��TL-!�3�����[*�C��a�
 -cT��Gܘ��F�=�zYi<sm�bi"�b��O��ec��s� :�Б�qi��a*h�xFm^�<��1���5��Œ�$SO��G�Z����n����`9hܝ��n��:�=�8hi{S���֮{Z���o��E?t"��٫)
Ӌ�V���S���ԳQ�h�x��6	��Z�q��n=�x�� ���kJf҃R�� J�UF�H���M���F�n!�5��;��ZX�����)�Ң/o�U�%�V���RFi3���I2r��������g�WJA��@^�̛6���l��\���<o�e�»u�g|��=m����֊%Qd��ߧ�IW�}<�Y�k;�\� (�5��$g�(U�d�m�W�u����0�S�7ȷz��SZ�@5^��>�g@\tT���1���j<+���;�|��2��Vⴻʍ�^���av���X�f���A*_���@ԙߎ+1d���%Z�bYqĎ��m`+�@�L[i%�,��1���(�|���7�N�����������v|�Pɉx�X	+�K�ү��i� @�x��Q����i*������L�{j l=�؊��3u���ȠŇ��d���Ib9��gV���e��j�z��QOy��1J�}B�P�X�#��M�0T_�Bs�E)�l�˫è�;�f3�J$4��ާϚXƩ�{d���I����*��+�.�C��ih��K$
C\WN6�l���Hw�a��o�_�e���%%��X�,�(�,6��%Za^*�I��i�|*�4�K=��jh�9�*GBmR�
��(8ޟ{�X�C����M��U-��kk��oN�䑊̉�u4j�g�}��H�4}�������"��֒�m�!�I�-�R��SJk�q�L:��[bw�`�Q4l!讶¼s�ȹ_�>:yQޝQ�!�!Q���]�����^��_�z����d.ߊ[�!�y���|�A24-���܁����-���Q�T?���-�U9J�;'5��R&huE�<K�kkuxY��o� 8�$ [85���x;č	����J���=�2�dpk��bu=-ϯz��&˳i�À�YX�NQCKZ<����&#h�0T�(�!:*�Wcޫ��	����xCtX����,3nv��b �(GJ�"Qx|# \2��<[p�%�<�Q�
~S�k h�6�M�^�pU$�'�a�83%��8�g(}�8d�����əGD�4�7G�g�0+1���tϖ��m��O�W���d�u�`��-%U���!iQ�"l�PXu`YF�*Ì��y�ߡPĘ�e�B-Z����E]���ON�'J�����%�1�݇"U�Q���x�ӏpV�˙z���&�Gby�-KMvu�@q ���^�r�]�=+z�� �p�	o���.���6�� �Z(5ʁ����䊫�ȝ]�.&��C�Q��J�O�"��I"�k���y@Q%G*'�zy�r�?g�^�����@I?����/8���n$��b�(*
�>�4Zg���eE��a;��"!�4ZN�|o�t~�ݡ;*��(B�}6�G�����p��o	��KG���uE���i������՘�����5�~���Sқ
ؘ��T�T�vDv��۩p�0;�&Q3�S�T�����s'U/�>��ㅱ	~c�wZX��h�O�(���������~�-p�S�}+��-<��&�<�]5�fE��b�϶
r��Tczl;��}�"~���I���k�w�9�����܍�&� �5�{�[���II��IO��d|�$��2�Tc�C�d |�v��I�I�+��]�.J����~s�q���qD�0�Ι)�����yc��9gR^8�l��O ���92`�r�3K��'2�J��G������@;XJ,.�9r4��<��ruѮ�j���S������і����M��]&��Խ�Q���Lõ�Y�|R~V� "�-D�f3
�z��L�	ñ����0� �=d,C?�t��x��x��(��L:�G�L,����z[��g����j��0��ۭ~��,5�1�o�~��2��c�想�|M;�Y�W�e��K`�6����gj�Abq؏&���46�v�T�@�i��l��`�X�χ9p���hR�R X�S�%��55�ym��|Ɗ�Y	w����b�\m�.��	Lp�X�cy�L�fG�L_T�2$�g�.���Sv���H�����vlӵ����C�j���K�X��ղ������81��L�D5�&�N+�"�F�;� F'}�`���VM�++�E6��Q��JH�(�{"d��M��`�(�}a#:6뻐�ϒ~QBN�(C}�A��X�'/�,�hg�y)��'5;d�)2�$�A��?hI�{ۍ��.�ʂh��ډg���z�Ęj�5�9�R{���t���^d|0�RX��S�ML�xMڤ�&��!h{��P��W@Kb��r�M��h������ĭ�G����{rjZ"z=?�"��%);7-���|���,NMz۾_"���!�}�����6��>>�ᩩu㥉S�J�(j���4 ��6�8 ��cX,ؠo�XI��P���u�N>��.�(,���-�RHI��!�9���L
���છiI�Q?���U�k� @���8�͓p�\���=�����dy�P=��ي�mZ��۩ˏ��'�ǧ�UMI��a'Z6�K�
<&�,-�芤��K���ɨ[�$%�0|�^�T�<�e�ۿ8� l%S�PIw~Q��� �DR6����FV�4�ge �>�tWu<�Qg Tn�1�E�t=�P�� d܆T��M���Yo���q���K��,K��<����L>��,#T�(�
��x�tv�@��5? `$�h��S�lk�%̓
�8� LK�H���ݘ:��h_2B��mx���Br%�!�=ޢ2D��W�`~Y!-PL�a�N%��IL�G���ݕ��91J��7p�M��_a�F��K!��ټ��q�#��o^}O��|�D�.�[a�k��ȍ�o˺��.���.�s(��y�BaժC�"7)�a��hߨ���ln�糯T_�4g�A�Z�T��=%
�h��:�L󨩚�xd�b����Sbb?�� ˃a�|V�@�t=`{|��rz�
����T��U[yP�<(�H�Kؠ�׋@V\�q/�h<��.������|(\����
�)z�m��Е\m�K��x�܈�H:��>�vs�<���w�q����M��}�gL���%b�j�K`2��b�S��ģ8_��9s.>m��\�"Q���J�������EW����r#�s��ǆ�5�Z��+IS�S����w�Q��-���z��+�hʍX-����������A�i�ֺ��0�FB�"n����|�S��^R�A��qhfqBt1v����٩�.�"̸��R��<��EK�+��������(eE\uK���iE+�?��-ؘ�X���{�ڣ(�?���8�B�K˿<�uڲv�cL�m0`M���C�Gx�=�u�x���KB�y�Qԕ�^�m��9��!�kϐ����;�:�9� �0I�ی���4/�#�w8�᱅4:���G�ʠ8z]k�J���$�2�K�oʁQ|W�/u!�D�-�(�����M�E��A�b�K��4ә�S�ic�@[�~��� �<���Cf"�§4Q��|+%|f�y��a��H����Z����Y0��������f��Q w��=+vm�v�x�����%N���0�ꟗ3�
5]�������a�誽W4�zKM��7�x�����̧��?�4<�<�Eebk ��O� m*:��['qT��s|�7�ߵU�����^^&�h�w�����
��:� ����x_|�O�b]j����P�3�rb	��󲇑�I�I/Ph��)�Zj���1��$�������se ⁗���^	�P$�(8ET�)��օ	�6o���n��#k4�	d�F����$h���;d��q4Ʋ�]��:z�P�>��oGjbL�[x��8�6_/5�d���u�����b�P�pr�b��+`O)�)�Iz�����e����6�y,�~�U���9㘎`�����Ɂ�?�P������d����o�v`��d�
����6�����`���K$���eQ6V�\O��䩨��q3ї(a�8!2ۼ�Ɗǁ�|to@u��q �2����zJ3�{
+<�`�C&�97Ұ�Q�jx�1w�����R!Mp�ˬ@Rs�l��x���	;n�d�%��ّ�jڣݔJJ��y���������0��ֆqZ����倗��0cR��p����+VU_���]$��p�����S���@(S��>w��=F3_�����t^s��Ε��:���Bve�T.)6�����-��X������NC����*I�o�h��W�clH��ي�W�*/�r�n��=״�`�>I�l���GS�l�Y�g���ӛjj�S$M��A�y��$�aH��1��'z-�>K\�Ȟ��,�*Ee}F4�2��<w������m���ߴ�0/�W����&����&���0�75��V]����Y%�]M:c��y2���7?�Q��%�~���Tz
��Le4m�x�g��Nz�������W"������?S�B�<f�G
3U��]�ֆ��r���[��Vr<�z���I��]�����؍:\��(����d]���,a<���q�-:#���L�<g���\dG����f���������G!��x0�f��b&���/~^�Fy��ֵ���}��r7�+Ԩ����*�E���Nf�~N�[rg��w�	5a :y�#�ھ΂�	p�t����Q	��~��yH��w�)��X:	�";���7�1���geQ��S7�SMY�>�PG�0>�#���# ������׍��8���$���c��J��X��c �^��L��.^�Aɋe�"���;��V�Ԏ�>��@��oƌ;�z�!�Y�+r�5�� ��N���A1j��x�w��h���Uc1�(���HQ��a�̳c����[�������ot�BQ���o��Pj)���+ވ<��e�wQ����j�������Q���Sl�v!��w��]S��4E�'õM�#�aD̪w�{��ȭa�&D8� �8~�V��x{W�^��3I��Z��z�P�P
��F��<�j6���w�qd���T w�-���]�sS9ʙ
I����	�V�Y�=����H��� �Tj�����e�x������⹷Ϩ����cECN���T1ȄD[%�x��-�ۆx�o�
":>|��r7�ӗ�Q;����.�����0�|��"mK�1.�=���~1�~^aa.�'\ϓ��S/�^�O�'���~�n��E��(_|��*��KT�9�|��