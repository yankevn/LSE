��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��� ���/M�R�GTQ?{���`��x�����pw����j��!�Y��ϕѓ=1%������v��_�H�-�u�i��_Ѻ��g��$<u�������~,����Z��(�"��Uxځ�!���2�,ds$�&d��eޜ�<Ǿ�I8u���0�ϩL4����{<����ޅ
�h�
���R5�I~�vTi�MF[�h��6�0�/�](բ�hm"�0���S�?�&6K+WP��4�����@H�8U��$R��Q�cM8�a)��Ssj�Lmj��xx�HZ���;���o�V��à-����1���k��
ў���Q��|�wԪ���Lr-Rg<z7��}�Ö0�h��!V#�if�yi�WT�hy��Yh����4��,��"���KR�6Zi������ϼ��o�lv��GX��R� ���4�{�(i/���YL�5�� ]qv�A%\G�QqP*;��H�[1e��/>��5T�9�`gN�D��7��'�:�	�E��s�p��R2m�N��{�G�����_��Ʃw�x�gԊ�iկ�9�d���Ζi�-� �{J&k)I��I��|%X\_NE�*����4.-�.��z����!XU����(�V�k-��
���)U�XҀ��b�YTŌ�P�'zpk�Y�O�������s�z97��R>|����;���˶0=�Q@u&q�C�O��>U�e1˕ט�[n D�j8�D�#"����8y��6e9F����,8+�R�k�I�X�e���k��x���\�)�R��'��L 3"TB����]s�F����fP�Q���A��~�2鹵����inzК*�Yk��,=�	3I@dL����ǉ������Y��m�]�l�%IZ@�	+�,�y�10��`����5F�%�����X��<8����;7��%(<����@��Y�r��#�������Ko�����[���7"�S�4��G����(�8گj�fna�;U�t���kF�K�C�(s��t�>Շ�˗)x[�je��1"b�E�R��)�p��� ��Ybk�?j�TKt�c�j�Z�3B1=r�8��})���r���1B�dܲ}�(�w���M����/t�L�hSلÊ��&1��\�[m��B��/��%�ߴ����O�aKOm?M4K���i�����(Tzd�j�1�u���S�	^�`�N�W�)�|�7(_���s��5���5z	�;���$�s+gu?"W�:K���~��b��F��z�P�C��FcQ�&��n��'���m��i�W��wU�"��屼Fp+��t;��s}�GV��x�A�$+���x��!e�71�n����RFy��zyc2�^��D^�}��ba���72Q	���(L��)ɨ���3gds�!rp�z����JV��֔:� ���d��Ha���9����[��fϣ�4�0
��R�}@W�яT���Y�y��Dۀ���^$��� Q�S��e�]�,Sꜗ��p��@!��&]�_a*���Av~5��j������u��s��'���B��8WY��*�?Fpb@p�*�KV�&|����/�#5�񢼯����ղ���@��o�>씴�Q_��w�)b2	X�§���)j��/�*t�#��f�Š%�^r�u[*Zf��g5��������,S:C��qZ��U����4�9k4�b��7������f򋔳Divy_ۀ$�,���cw!.e�C�y��U���Ÿ��1%�gw_���Ӏ����}����c/�(��JÕ���I��B4����Y��-zqᾋ�(��;B`
.���/������%Ŗ����3C�^V?QrQ��a4fM.oe���z@�_��*V�؆s~����^�{�J�z2�w`�A&�0R�$��a�0w�o��1;�E�j�Z1��$�5����X�]���)�}*�JS�vw0�]r.Bc�`�M��~���	C��UQ�n��ܶ���"XWk�e�o?��۹�|�k����UW�n���鬣p��nI��?(�A6����r�����*o^�k=w^Zf;R~�ؖ��VP��o+1�}��d��;��oQ��&�G��� �8�tI��O�\ⲷP"X?K�J�tX�������C����vg�q��F�ڨؔ/��FG؝��R��&<P���ݎ)%v��Ks��֦��H����fh��"kI������M�����	Ȗ��.�uXm*WW4놦Uz��g~b�U���S+
W@�t@���mTl����������|��(^ל#Z��Gh��{Ւ������1��$��pl��	J}sG&nˉ��9���:��_��?UMw��F�8�8נ/��I|.�J�GP���X.h��G�,k?�Ud"%8^m�����s�I�Bii!^�j�Ԝ2/�@4��[�~��-@��9�}����c���<R����}�#̟�Eq��Sɮ��v��������dN����SD3���8���`1r&���]��|<հ��d�ʜ�q��C��ޜ�TP�:qa�d��jB��;TEa��2��i�>õ$f����V�V(��UP�(�J�R�!=�{�����SD�K�A����"w7aV c-���n�4���h�"����m!�d�Q��i�J��'M�de������@����Ő��Xp�~d�8�������{tkc�TYF���& �Y.���w?Z�׬C��tbi<5I0X>��6:_*����<��.�)�P̗�PV�`j�%��wz�Zj�QoͶ�Ʈ~��m���f�+7J��툮 �~��]8��F�	�\�%�V��M&,�OHK�p��t7>o��������E�[�;IL�7V��K�S"Ƴ�M�z�P/��%�R''{�����2Qг�.��1bb�gIͲ`O�6�'d�@���ё�a��S���ӐH�F^�~x_r�]ʏ�#T���9���"m�h��W��9���ď�ά�a6p���{����ƺ�R^A�j��,A2������iч�3JNW���ז��>S+b8$T[����EE��4��=���ծd W�Z�X2�N{w��;6[�+n=7����
��rׁ����權��.��!=a`�ڗ&�)9�\���Vd���y��h�l:r��$9��3�00W'����}�j���%��޽�B�ǵ����N�׾�튢e<�@9�ic_����V.�1�oO�U�q]�k���:�]y�����:�	�/������{��5`�	d�����04Y��h��uO�%mXe5vuch�M;D�!���=/�
�������~��p���������������a�*Q��7�	/	I�0�����?	��������+VH�6հ^�r[���E�/�[
�DJK�qJ)y���m�i �����K���nn����f�Z����9�g�3\�Wf�T�E���[�Lp5�]��	���@���]�,0 �#g�x��I�$�Z9��'��O<�B؈9�ed�4�u�F:S�
4��)#�(��O" ��$��ͩ�$�8i����̨k3��s`-%��ak��a�j�/Π�=ױ�Ywz4LS?
XO(G*lַ�֤�&�?��j��1%��G7W���DH���`�]n����@�9�n�jX� Ci�BO�zRř��A��]�1n`�����u�Q���#�q0���5䮒<�ᚪ���
c�V�'7t�;��L��|R;����	`J�;�9��d9p�/ko�V4][��./�e�&�_����w�$�Oο)���=�� �k�%9�1���@�]1+�"�9hw�b�H^�u`d��h]迨���ٽM&��;���V�'/����|�Ɣ�%$�D�iH�� �w�#�ܐ��`ۊA���u�	�������zħ(c��l�U#U��Sf�TWvܖwΠ�y�ӗ��Ίk62�z?�X���]c��Ӷ��r��ec��0�`���<�u����zj�RھX����������G�֢TVd����������$��`K*]� ���垌&�֜��9(?����(@�{z�~���O�5����t���5:�Fc��s�֑�����O5%ZiL��r[�̃�_�w˓%�H�x��K���ӳ ��������7xFk����R�ұ��&�ڞ!��{#ҿ���	��lt0���k��ņ�����CD�����&��&%	�������	� ���H�_��a�x@-d�/� z���p�K�P���u2ٱȋp{��d7��	p�K�go��ړ��q	+W�B4��)�q�/sڷi�������N��ձ�kʕ����#�N���j�+��b��n���g)
��p�mr�C*#۹ ��ջ!�JΆ�}�ӌ���/§(�i�fA��et&R�.�hfg��+	�z�g���M~C��R�B�x6�+�ވ�%��+䄕��S)��GbN�B�\��0S�^̙��jDy���B3lfRO*ۼ�������F�5�m����^���SD�"y)�"��6W�U)���|�^.�[\+8$ ����5b8�矓 ?eX�h��-�~Q?ˀ��/�Ai�o(��]O*��?U�&�������7���G�(ɤ��⺱Y3���dOi�^Mͣ�=�c�T�F��FHJ�*�����:"��p�'����%\yߠ�� ��x�{�/�/6�@g/���ٸ�t+o/�S�S�:�\O��F�����]�^<q9>u�*���6�n�4��8=���5�U ��e��x�H��O�G��i	����^7��v�S�X�U9�'j~���N��˼�~�Q�Ͽ����LD��b-� $flG�H�ֽ35��}�;*����Š:������X*r�/����(.["���zǘ���ѵ�4�~����VyEsف+�fs��\�gT�����l��T��/�����˷2��:q�M������8 Y��Y~����b&��?y}�^;�v�O�<��Y�1��ˎJl
�t 0��w�DÛ��޹o�����o<B��2'�I4�+q��	�[9^�g0��gp�� ���͑W��o4�o(��Jt�w_Vv�t-wNx��{��%鬅d@mQ��
��kn.���W�������}�b������kT��R���֏�.�%�;էe�׮�G��:��杅Yb��2�#��`�v���Ѫ�"��u�r��6>�g��-zd`��
߬�j�9o���ԉc<�/���h��nX(����B�l�#VI��A2PzUz��S�'�F%$��	�� �8�2`j2n7>��mL�izD�{<.�Z	\�1q���� ��O�hݨ��AX�ͅ:�a�<)�`��Sa0���%MH{���"��_�߻Q����I�R�U���1�P��:�*Jb	MO�!*�4�	q[T�|��hmt�sd���>"�y�Z{6c#k�F,�>3���Z̾B?G�T�rH�~`��|���EKP>$"{�Gq3�zϾH�(S!)m0�ݏ� @Wj)s7U�G*D?%$�b�Y�E9r��o��'~G��5�YC���s�ԩJ�z�u�/#わ�Q�ei��h�bysɉ@�!���:��	��e�3)3&~'����C�'�R����P���W�03�F�����|��fV���w�&!P��ȏ��8�J���V�	V�����5lO�`�C�������q�;��Pu����*p�1T���`���oN|������H{����ʂ?���_r��I�(}T誐B
Ý�#��̊"���n�5(�.%�!�Vl$v�x�1n�������HuT~��<`����Ųȹsa�7���E��횻�eiO��������
�0���@þS�������I"o|Hg��w����9��a)H�,�Y8,u��/R�Pi��n��b"Wa��cP6���Z�^�+⋃�a�>�58|�VL�)_b�����!�	sd*6�Z�#�7 ���\Zm��i>n���W��oPJ�|�ǃ�W9>���`�)qO$B�0����2L�=|��(�1%�I�%Й'ɵŗ��z��HRŻ>n��X�0���}g�*)�a��i(���b'��Z��Ժݏm�M-T���Gyޑ!aR���\Ά�ơx~�YN[��B��{���,� ���� _ ���,�����`��D����N�:Q�E�WF�9�����Ho�.����3�������&��=�2�j��az-˝�Y[�>��p�kj��EBQ�A�vH�{�m�#E�존`���+��ҴN���C��M�|��%e�,���/�cCs��L%���ϥ�nc�ԏ+���\=i�`�a�lђfZ�׷��~�Ү��Fv"��ث��ׁ/�R�՛�!�[1��3[�{��&��"�\+��m`�yQBv�_)�,��x�T$�t7M,r���.?	�uAk�9Y��MDMZ�,�8�ݧ�O�ڟ�\%sA�X�\�ǉ)�3>������8w���F��JOu�nC��_����]8;�[�"GD�М;�)�̱'� K��$f�/���-�Ն6�J ���/�r
�2���ҍ`{-j��E�/'s7���i��� ���-���"���s��kD#�h�hy0�jd�W���%��=�CoU�yZ ��<J��R�Q(�TL�rA�����o�Mg��+󐯉fZW#���r^��q�\؞�����gR��,��UQ���wB�I��h���[0��;��C$B�ZA�_=��<sl��k�
��e��<E	����X�T}�kh���b�եT�rw���u�8T���-X���Sl�"�$�[��� �z+�H�bdZ�AUq���v�:Y���
��ڂ��͉6ǝN�8�ç<[�s�����H�����+]V�c�@���%����)���Vʆ6L_����T��zA�1C��b��}�+oY1�	�Q��yRE�\�)��=R��{�1���ˁ�˟Y�7��9�e&sf*��*��n��2�Qg��*�Y���ֻKD�Fiw�;Q�
fv�
�|��W�z%��2N
6'�z�������7 ��ҙ�n��?$�^Q����2�7W�΃�`�:�(عJ�� �W���F�Z!���� �VH�N��bn����t�ӷ�~x(��Z^5�N�~�Q�j9�˧Cd���=b���0���eg<�%�����
��8��v�+��ٙ��W!�<Gl����0���Sl���i0�v�s~�M��c(Ճ��I�3��i+�+%�6Y�Yl�fh���4�<��R���[��~�Ni��'F<�f�)�$Gf�\Aݞ-�K
��;-�#S|��T��NX
j�.�}i�A?A7�l|ɉ�&� ��$f����-+�?�&Z,�Y�[8�e����F�`4p�7��kuܳ�o���k#D80	^�"��!g��*�l5k\Qo��Y姠��ґQQI�,�;��L��rr�\�]ڤ�_!FⰘ�yC�魵Vϔ!q4q.T�Of��^���LH�� �v�)�˥giS�CƘ�������	��H�{X�vP������s��=٩Kg��0M�0p6�����<�/%W�b��_Q� ��
���䤠(�nk���Wq��Q©����q�|��\�ȄHXnu��q�|�ΤM�7���}���ُ����I�[f^.]�(B����m�.�y�Lh�R��P�H�g���	�+E/2T\>����'_iD>�� 	-b�ElHM�9�طY��׺h$��5�[���u ���l[~�m�H04f�fe�T&�vUzԾ��:H�gY�`%x1�a.�O9��X��.l�8��6j�E�-����?2����6:=[FtApq��f���^pҋ�(�h�`X0�S���4"]	}_�h�������,W�h���*�'W�fzW~��=�����K�՟iXgL�H\����o҂�Yt]����kk�������&�g<��]�ݔ�/�	P