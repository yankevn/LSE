��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#�������xڢB�߉�u�=���=t��K?��W
�"dm^ 
�a������^��7�[������^xf}�!�0�U�'#��sǫG�Vꪇ�|\��&��$a֐�m�ЁAHogķ@MzL�ʏ����iM5��N{��M�h�xȈ��1c�'����]����戄V�E���(�b�y �Z[�]�@[_�k�TNI����TC�	�HK;��F��\O�V��>{z���[�1��*�M��x=�ܺ��v�I�~��Yv]��l5�Q��9"��r���R��Q�nB����� �(�r9�ҤN�w�h�t�)����EN�t%�������ި"�2k)�4ٺʺ�����ޒO��iQn��J5�;I�L�P���6�	,1��y��V��覶<
ˌG�ޞ����"#�h��<������p�C�g1u�2�����J�*���gmE�+*`��/d6>��0�.��\8V`�=�5�3ٷ�M�$S`���:�4@���V�>�d �sv��Mч'��r�xb8�Em�*��R�J;c[�bj����}v��EI����8#�SĘ�c������۲��	R�Un/9�ɀ���b���ibz����&�}���d����.ǆtLG�4j�VB������ئP������}α��E9�����?�����=0%��l���-������D*��݁���:�2J����&J�4������͕�����3Ͻ��6�6�z�8{^�.Ea�K�E�m��-�,F��]��R��u�6��P6#��G�lS���Xl�ZV�).C#���2W��#�����̷��,����%�o���d��<�,�F!Ҏ�Fw��	I������� �B�?t�v6�9�=l ����mK5/U����� <]��	���o?!
~�֕o�����%�GW�v�wrK�ӏMM�,���,��U��ȑw���S�E�f�$���F�.�]��}M� y�����N$�Ԏ��h֣{�"�wu������}&���������h��$n�_g�����v&7�ح�O(���(K�I?ߪhy�٨��|H��K �mԳ�Ss݃��J��!r�(��,��>m��q��(+��� �ؔm��/ɹ�Ĵ�bݼ��-�������po�ðFs���Z�g�u�v�;�Ys8��Cx��E��
ݦ��h/%�1$4����į;A*�t�AL\�T[�q0��n�J��f��h%�I�E��k�g^��uZpݕ�eޞ�u.$�Si�fg�R�x���3N���t��1i?#�x�c�j��F�݅"�*�h"����޹�#�IA,�~��Q�T�u�����mW+�zC�=UGP�	Cf���{xˑ��?��M�/y��b���rC^0ŷ>!����岵W��Ʒ��Q��a�+
.����׊�v8/2�~C<�ۑi��ƅ�
��:q6��8���rM�C����U� ��Z�a�I��ܼ�(���,����@Y���D�[HA�ئ�㊟��O��j�C��`�0����$�S���bL��-^���=�k�7�[� �ʇw�j��W�l�u�M_�:����-�Tbm����b2�a-]b0/�Χ����l���;����;�ʣ�*������<$q �Tm=OH��u��:����K�+�u��7��2�b�w��.�������'4ت����|$�ސ�^[˾��ECn�N�l�RSg��W��'"�?ZXCAτlqK�TM�l�%M��4�A�+�d.�NOTj-���No� )7R�H�E)�;��C���r��н��v{�������C;a2i��U^p�[�~�e�Q{'M�P��(Ql!��Ŋ���H2g(<��&��ئ��y3*Q�~�OUX<Ls)�K���q�q��Z���Q��K�4݅��:�Hj���@>���TO�����oa�T�O��L��8�L��vj\Dp<�7��g
���~��g�3�#���,7�@��v�]Ӳ P��Y��*��He�4�O�y<C4���*0qQ��#4w���������x���0<����y,�b�R���{v��x�����.�J?y z�s�hz����c���fŀ�H�4�+�|�w�F���a ��ۭ�����<���N:iY���/M��a�n�2�z�ɚ�D8��G�C��^�[qt�F$�P����hB���o�83�p��$�<���#7Ƌ�����ALz5>A��^I"��0�!@d�nZ:�ާ�ol�ZsV�-���E����lZ#�ng�@�gZ�[��-�K�#g�����j��B���d��]�~��';��L潑z�6�=f�aEWa�Mm�DQ ��,,��
\-Io��,�v��/y~�4��}��Xn�
D�c�p:�b6Z5��,N�Π� ��8��.:ZH9�������"@��&��>EeI��hI�4����fW������-	�Q������4������$đp@p��,3|�� ?���R��e�ݍK�[�T����P��=L; 9h�_��ɕ1��>���S��RN �%p}�!��Ģ'��Y@�ѫ_�d��� �W�4�ъ�{T=l��W(Z�G`/�t����{�L�7�)t�v�|���Ǖ�_Zx�!y�A��"}H���"�4���_+�܌1�l�w<4���M��}������^�V�Z/�%-v1JK�vSn��&UX`�i)����ꗈ�J�{풟��q���g&ė�:�ۃ���θ�*mXw=j=ۛNe����z��k�*�ߝ�u}����?tT$Xʰp�7b}����ٸ�)f4�e*�Eb������n)$����eR��(Q�\!^��]w��##ʸ�~�U4�$�c5�@O%��/��SD�y����,BKSD
�c�5�pJ��B^g|w'��I����TB�ԡ���ݏ0O�o+S���.�-=�Z��"��=˲�T׶Mm�2AL��������_"���Y�)"9!����_->��Ĥ6I)���u�TJ����t��%�T8�F���à�@����q$S̀�
MO����\-b���{,�������_�O�)~�j�$q��RD�7�d5����ձdvT�5��e;��XTA�R��v�9�?5.5)<b�襰�/a�*��cg� EL7Q���`'f.K��͢�h����!�.V�[8�}�������u!9�RЭ�=����6pC�'�_��9�V�\;<r5@Y�@��2�����/�=(8�MF v0���|���E�0�{�M���.������R8�Unf[&�:s�?'Q{ $���T�	��;�a��w&��XH��������̒r�/ɝW�΢���� ��Hgb>��)��,�4��a�"�aҕ�6|1�{wh~��	=CO,;��h��o$R������6�	���Lq�7�]kRQ9<:�L�V6Wn��=�F�eDF��m����V�T�-��Z��B5�R��c.2iR����<�gh:�ޛ�&w�~]����a�wWŭ��C����b�f�G=�	��Gc'<���0��`�GĤ�u�K��IE�_(K��(e	�5nܭ��g	?���-Ia�3ɬn%:�����x�/c�RQa��@�F���b��DD�m�w��Ŋ�<>\�s�;���R��:{�rYE�ڔ_�� ���iW�f�ߗf���S1sE��e����SBã���*�Ҧqg���'EG!����NUu����$����YiH$��:��5��/�d�M
�0�Zo�(�'F�s��sK;z���ڈH�|�� ��5���T3�����P`U�ij������ōG&u��P�)@2F�J�,�M�Ψs��m�dUq��LIɪ?��Xֹ-��.���.Ŕj���MT��m��O��ϲ�@{mL��r�j�,�Y�ƥ\Z�R�i���M�ɤ $��&ƞ/�LT����7r���#6�ݶ [�=��ɗl�r�#q�Ҫ�i���E1<,��wG�x0)�X�9q6t	*1�RL�����������v���L��Ѯ�>�0rZ�""��on�
�BY6�E
���V^�Ӵ�����{Y���N�o⨒��%e��������ߓ3� � yDӝ�$���KH��4٧�i�\�Ja>���'���:�������q�B�����eeQ�� �������W�ּ�c=�cIO�|e3���X6z�ז�mP���BR�A�.SVj�Ɯ�X��5v��,���#���HeAP�?

��DR���b%`?�k���"�Eg?]����2�����޸��y��#%��K�8A��,G�W-��*��錕�6isW���DD��aCF��� 9D�|�x��dp�f��!(ki]>��tE�^b�r?-���V�}c��i�$�RS� w�4�k�,�S�;����n��o���#,���&�<=c$h�M�_�7稻]�:~��2�O����=���|����U�ڣ}x��A��-�q`�A�����*�D[V���ت+�����nG5҅�f�А���Ialև����K{\�l���v�]]M���p��C�{��@�/øOf�S}'c�Qmȝk��&T�z�_ ��W¼p	D�aC ��RN-��	����^�ThF�ݳ���v�Ƒ��ޙ��%+~mqk���Ct�{5�Z�������ی"�@��0Q��Ӧ����J��P�a=c�/Zj�\f�<��R>�-N����WF?���DJ���:�5�!�$�;�f->|,DK%���N�i|
�Ь!�sį����?)�C�q�D�Y	j�	C��tWg�V���rn�����V�=�������m��c<�K�OvtI�L�oI���6[�ޅA"���b�>f�RIB���я��R,�s��j4���ts���&)ug�xB�5?;R]��t잱�"��G��祆&�'���BmV�6=b�����@+E���hpӄeNû��@�ih���,���Lϙ��$������斑"��^�`��]j�j��f@g�|>��/�/I�^�̻7`�A%����j�3�q֠��0��a�Ss1���$�2��<��U�O/��an4{[��B�E�;����ij^Ǫ�&^ۯ��F��:K�A�N!Ї�9U`�*��Ɏ�D��h`�Q�&������(��5�ب�[��_C��-j�f�h1�+���X6�<�X�@�ic�?��sA+���3��?Do�Q��[�..��!gx;4��x�wel������ߘ- kКѤGZ8]5�a�1����"a��Xx�S��7�Y��d2b�)9)'ûP�F�Z��ǅɫw���.SPJ�Q�Y?RC�S���y����!^���g��$H�k�O]�$c�B!����UU�1Rxpu3����b]Y����q��a�A]9�bcQ��A��3�=�A:%����Vv�N���� �a5{V
k}�-�|�� 4�%h�]��]�U��]�\����i�^0�y7�3|��^�H���P;L�Z;�<����x��+�̜���b�ܭ�Ȥ�o֓3z���n}7��!�$��<7*A�\F�*%j�6Q�Vt0晘���.V%�bR���N����[�������ȇ����3�i�6�\����:��I����<�)���2{�d��&��2�uf�=�eM�:�3raHt�\�rE�:���?����,!9kŶ�t&�9ҊB��J����`}tM��=; ��/�|8!��v�SL��ċ���Y�<��o�$����O�ME�n�C/C�-6�[,��KH��-ӳ ���^��RQBc�LP��(6i�V{-��������*&2|��V]AR)K{ʎ>�V¾�& �X���{��!�v��6/z�-�y�-�F��݆+��*@�T�B����D��j�}Z��zVF�Q��^r�� >"�#�,��ωu\�_ILL�rc���a��K8�nVkN}�0�Ȏ�zF��*����U~/�5��c��~ɀ����蜍�E���	Ŕ���=R���1t�ȳ���w�wPmk���iJ4�GV���F'�8��7U�UD�4�}6Z�M���DC�Bpq�e��n�.8����_U�b$�J�y79���q =�B �4n"��؎�$Ŷ(�BRj��2*S���m �	��}��)�;�$1��bO�+���p�����x�6��~��a���շ�nF�^g2Ց%��bGeϿ��Q��1a��W��p�p�X���|6ӛ��Wo��U���7�/u�|MS�@>=A�w&%�a5J�S���L�Imq�C��B*�_�A\űHv�+LX�Vٟ��-�'|�"��\��U1����kͱ_M�Z��+�Ǟ��?�l;p\�&^��rHk�C��)qhW.Ě\C�ow�@�)��Q�������o#��5 �p��b�i����O��<@&�
��7��H7?PD�R�(@V��ɫƹ�i�ǰ����c�_ƄH�Џ0�UX㎋�av2�6}Iѓ���bK%rvJ֢F�����������G��y�lZѮ�a~��0J	w���W�k�|�^�->�e��ap��=������"��4��4��yd��nr�
SW}Q��k�݆5(�a:Wk'6��6}��P��*�9��'��{�5�%�c1��(/��1��j	����s��P�&"��}O�i�	aT��Nǟ>*w3>]��N�4�@9_��n�4C]�8yЅ��n�5��v鑧V�:r�2�锉�Id�4�>_[\�p��'�9x�D4@��QO�q� �?���qU�ߢE%}߃��(ׄ�%n%��t ��8H�̕�@C~>������2۟�x�7�!�l��)a��&{m��E	"/�\n��;�a(��a�K~5��o�j`��6�"�{�<�c�F��o�>0�t��&�1�n�J	ݖ��y�G���aŀG�H��5��L1��ծ>���B��������b;�^�7��;5��u�ԫ��\BZ%#c#�|�����P����_>�-;=d��A>)��Q��Nʠ�U�h-_����e�|����A�󛊢>��Yw�L�����E�����Nq��Cᷗ���@5j�rn?����T�5��"���-��m�I�ψZ��Jg̠�NN	� ���Z'Q*�*��������p�R��h�&�C���m��At�2���JZ�o^oɜ��äU�k;A*	� ԒBy�#��q�����#���	�J�ǔ�	�X1�N��{Br���z����+�M��[L�2m(���}͡p!�*�¶�z1 �^�<̫�d��+n��z^��9*2j�rț`�UU6�1�c��	��G�2S�|A0Y�@�m9�x��f�L^x�0B�c�����> ��8!����ʷ,��>O�KQb�s+���7�؃�Wk�e�6���<c�$�����I�ͼ1����17p��|��OɃ�W��K(���g��-<�@ߖ���򥜆#B����n��]�o]���(vD^v�t c��}��cI��k��Je��7E����j_@�g��K(�1.��nH� ����ՠ@�N��*�t�2I_z��{�!"Y(���`�'�6܍]q�2�����Dnٲ�z��o�e�?f��Ǐ�>v'����������Q:��V��'���xr���*�P�ސC����7�4�"Οh'Hn0Ι�TU�x��r8����\jB�^��5c�H,���r�+�Fhd���ެ.%��dA^�(0�A ���ԗS�o�=�ҝ�CV "�:B�y�:Ϩ`�%.��}\0U��gE{�C%bL�u'^
��m���}�D��\8tɤ"Zv�y����˭\�E*����o��jR��-H�qv&��.���h���\AD��\�3g�﯀��,�6����w�P1D����7��2��af�NGH�t��k!ԍ��/*��n��Ĺu��O��38@T��i�dظz��L�Y;&����R�s�yB��G��o�����Ξ�Fo���,$0