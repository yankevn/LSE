��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�d��Lx����D�~�dE��!oC0���ñ��t��!����ε���}�V���2��˘�8_� �-��Q�r�eH�<1v��b�qj"|	s�z�9�q5�|��,��x��"�Q�z��Ml� �(�EVU���+�Qր��@���K���o
Ԑ�v��y�<	��U�#���Þ��b�,H�ג��R�q�?A$���Y
��-��æ ����i�7p������/%Ŷ�W�Q�Sf���M�'��P���M�@6��]Ddڀ����|�>���r�~m]��o0H�f�&b��	�C�����G�C+��s��]�ߛ�B�Ƒ
8O��wCElO>��:�O:_Ѭ]#�r1�W�M+j"��7��H ��P���!���I��.�5����MT�6@�r\�O�������hJ=EjO�ڼ��?B����J]��oO���E�Dgϕу�!C���$9����}{����_�47�Qҧ���0�,s�+�7:��T�X�u�ӵ�D�֪ W|h �!�k��'�gq)5ɠ�j���($j�nDQ�����܊�N>/7��z�h�Ġ�-���$W
�[�8���H;-�BH3�4��]�B�5�
{�E�:�l��0$"'��jQ��%�O��m���̂����N;|�|���ӯS���J��?�:b\�a��ӳ�,s{|�yU�a0m8R�!	�O�ů߈����9Us_��!�>�_�x!���جǶ�I�T["�p��ӍvSw�&��T;�Ad��ʭ�D�+�'�j�PyN�2j��V�"����ޭ�y�ht�Sa^���h���ʊ;i��� ���H�u8�Hl:s�zW���Њ�e���m��٥Ԏ�hu�o,e��P��t�.�����$���P�r���=��˒�aw�I�XXu}s��P���i�M���=~��[ 4'�b�Ί�iR:��7����Q���&��eI������t/�]n��V�X}X)%���w���S����N���� -3,p�dYd0u<a~+7�H�� ��eI�<��39���u�~�Q{CE2��a��n�um�v�x0Y�u����Y��f�7���RT�]�+���Y�>q��J��z���?	0�y6������~��$Tg��"��;|���>/ ��hn�{���Q ��f![��~�8A�,8o(�u�!1�D�#�6=,W,��X�0�ל��6?%k�|a��!�ƕ��N�E]�3�k)4�FOhiU!��x4A�'��q��}a��B
ع*��c>Z�z�ͲE�Zi�����W�q~�b�y�{mfح'�}���8��8�䦆�X��o����A�۲��?��O��Q6����w!h4��1�t��two�����	.˶7�d�sCH1x�����cZ�p�{���`��:����vܣ-؆� �M�E��9*���x��������9�zn8ɹ��@��=7 ���&��E�u���TX2l�<�â#��Fj����n�!tO�~;X�ݐߡ��*�.���q׽�PQHKZ�K�p�#�I�%L�T�j�+��;~x9j�@�w�⢇�M�^4��xto�Il�עl�'�����ʚ�"I(^��̾&���%w���s�����ȏ�Q�zn+H�J�ת���AS�~���7,k�Y}���!�g��fO~?��/�=|^�M���{��DA�w��
c��̍���R�C�U:���!���\&��*O	Ю��_�y�	�p�[�/+�U�ߋ1�F��n�J�^����KA�6n)���)If��0?���[�]k� L��!�{_g S>��+l�����9�D��o��S���HaТ����%��!���� �V�ސ����)R���N/j�<��s���L�ӹ�s:�VQa��s1����u��M\����0�������Qwlv8��I����Z� O�%Ͱ-���.�TkPQ�X�� ;>"�4״<�R'�!,鱽s(k�_�F!������Y[��s������a��[�Y���/t�6��n�6�ɳk�s����z�3�^:��}o�dOܬ\�V
���1Id]T��'#��&��F)�1o���O�1�>�`n�[銨��Є�@�`��ػ�3���ɂ�q �-$>P1��Hf$y���U�EF��J[?�g�N�H�G~��^Rۃ��I����0���������X@5Դ8�s4�:��щ���ZY*7;��42���T$~?�(����6 n����Qe�[���:%��d���.NWJ<���{&m��'TrV�eu5���X�P �퀐@�.\.�<��/B��/*�9����M��ˤr��{uL~W��{Z�PI��}�8s�a1�l�V8�/F�����j�N�>F�H���+��A�>�CzZ%3X:lS2��iڊ�� f��`â؜�K��y�Λ�q�ȤJ��e�{���iN�r{c�(�ͣWZ7��2%|�` ?>�V
O{W�B�>�fd͊�$k�nP�Q���ew8�@dŤ����XW}��%�Ih��M�Ƨ#]�)�vy--WN��o�qs{�S�x���$�n-�*Js�ߋB)�x�$ ��ʂBo���e���9|�,�fjCBM.��&�jEZ�ˢP�rŠ8�RC����/�N�;�}�(��&R:~+M��ڄ?��|~{�:�4e[�dva���"�a��ի�l
+�����JˤVkL��q�¬�k�����7s>�����gl�N�q�ÁX6��J�l�m&n��%�����JZzv�z�$�͐�?)�JA����s��T�ċJ��ը[R�$��(�٩�4��DK%AT���V��b�q�[���դKEk�°J2��m�[�}{��УBg����ĵ^jg�4#�^�`��a װe��,��H�����x�E�,��Α�|e�n�z�S�am��Z�ݳ��+��w��������ҹ.�Z�hݥ�!g;d7J;��ێ�����}Kv��#������>7�5���U��qE�x��n�3#��6$�wA/4.P�>Qs����zP0�nl��7��$��/"u1���t����ez����-�q{���%"��I}z[��Ie���*�����3���f�a�r�WO��oz[����A���]:�Փ�^z�M�<�&�@4z@���Y"�.}�W9+���<º��m��3,3�6�����1��sy
�b����|���Ž��.Koxڀ��3�X��U�2�Ҁ��e�U��2T��~`j t��JU�-�!��x۸-�����D3Q�p�sn;A�#]õ�j��Բt��~�#͹�E&!aO��^�)gG�iK��a���	C�}8�?��{�V�+����ϲ������,q�E�|�њ`�Ei��C�#��#৲��|���wWD�.�b�zt���@D���َ�������=]m�+��Oº#��yZ�?��tR�J(��Y�F�׬Yܐ��84[���t��l��%i�{��E4٪"�A��X}{g���4KH��������)��!�G �fl`��1[_QӶx3>+�����uE��2��-�j�e�<S��Db�%L��5a�
U��-���Y��a� X#'��v`���{�Y��PP���g�$/1�S��c�������4��y�@M"FI�ӕM�Y� ��>4k��[T���Ap����)�Wy޳��ߚD�|K�d�/0�{��RV�<r�u?0ւ�8Q�m��nVٗ(���XH�W�&�x�H�3�}M�b��@�a|@Oh�O@��o����nDT`5m�#�f�"�������s?\u�u=�c�⹺
�G֝�,Ѳ<��Iw��^�̥�n�0�HE����|��%5��2I��<��C'pja�r��YJ����jt��I2�@(�(��b��B�^-��E�k�OJ�r?��%��5g����� 1ΓĻ�!�!�|�*"#\3���V���`ֈP�>m2C���{��P��I�v�3�p�'z�F����hp��k�ޅ�+|�r�uu�dPU=����0v6W\�Rvg��`���Q����R���(Gz�{#誅B#�s�E��F|!8�W�p���w^����Jޯ������e �(��j��V<�l��bW�5xZ�����	Q�j���_�5d�'S���7���ٗ�M�ߤs�_�����x�AX�
��j��3A`Ǳ��w�pq�a�ӵްv9��(^12~>���4�($U�;,�޸Z�W��8ۛU_m�yRD�4.
Z5����鲯h~�<��R��[\�t]K!#�u`ΙF������9�nA��E����a�e�r���e#q�D��R�,���f�㐐�|�@�P�@w&ȣ�_��VnrߙQw��[PÐ��N��J��ȺBQ� B��E�Ҫ��K���R�<�rs99|ud��Y��2��QcL����r�Fa���~�hI�K��`x�^r#[q�?
�z��)�H�o9J}��\|"�X�����C��F��礮�r}/�ūP)���.GύQ��7�~�A���ك`�6�ss�\$?3��{w�I���T���\��j�����.)[Q�7�&�\��xWϠ����~���^��h�4q4m�p�P\���;�?q�'�3jؕY��g�c5���I�C�c|_���֏�cUx����2�y/3�R�~��ڦ��x���`�ƈ뾎9��%�63�'Ϙǘ���R�^i{�!!-&�4��c˨(`�˦y��6�f(��O
t0��E�*:*����WO��nn��J��7��r�m����	Jಶ%�����]����`{�ɊoF7��f�xK�l:^IS�r�O^��v3���[�%�h̖dݺO�٣|���&�V�pY�UH�m:����(Q	���5��ñ������e���2bkPV ��q&��WT�"�����2a�`7�=V�"+��07'*���e���+�m�՛�-�$Ny��G
��v(�Qv뜶��(dc�cI�)Ќ.��.�a���)$	A��>gk���:���[35�o���a��6o���� ��L�m� XUi�+?Hz���&z���l���ׅJ\�HBe�H?��e�L�(h��:S��'d�P�3��%Ȃ������R�˜L�e�>tvIz��	o��& z��������q��I����4��m;Fp��Fx|�|�Z ��_Z���^i����j6�#=�FE��Q*
���H�4(fx���0�t(^���%�����;�-Qg�.�2�DC�o�����ˠ��G)}h�ͭ*�Ѧ�֪1n-�|��)'��\��yG:��d�[_XK�7� ^e�Z���~-�)֯����z	��إ�R��WR$o2a#�#���0����R�S����ݘ��9D�1 �]�6ߠ���X!�%K/��,�fL�RbbӘ�)�a{|5�q�A1�[��|��l��<qԯ�n�$B�E��cAy��wj0��!��&5MZ{ʖ�0m[øek>K0u�}e����Pr�s���1�5��Jѧ(��G-;�e_dW��La��+w)]�l��p�0�ЙY!�;�0���2���wؐ��|��	V^��EW�}�3���LB��ώ��k�v�U��@�z�^.� �]/���@{�<�!HY�F�O�#��ap>7�h��>�ia�V�5��Y��Id}IP�8��B�e����"�Mrp�V�ưiV�Mk��f�`����l��[V~���w��0��k�|plTmv�r���kr�Gv��q=��/���E����j�<~���>�w�2-[k���A!�k�ۅ9g,2���fU*����/S�����XD@���8�aL��X�v�?�@K�J����ǵ=�UZ���cL������뷟ik0P��@�}G�K��C�T�t�>�.-��&b}�qR�db�����0����P�W�ru0DAEi��6h��zP$�@}s�U���3WM��=�#�`e�g"��XiM��c��<� d�,,��P�A�b֩�#��M˛�@e��΍{_ 8#�z'�JD� �dnm�!����406S�zm.-��W��W�3�o��A{�=�����JE��h{�����b/�|.̭.���.k���FJuji8ǃ��4!��Q~�f'�,u!��� 'ND��D�f�?U� 9lG�����g�:<�k�}�[!������OP$=�+n��N8�E+�[&t|���<����J`�]\e��')�Z3�D�~d�s��e��nYH���#�C�VĒ�!C|z����u�J�DԽˀ
��kK#=��lcV�sI�#"w�@e3�����~Y�0��zH�=��e���i\d�'�^�S�qO��d�Du:��^we�d�������}���V��1'�>�:�r{�h���g��c<�S췚�S�vL�xj<�U����r{��Xe��y$�̍�e���P@Q"q�o^��~QJjB�7���%dc����0wr��s�rx����&�?�%�3oˎ	��A�.4�U�-s�2��aJ)���4��iT�n�n����-�>�I]%�N���{�-`;���j���i�.�M����%c�ی%��c�D�+r���t�1*�e]'84Q-�Ϻ�U�=(���F�	���RnE�������Tu�MD���"7�Y�}I7����A*�Upϩ��Gk�^e\�X`��y�����ei�@�aH���{�RÍ� -��TkftQ���Y곐�0�QAW���I�]Z!pDL%��&��)��P�kyQDˇ�wD��y#��w�3f#���k�g� G +$g��<ښ�ƒ�X�y0�F��VqK�Qh��5�Խ� I�*��>ߩϘ�FV~�W�c؊0K���&�bg� <ΞɃ(o\����Tk|���s��[iv�I ��b���G;X����`Q�P_;D`t�f2�d�A�"�f�r+�r7�Ƣ�xؔ��F���������3�V`�|(�:T�$�t��t#u��B2��!��	ə�`��NXF������;��?vlm ��<�����^<)���D����C�}�4��f�Slo��U'O���q��F��`[*8�p5y�3KRG��%t5�b�w9HB�G�o�=|A���G���IjM�4Ļ��C��F�Q�jqn�~���-^�/��sJ�����oW����*:�����ƃ��"v�ǆ�è�\K�tW�{)-��������
��;�t�U�I�J��V���9�z�k��8�ٽc�X����!H�0:4�����t�d�����(!�QGm��F<_ h�<7�|�-�v�_�2z��7c��a��Uc��߸�1nLJk�@f]����T�i���m�}v3��~R�_xa�s{n�b�zB'D���Ơ�	X���T��D�+�1��;����+˸u�b�%�:�q�B3�E>я�#�}�.Zq��60m��P�u|�B7����k-������@7bm���Qn�p8�o�"��ݼ���F�Q��IH�,۰F8iCNB���v*j��s=[�wr��!מ�%�w�d�O�ڰA�̓�
0��Ӝ� T��Q�/�a���T�c�'�k^�3GQ8t�Y��9�Qw)g�����⣘����5*�M�Ό�W�V/f�!^���9JX�2�Δ��k�'���*�@,j����wz+m�I»�ơL}܋5�o4�E�aٽ9�$�О	��s���^�T�|��ZxmYèҴ�MߐauHW0�ofs��w���+�*��x�`�3�wܸ'��O�;5��N?�Y� "G�f����Y�),\��+X �F�Ď�ƈ~�uH穋?��L����YrI��ۀ�%�f��3�"�B��}x���Es�9Mv�� ����u%�z!j�H7;HY\h}o��} K`����9�־���1?�uq�x�j�'��FqF�#�&|�S�c�'���vp�W�Wj*9Ţ�Aէ�0�G#÷�B�����C9�-5|r�f�,`53�-Ňq�	��{s�*�,�"n�#&���q�Up������*��KR���=@o�hoM� ۆ&��K�h����`���.8���>ſ l�殧�9��x���;�|y,��:@gc�}	��o_4c�O��	�_�� ��Y��
�d{w�#XU��A#[�+�F4��(���K�T/�7�N��\��<�_�a�w�-�I5:�!it.�z  z��j�][�%�[D��_�k��aɞyR��0TX��Y+2��OMo�Dے��-��5*�D�Ujf�s�06��vk��J���&˼��)�0�>�k�$8�`@�P嶲F�����r!��1�����3�D��蒗��/M?Eq���5:%�ƙ6�8��.����xK�Á���������dPLΞ?�����p��D�٫Bȃo��N������۩��W�"���8S��u��H{�Z���_P���a`GJ)�Ȃ�X����{W�IT�V�v��8D�ˤK����@X� g�	�_9F�:��*�L�����0��8J\F���Kt��p�ᷰn�x�E!���Ӽ[$"�XB�r�̱�p#Dd}x ��X�D���23�<h��������p�-�������,=���_:N*�Ϋ2P_�������Uظ����5L��@����ma}&4�<V���:i���:��g5�'���S��A%U���lWi�	�-�ٻ�-�/G73I	�w�Y��l⵻�i!d�2
"/�L~�>������ufo�0�����
��)�����f�˃�Ǻ�fu��=Y��_�ݓ�	%��K�U1v�+�G����;F��c�'z@?~�x���I�!0��[�k��:9�&R���zIYËi&`�:��$�Ѷk�41��������u(k}��"����m�%�� <�g��RJ����d�8��F ����=�0�yH\FߐPP��dau�z
\����>�;����j-Lԍ���=��~a��pD��~ܿ��Ε1�|��N����5�pS7kvo����UD�e���]�1�(ד��i�nM:�.� ��A?������c)��o�B3�������~��|������>�vW욤���p��!���{w�>`����߼V.���;���;���K�DQ�R̴1�3��Ot�8�r����k�7ЌeUQ)��D;�UU�	�u������m	��{_&	����>Vv�^�<�ŋ��9�*�]����@	
��V_�
(�I/��7�;���yc�� 2���(%g@$�;���tM�tg�ψZ�x�m� +f��L�89�^s�A�A��z���T�jq��Ѩi�̑=H�V~��)��j�Q}�q<@^!���f�
;落����C2 �ڸ��������}��#��:�)���n���� �/2�J�5q�����m����)������ƹ�9j ��  �{~���;��(�g���y��z(L��<�u��_=i�mn�U�#/�8��ղaU�aH���d���C�Z^l��ݦkH��m������ʈk��`Ip^�{��Us���.�otU�۰�P���X����=IM�C+���QG�E U��
���	��l+�]S�y�F�������R4�Pv�7�u�>�G�j�����J�wg�����θ�RlWE}9�Z|!1^)Y�7���H�m7(���\i�W2/�,m��	��
1e���
6��x��y�gA> �׷ 2�j��~��A �R�I2>�(�@�P{ʙQ��u�ل[9>�VK�`Q�%^x��
_���L�e���#�Q �?�.\G��I��T?����Q\�oN n-�.+���e?CU��i��t�l*XH����cKpk�{"�2߈7G�R�]g_�e^��u���9B:X^@f�%����y�@���6�1,/��T�O�m�q�7-7]81�f����@�����S�ݛ��@�I,��B���6/�L���*Aw�+�QvSu ]'pª4N�o��`8he%#��B��:�����i���ѧ�O*oπ��)BTJ�7J���r���\O�1R���ѓm���4�t̝D5[�;�:4� M�����L��Rcs�I{eF���h�J:�d�ޝ��<ރ��ڏ
��@���{j	�6��\���JȧI�
��JkYz�mTyn$�������p��g0X�������9�$ �6��\�t8�f�ۂ_�� ��t��즜��oY-5O���	�a=)�7����~��A�ݬ	�J����0H:�2b͋��D��P+��#"�޼��F����_`��h(��hqnu߆+�2��
�=k��/v�<T�{aco�ntn�W��N{��5f����Z�V�3v�H䈤�Q���Be��AR咿��_�]�s
����\V��[�bp��H8���'[���.r��c�ˆe-Yy���=a@�#]�T�N3m�+;����0LO�>���c/�\�f �u��H�� ����U
�]��=yI��-�
�I�x��Hь����_�X�̲����i�տX�i6R�?�N���W����!���Q�!�}�Ws�%�c�����L�a�Z�q����pA��VrK�{S�4�?a�3������e���	J5c]'�N��ҩ��{Gc���(���W�ܭy����@�c6�ʱ"V2�j��ÏsEl@]��D>+��E�L����\W�f���=���8�����RP��zUKf�H\�������$j���:)�t�^�ò�}'W��%C^�"��!�V;�Q=�E�����<�����mE�J��J�M�N������k���{`2�u,�D+����%�+�1��8JM������Dd��G��s����:a�?�d�j�]�Ev*�����pV+�I��������1����N���V������-�%$b[|��4�y�U�jz*F���G�_eUڧ.*�̔L�YP��Ӕ�WS?��mc��T�?f�$�����h�u'k���'�~$E=�̳.HGU�*^��-N�:9�+
��iFyQ�8d� zE!�J҈�� �i��mi�˹��� xF��^�Ͱht�M��xMiÄP}u�0?
��{߹�@���	1�����aF�m����ב�Ĵ8�J���-���-Q�_��ڑ7�(��ᘧ���c�&&)g�O$w��>'����^S��4�u.a��U�&�K)g�k�zP���^�

jUfr�5gެY��>������n�]��S��q��PA�M6�H�D��I�~������Qu,�����?Ұ3"�ē�Ƥ�����E&QDe
���L%�ڒ�c�dDu��K�.�h�T����貸e�R���y�	
��Y�o���ݟh� ��o�H�)�,��LW��&���T9C�Q��B�­�	O�C�	��9o��qѐ^!��J"��[#,�^��W���^�1�P�N��'�T��
���=:��A9�J`�1��G_<�,er��B��d�����2MgnB�߸C��L�?W�JcV!mr�<�y/d���Z��j����M
�[z}��/���_�'�Yޏ��5�Ɯ��ڛ!C�of#7c"�N�"3y�v�����Va��q��3D�d��U�A&8��)r5TT������z��K��s�krw�n��N)y����.--夣�=�3����*
 Fn���嗠�>w==ch1ޑ3W�)�NL���rF����F( �nk��,鐮���!�W�;bt*���vzZ�J �\�[�S�RS�RB��Y�>�j���'M9(Y���ѡ�.�ǘ�(ޚ֨��sL�rU�|Δ�̷'����s�G����o@C�R���E6nTd,a��0t3�^c�p�+�~<�����?cf\��ڕ���p���8��g�?蜅�ad׺.��7K��0�u�S$��H�
>��A�&�Fwz���Vm�jD��m�Z�D�����0��\_���^Ԫ��=;��A$�)��}y�{\sR�w1�������\j夦cG�+&�r�r_:?��V�Z�	�����B`|�PPf�ĕ��	/�Bu��k�@]lz��Qч,�d0\h��8���;��������ҩu�Z���c�=���J����^��վtb/|���R|?����L� ��D�4�1�^1������U��r��s���`D�[�%���J!@�]8�7��C�ћ�j�"@�s��H�s�+C��ѫ0��]���{p޴��G&2xeͣ�!�^�>&�IAX�Z���鐛�e��SJ�΍z$��s��	?��؄
�<# ���wK����vfވ�Sag��99������p�Z7�Ұ�s���v�Qe4b��pvi#/ �&� �1f�����
��X�O�`��F�,I��w�?��fu�17+X@�7�x�Uֿ���x�퇰Fk*g�.��_�����
��a}0O(/iN��x]rX��ao�)�V~���T[\�ߗ���"��hLp3��7n���o����J��4,�+A4�X���N���DKH��(q{H�Z~�9���q��y��y�KFR7\�Oݹ�m9�魑6�P|C��}0.YcP/!��5���N3���Z_x�sՋ��LD���<"�cK,PZz���gS8���,�.���2ԂD�]��`��@(l���RJ�qɦ ������l��ݧ��ڏ�KYX��9.��]�4Ex�$:�q�1�8K��<�2Sx`���b2�̆z:n�0�'X������fL���/�Bڣ�Xo��E�0~���~dڤ�\n�5�Ԍ�l�ܠ6��	���_%jy��BFJ�hXM�A�>��CRf;��^�=LP��5)�IX���Z�����(�y��n���������>�k3�gj�+7�B�T������f�f��A)M�,�b�.���8#8�n`)�ׁ�q��n&���^�7���w��*I{Tؿxx�-�0�@��ϖ|��.Ol�b��V���
�K�}�o&L�n,�� b�[zzrTԎo^*&/M��i���V��I#���mUD,4��y�m|گ�T8������N�S�߭hb����"�7���-�5A�Z�l9`
	}>(@�a,荺��a���M���o�Γ�Rb��F�o3���Ӆ� ��	�����'އ��C��X�q��J��q����V�v����M�	�V�ӛ���q�|�����%L*?_]��q���Ɋ>'9_i��$����)��c�3L	��Ă����2�>=['}?�d}XE��t�Х���gƒ�֩#D�i��AY ���)���t��+*��������kPe�.OQ-Q��*7%x	�o�IҖw�,['L�o�����$ɩ����c����o�I*f!��ބL'�~�fH��x��3m�r>����aݚzΡ�/�,��np_3�,�6�4��̖�'b$�u�R���yƔ�ϖ�~	T��!N��%nͲj+��:{����"��_Nٱ� �< zu��GQZ��|�=��:�7p�>l���aO<�,��t���P��<
���Ò_�I���+{����@aTF�+/���I"4�0��YSa�3��y�;�xX ?�6��&�nL�I$��l��F�n5��_@¡�ɢ���P�-c�&G�#E�����ƺ..��3����!��t�{��}z	�4~�@c-O@h[��?=��*ݡ/�SŌ����?VZ�gĄZ�P��Y��#~	�u��n��p�� ���|�'�c;YS4Pܦz7�Q1�x��[�����<���@�/p,��֮����u��LM_&X-���ȹ�333��	wnl�KKJ�o�$3�c�?��u���ς����,q��!Fk�v�6�� pڒO�h�V�^}���	\�)�"���zU�;R:��t��U�c׻�7O3>=_dl��V�A_(;LI�rGt�V���+�n�\�i���-�#x��)���(Yi{�)�[�FD�0[Y�k�y�,T-�习yԟ�%�*���P�<g�h���Fd<�<�D0�l������d`�8�G� l Vu|�0jT�]��\g��S�ޛߘ����e@C��[@�)�i��6��Bj�MAs��94}Z0�w��O�##A�2�|�=oaD>I�+<��2E����
�nS��4#�y�Ʒ�Пkl^����d�M�͡I�+���l����X��Q�4LSnK�#�`~['��T����@F�� `��䇷,�_�y�R`��Qo[>���{E��Q�f"��� z����fH�'>�HD8�(����>��@Oe��dNH�Nq�|`�z9�X�w������ZF0c�����3�_[��4Ys����!�1����'d��v�F��}�(�<��OXO�.��.$��=�>�y��-�>��Ϫ��>�|��dz�?.������qE���\�Q`��`>:���x��S�=�f�I�S=�W6��郻����H2�%�>j���% �!�E�H���w�7�%��d���k��r�W�� ̄�/\��X�b~p,���jZ�qL��W�ɵi�i��=9&>�x3�+K){���{��7 �EmAhٶ��"p�&��7�i3��:�*y�dBʪ��|��Z��/��PW�`�5]�4��Y����O�n���Rry�u�0KM!4Y��S�g��t�󿁳�gY�IC�"��|�p��"�8=��B�f��/�)����~��Rw��������TH.�P����o���\ݵ�����b�"��� ԠB�9�:��1>T���`J}E��q���V�%=@ЀX2��U(��RDΝ�xc58�� �l���1\l�i���$�aեDl��w�*n	?������u�Cn�0\��~��H�ù�nM"�b�=,\F�G,}��Î�x��g�0M�(�7q�(��[fZ>!�SЁ� |�ih �k�E�|1F�4�1,���)�`�C-����L~�9�e��xX=��g�8D}��>T����t�B��	;�B0�Y}���Xq0�ˬ&��g� -�P�Qx.��wq@G��0���ސ;�=�NV(�a���2U���%~[����D��U�{�~�neL�J���~,��iw�f�����~�~\����L3q��yũ��!=��9��Z��g]N��M�9N"+]�*��D�/cF��ϡ���G��)���r]J�1w�@���WS������U���<�M/I���f�3MjP�d���8�t2�#����umf}lʣ�$����JU��]������|�mI�U_�	6%=>;�W$y�=��Ra��p9��)w �h�[�b�-7m��0�A\ ī�]�F~�,j��,�`ܺڇ	 9.���f�R~�$@��AC�<Z��ÒG��teNĹ9����(���;"��'F���+��4U<��E��ݕ��,�U��~��ΔȲ���M��_�Å���Eg:��n[e!xZ��Ͱ��=��@ �{��}bRNc��b4��j���{�Ǉ阢�4�
xm?�HA^е����j?<�
���0���Jrz�����ư�:�Zyvn�����U( �&,��_�v�{^zt6U#<7�8*]��r��ǘ�9�ڹ�D�h��\���c���һ�5
��g�?lx9v�]4f�/-\�8m�������<��cJ!Ɯ8�V,���5�&��h����Y�^����=�T�����R�
�_,�
�v'��X`�p��C��(���n����������Z	�;w�����uU�]8�A���/
��bp)1�e�.X��+��H�����%�X�;��A������$�Jf�3�&�'�4O��
8�r�\P��I<�$���U��=�DHb�o��u�o1�3��Op?m��@+��N�!SJ���,,"W���Z�̐�#E�`i=t��E������k%S	|t�"+�G*��k����f�Ȅ�l�9bD���8#��ê�vwJ!eϬ\;Y[�
�m������ȯ'��$4���%2!�u�R��1�Q�**bp|���X��<||8���xXc���vO�"��e�c� ��Ż���xvE���[����u�^����s���-�$��b�cP�iN]�J�TLO+ފ�Eփ���,p��e�!7�}�EU�8r���-q0uy���$):!]��Q��{�#����M �X��\��𸄘�{iLIK�w���~��E;�1����5��3�	�M�k���3��Un�W|���&u��ȱ"T|�o�QEU��N�z��A=�5)�RJy��`5����j)+�
��$j��tH�=Pǎ*
�Ç K��Lm{��n�/Cw���	����qPdH?`��%���v��8�r�9�PyZ���s� ����w,��%�-j#~7���2N��m�Ô7�=�"���aZ�F�)�4��>��	U�-��7������|�y�g�t�ϯn�F�������	����-&ǻb'��u��Р�C&1` �n���J�o��m�v��k,�O��y�Z8��y���څ]��kq�
���y���<�Į���K_���έ�M��7w���,��0�fE���xi�,���Uä�
��|>�>"F,�5�u���ٿ]o.��˺��^�W.HBQ��^B�J����!���Z̈́�rO�R�.��2���ؙ��L(Y��\SaMe��L/�l��>�>��
�3���֨՛�� ��IޤfY��'��k7;!�4�u�ky��lȻ%��T-Y덭Σp�ò�B�����A4$fi~�f��K�@a��x/W�Ui}�X� ��!,�a����2c�@y�"��Cx��o�6]��WT?�R��!�sh!_czO�����1��#fQv��S�<���&��S���fK�J�2���;@�M5�M����n�	U߶��1+|n�E�GeZ^�����-'��*;^�.c�D���"�[Ս�6(boz$�_��G
��� 0'�K)!�L�q3��'���m��0�{��=��ö��]�Hc!E#�iZR�/�G;���P ��"܏�u9�C������"�� ��*f\
�h ���Fd�nڨVձ��������X��T�/�5�V�y��~�>)�ͷ0�O`�T�]�I=I��]��sB��ax�oSs����$<cv��?<0��?ʾ]�91���n��g��o-:��k�@�2~��slM�:Ԕ�2�ͺ`[�8��U�iaΓIY��y��j*S?�iv�0�4j�qg����]�D��9�n
9ĝV��5������_�ɗ'tH����a��L�"���G3�����Sɱ�Z�](t��S��d����%z�Wd��09g�|�h4Z�>_5H�C����úP?&�r<��̣�!��v�a�	 ɟ&/*� h��&�a����a�8x���!��>����Kd�MI�(��$]�����r��#9����4��}�������^�=/75W�����9_j��{5������C���XE�n,��t.�jL�x�g�E�ƑF<��q�\�v����K"(�s�!k*m��>�L5����պ����p<���a����҇W�;ܭ����p!��tf)+Ҟ˰�ɀN!�cZ%�Ď�;��îx\�<�+똝�
����*ɦ�[�,p:M`���X�eC���Wp?�J���0}|u؏��͸�7�f+a6��h>����?�tA!��ΰ�=J#�w��ь	�P��t��ڼE�࿵R����ui��*���ԟ+��_i�����13�<ީ��*��V�&��T�@��^@���y�m:~CÕ�溲oz�/�%����/=�B�!.-���<��-X+dm�N�xZ��v�q�~#����*?�(����ʾl�!2T)���Y7e�z�Dk5��7�Jo�H�8eAC���7�i��^�4Y�,j�A$53w�s�޼��77UE�g��ҺU��N<��X���<���0��Z8Z%�D;%�AuQh�k{���Z��X�V�=�HI���N� ���#O�S9�:Z�����*[	�̼-�6�1!��Zg3�8f̌����4r�dj�9�HSP:�o�f�j�l���y��n��
�%��Q�:�U��.����m*uHȑoռ^o$`���8d�EQ0��&�&�X�6�fZ)�q�y�т��qRO��55j���n�� $�*Z,�F�_:���r�a�.o/��./_��7w�VL�1g����o/X����g���=��OZ��A[&JG��hj�iZm|`��[& !��j翩�M��(x������1(;�P�4��%#%M�$�9L�ݨ�Ы�ۊ��?��ʲ�,U�`���ؐH��A]��gK��*�d�n����kLޗg��d�7E�ļHԕ�wu��b[�S������5!/g�{e�B�ͭؖu08�?�A
�6eM#�����kT���@L�T8*C��1Z�������m�3_�CG P3CAp��5x��&��
5�����z���̮�t��yd|	Y%}���7]�tn�h����Qu��{�����&=�89@��B�V�?~���u7������ͣ�k�����ɨa�܁Tx��KӝxOG�6@�B�qyH������ºa�+<�x��*�''J��_�TUN�L���sƤ:��n �|��L���P�sjF<��s����Jn����["�C0���[�~`��!C�g�E�_�cm Yg��62
�[�xp
D[�t��v����E4�.>cy8�i�ab{*JEش�8������[!y�t���(C�6`Fr�掜{��t>�`�Y%����N�?F��[�L����j�w�/\�]�`/�܁��\<j�d5ı?�,�ϱd-��un����QD�Ɔ~���M�3�T�����>�!��}���r�D����0	�l)�F��}j,��{q��퀍��O�mD8ů�br�	2��8B^��7]��\f\��2Ax�0#�+�r�ƴ�6$��3� |�)����c�n�cp�mЩ&Ɯ���-t�.����|	�`��!�o׾�lxV��)Op��bʽ����-љ[��%;��1�� ��#����W��Dk�O!���E׮�v��n�2����i�ư�G��]9��q�'a�,�����vs:��N�M�T/"<�����/���I{#1I(\8�N��O,���X�g� ��g�����3��f`!���
U��';�����Ph�sŏ� � N��A��=b
��`�����������3�Ȧ�^�;��P�64�����|���9[�g���$L��g1&6��f��'�8k
�3U9���Z��N4��M
�q���3b&dm��̾�'�%��Z�lf�gʞ��y���a1�L^:4���a,;0{��$T>kO~�jĠ6��g�����l�6��c���E�1��f7l�wZ����UAm�#�$NUp�4I:7#[Y��ʄyҡ!*�4I,[�{�Gl'�&�GV��WǊD2���4	Ź' /�Aүt���ʬ�B<��u��O_8���<�H�w����� �-l�8W��LM�	SvɃaIZ�娷B���Y�zca��(f��'u�g��	J�W�<n|O%�iN�4����lH9�:�i�ݣ�k��4�X�i�34�7(I,H"�_�?�CA�w��]���� �ikb�k��,�=��.����6\}�0}-����|�l���B���Wٔ�)=���D�zp�*�Մ���$������f�"���u�n�y&�F��O`<�}��F-�<��_�]yGnL�4���r���|���8Cec�7�ŧ�qB_�.��Re�'�O��1�����;~�t�c���A|�eo}��U'._/-q>���)�=_���r�Ġ���Aߜ��sJ��&q�g�a]�̗��=S��(�ʆpH���c�q'��9�K�z�����1AY��3I+��M�����TX�fa4�����(e[]�	�r>y�F��lp�~C�;)����s��_u��O��M�;�o�B�K�+�-���<��T9*�Z>��2T$�ߥo�ZOޟ�;�l<-�e@�8�Ӹ03�2js_�
b�������Ɣ�Wu�9mMI��\�����(漃!�]٨zLTA�E��|!����(�yl���?嚿�R?x��)*����U3?}�M�r�d�8�2˱��&CgH:KU�PC��U���G��PK�T��U<��4��f�{�����]?$���d�Ebֿ�3��'M?�W,r���S�x|��b�Kw�uL��kXn�r�^x���~�#����6<o�P��խ0qb`I�� Of������"��ӁP=��I�0�ύy[�Ά�;�d���m�_3����֤7ïQ5z�U�8�un�1<Fo���L�7b��%ϒ�9�{*3��4O�� ٥���.i�U�:Ǎ��
��x���RŻ1�<H$TK�},jW'�%�&n��c [����^nji_�R�Yӎ}%�s�'��Z��D���G����)�����ipR�2��Sl����N^�L��`�`1r��ֆc�:����.R_a']���A�5�o���i���R|�!Sx�D�� h�q��d���мWV�d�[@ئ+�O��
��Vܺ�UG	��&lRW�ߠ(���ǯ|�ob}{���br�����S5وel ��R*�k���e�uG;V�������I���ƘE f�On���ռ1���w�4޽L�3����`a}�$tW����S�yx��L�.�H���r�5�xi'o��>Ţ}�|��''k>$��H�4�m�!8��!o�r����z0Ȁ����ǻj��S�lM�Х*.� -z����X �Dx�~? ̍j��b��d� ���%�_�t���$7sW�Q�Q����\�m,��CoO
P B���Z�~[�r�ѻ��d�؂g5�Ve���f�9z�0�\�e�U�V`�����u ?54k@7��� �����!87��]YGJ����)�.�P�iV��G�B'�CO��m��ѣ9l�@x�s��AuW_%�Mscz��Ɣ�]��-�[��i��L�I:O.Yusf&Z���y��d��N�0-��$�Ѽ�	ˢg��>�!�B�]�}b�Jk���߭����>y��݀�-KV�`��UV-��p�R�����`E��-@G�ӣy��.�"lx����[���?Eb�Th�BR���d�!I����<�6@��ϲV�e�|�'\≩F�UqҬ󛗇�&f7[�q	�\��|�-��wt�3SQ�h�s��ys8�����J��5jg��}]�i�t7�D�6��AJπ��E��_&�+�[p�*�eà�,v}"ѹ���j�g�{���#X�!����dߕ�K!��e�7D�`S�0����p����C�t��u�_@���z�l9p�y���W��(R�a�O�A��� G[$�
A��<�F�\5mpw�y�����`a�b���l>�x��R��U��x��ԡ%[�Pm�͞��ͯ���F�P��Zq�d�1Ih.C�Q��;[ �찼i��Ⱦ>�n�8��a.��6iTDL�d��(�ߙ�]�Q���fW���Q���+�I�5�ڇP�$Ȣ^zP{�u���(8����y�{mF�E�mH�N|�����%�=�Q+���5�@�k����{�	l��a�.��Ҡ/��5���:Az�Q�V刧���&�b�$~�����5�a���ˬ�K&4�6_�߅���}DE(~�_>��w���]�<��� 	څ/�U�C�Am�&�IJ�;�,�5m�_P���z�Z#02� ��`Ƥ��I����[mW�Bbp�T 9�͔��
���?���{�9���Gŭ�����gu&����S�&,$���-�Yu9/C���r+Z�Vx�l�zq�{&�{rhdq�����Ƣ����[#�#�I��Ew�66Ό�c���Ĥ�;�1o�y'f�!�u����]3A�G5Լ�
���C?�������r�Ǜ�����F1�<�O�~���5�K�[.� ��^��5��q_��2�2s8!����5o]�ךHQ�n��&�ch�^�6o�N��87xІ#p�=��m���I�=)h}x%Da�I<���W��(�Q�Ew-���Vԙ7L�,��c��8��>FZ���=��`����������9����3K�Τ�}��{X-��d�e��$t���=���i�| ������I��R��"�B��'^7t���
��}S��s�l��4&ـF�R/�[���L���ΠDT� DK�zR%<������/��v�Gж�h����4#;�J[����&Sn�[��~ސ��D*�h�A��5G�.tkG9��ɇ9��7�8��c�R��3�,j��@�~���!i��z���;�E�vIg����#��=���*k�Tp��:���CJ�뷄�)!��S�A�v����ԋW�����9^��-ڎբ",�3�aa�n� 9tY��>�2xܐ���pm����
R�N�@J�<��C��!�`R��@}�o�����^�ΝQ�����:�����Cs��;%ԛ"��%�=��@�L�\�f�����+��n
i���o���\�Aױ�"q���Q8�m0�C�ODS����Oa*q@��eS�<�x�	�f���c�ڣ�d�(��}0���jA�^)�n#���0��N1sڦͨp=�D����ŗe���ڀK6�h�+d��r��g�"�Ñ�+s;"�KD&lB�^~މPrQ�o��Q@)`�h�w^+Ă�EMFÄ0���m|�g�1<�����]�m5����u��H���#}ݦ#0����i���>6��&�㡫u���R��@�? EޤJ�W-|�TBUxc�+��=z��E/��#g����*�D�^�G���q|�(6 �R�g���U-ܨw𧫀�6��=h�V� �����2U7(q��@�JS��Ϛzo
d0!=���x���rQ���܅�i���9���O���v>�3L)l�1������n�&O���g��qO�����#��xК^\9�S�MhO#�W�d`��NR���^���Y�$lf��L�I��ZX��U"��s�;4�÷ڣ��HY�1����Z�w�;�i���S<�0�䮏iF����W7���K �/k�E��po���ҺT��k)/,9a���\.�,�.?��������|7�SH�E���`�Р��xq���k^�\6ZU��ѥHw�_�g��=��t�L �,�@�dǂ�#@��嫫�@�r�Y:�)p�P�R��V�"�Bd��o��D\��\�z��jY 43#�z����ß�Ջ���yUn�#���u�{v�)�rDS�6�<W���i�LlQ��b/�j�Ʌ3��E�0Z��ht�*)�M�
LX�	����e��