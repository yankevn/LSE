��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����x�j��ӛ@�G�C{ �`�*��k�Y�u�oM_�#�,���ֵ(v���?���!��ˌlo��V��٧���7Slh�݀32�)X�"�#Ţ�� ��͢ڵ�z�Ґo���	d� ?�ШS`60�3���6�_�F�L׻���1��� K3�mQ̴{����&抓%b?8E:���N��0w-��	�BF HP���1�p�@�.>�6͙�K��(;�@���/�C{_���ڴ<!j��O�p8��%'K�<��k��N ��h����>�<�` �s��p��P�r�P.��I���,f@	#m� �U���r�b�g�I��R���2r��U����1�y��@����?��[�ב�@��Lw��Q�qJbOm�[Un���D�oW�rr[;2�4<z/e�Z,9,2c���ۂ��`ˆ��-��[b?��U���e���]�U,�̙�KL��=3�d���W)��y|r1DN��-^ >7���)m���0��ޢ����T��Z������+�񎺀c��bj]b����Vz������Ɩ����f��v��ۃ�;/[f�{'FVu�lE���RB��|��&X�|Ka 4D,ɨ��MDx����T*�K[Q�@��P}��]�K���
��Ue�S�ex��ɹ�J���)OE�6M���&S����R��k�l�O��"z(�l0�ƃ�Wqe~��ʛ�amhi�ˌ��Bmnw�x��R���'l*�{��F�S�{R=^����|��������N���6yw��nK��2��z��x7��V�â"+4~�+řYiꡪ����U����/�y���y֝��-m�$"D b>0hl�M�+��Q�BMs��ಠ��J�&�.�d�2k9tF��u��ڱo����)�5��fG�΅R�'x#�y
WǨK�h��� �;R-E{l"�]P�w���$a7���������8�O4�YVy���U�(R�i�a���e�3�T�}0D�s֕��شx)}0;��M;>sw=��y�����P��e�!A�ӳ���o�S�Q�6����]�.�/�۠S-$���"XR@�߬�t��u,��2B���U'4��
��1��u�_��(���h[q�5`�9��6������Șٺ0gȵL'F/|k��!�l�"lo���B��A=" �\�Z���U�6����LV�unPSV�_e��c��8�1�ӓ�J.UH��%Di[�ˎ���qeW��g^TY��,x`�ˈ)d|�(�a_��ꒄq�v��2�GN���t��Df�u�T��nV28s�D���`��(���{��e���������jD� �Jz�%bq�PK��#�]d4C��?٨���f�B�A^"�����(�)N������TI�YIڑ���FeX�YU2���uA7JC�@v�kZ�oG"���j�=Z�DmF�P��K���U:\aj��/�Jr�µ�>�Ez��9���A����Pt���
{�#��(����C���7�Q߽
+a��Ĳ�4`2eAp�4ƈdD����#s~��.FƴęA�4�NG���:�C˨{��ۧ(m#O2bsI@���>=]��&��B�����u�r4:��0�t|��=b���]ٖ���'R�Oe�Y�6�h���sY�sCjw��ɚH�(I�֖�{x�w��N�X¥�X���#�6�1���ќ�� YH��J +G�ÚbZ|D�;����n�NR�32�H��s���
%��6����\K�$L*��8���&��$j���W�m�vV��XÜ���O�d3�"���$�jܞF���i���H�˽�!�	
M��o�o�o:��F�DO8S�:W++p���9嵨3vn��]�5X7��]�����#��"�$9�(qV��)~q!a�H�2D��g�+z��d�s�9Sɛ��*S����b&�@�;77� ���4�����4r�|δ��9�mߨ�ۦ'�S���7d�'��2C��w�TO�X\�G�>�
)���<<8X��ܦ;�U`'���^z��B@�[�B�l	��j���˨�zv�E��l@�e�T ?���-��a�u���?2�$��f,9	/�	�kΗ��R�\n�Ejpڴ����1�HZ}rQt��r�np�B}#(�?D
��SX���S�$�7f�b$�c����N&��H ���;�M' w��X�`�7p��]GK�ؘ� ��̘�V�h�b��]�(Ê(���h���s�E�����٤�RLڹCD{%^�����}T�Fβ3��!!��<����e��|��O������v!}�!��z�u�@!��{$emw�X/����G�wqt{���ڴ���$�ZI9r�lw9�=5FKĉV��x{�%�gB*Ʋ��g���ЌA���ݩ����WV�>~�%<��ب����2,���3O��X\�B���<�ǜ�'�AE��u�=Ǥ^���"+K$���T��{��A�N&n׹A�`(uu�L9��㚄�� ��|���`����#���$��b����(K�$�~�2{F�$/Q%��v����������v���?_��z�8�"���8���`�k�0��|Nʬn��8l�͂������c4��,�$Q��Y���O|���)x�Ptv�~0��G�����u���a/�v`��&���.�`�l���0ݏ�=�ڇ0�*�΁�1܉�t�F�6`t]p�3ʖ/�G���*�᩻�V��&n��6ZT}�\{Q�v&x�Kڪ����EO~/ud��v)m���b���qh�A�#��^P��c}H8z����V������rq����w8y��/̳��|l_H�y��≾�UclL^�r9�d{�(	+��t���:c���|�KzABhd�Du,���s�,��Q���};���`��� Gmd��t�W*\��/ꮮ :B��J�UtB�_�N3>J�/:�T��$�eEv7���Br����IT�4�5O2QKb���R�{T�@s�Ɵ�;� ���Q@��{�S�*K���2��觩�A2��A�ך����|1�WM��D��`�T*%�#�ܙ�u]�,Jpj�^E�D9J���X�O�W��WC���bg֨C�]<p{����(�6m��h^v�DR��4҈��#vSR�p�aRW
I�g�X(��C5X&;���K�.����O3w˖8~����]�r*6����1Z�~�@��2�S��[�!;�dU7��u�8�1�Sk��l_�y�n>-#�$��V��_F�œ	I�q�;��6q�.�]u!�D�8߅��de�t2I�-PNā��V�J��BA�o'e�8#OX���{v2�1EQZ�3�Ge�T��ܩ����jI��Е���f��k�]L���� ��;X���).�r\�_i���t�k���A6�9��҇ʛs�̐�ՀY� ��A�P�*Qi��o�?*�S��$�����S�c�Y���^r�Q�rDʻ�1 ��p/4�5��V%��`*�x-��:z間ĕ�$h�t�Z웸��Ǹ�P�jT�ER8Wx���]��Q"�4�8۫�T�s���Ǆ@*ܩT�}�-&�aH1J���#��L�}*0�Q�AN���^Ts���ibW��ed@n�_Ef��R?ʟ��I�_�`�w9�/F6�zQ�?A��>�����̵G�xc��\Ll�>B�rvh�f<r#9y�Ks+�1.��t�ў�⣺X1R�6V7� C���Á����R-�Œ}E����\�
����� O<��#��8���]��u��n+��;u�꺞�g!��O�*��������ZUQ@��d�����h�}j"U�[�B@�;� `�T5u���e��D�㐃��ac�8˽��C����D������\Q�lږ���FP�R�$�j�"ܥ/_�
��uϳ\�	�a��}ab^r(��3Rx�Q�L���Y�ϛsX*�oݛ{1��Bb�?I�we�r���kS`mr��_n�4��Ŭ�����j��zkÿJ�h��O ��?EE���r��XeBȲ��Z�"^�Mq�ӦG�J��	r��j;ޟ\�� ��Nz{$#0�Q��2��'���6ث����_�$�9��M$�PhfKiO���R�MŪ�^��Tm�M���{�[��%'Y���x @7m�b�C,e�包�晷����$h��� Ӽ��̘*3�y���!�����`���E�],��Ґ�Άƪ{���$�s�p�,%e�6�[��
��5����<B�f���%fZ�>_�RXBr�ͧ��q>��V�t5���q���o��S�X���\v��/%8�	Y:<"{yE�Ս��*\L���N~�L��Qjqh�T��*%��.2���D�Z��aJF�UPww�R���=&;��.�⦮S�;���m-��u�k���ʪϕ�d\����'H�Kŀ]�$�1�\��-�VG[w����`G2�V�ꎠ�ۡ�.��A8�I:�>zڨ�r�{���=d���j�z\!�x��'�jp6���`ה���ġ�FZ�s�gS* �'nQ����U����R��g�$������<��=Z?�rx0�Q�Ur���C���㳓�C�|�[����>�_O�wM#�"0,Rʙ�İw�0���&?�����"���,G؉M7���.<V]/Ҁ$H�Am���g3�T���M?=4'�lD�YM�9o�a�؀oV�_���@wx��8� 婗#�߷R��\�i� �ں��\I��A*F��ujc�&�2m�%3���dv_ڌh}�(2)Y��<��~�
�֒��^��$S���$~�<N����
��d�y�%C��{��jF��9�d3+⤃��d:4Dg/�������7e�IA^�Ym�P��/Ȩ[��0:�F��S!R�ǎ�W��m�sѢ��[�ѳ*.��D�z�x�Q���6U����5,�S=��
���đ��r�'�ں�w�d�k�u��h��Bu�Un��UZa���|\	� ��.�?�(��A�nx Z5�=��������\�S�]>GKҚ~���2�鑗�3�©��U�5]GB�g��z�<ᦷ[��s�̩�H5�No��vZl�b��J[�}=��V]�Ѩ̖�)�"1&����Ä����Rj�J���[�.�Oy��Մ��T%�'��qq��v��y1헹����}�������\��6�@�K���G�hXy�J�
��z]��Ӛ���^��[���T�4�Q��7ub����w!���Y֐E��`)h�\s����� A8N��>���!��,��s:m=�ӽ#>u�.15`r*, ծь��@`����f�t�$����8� �������K�W[\�-��"!���|x	޳����TR}fԽ�J�V]�� ҽZ�2�F`I�?��V�L((���6C���o�q�}�b��~*�Oy��j��32ۂ��W��Pz���n�_F1�Q/c|uX�D��`6Q�0G%	�V X����f�ϫ�����sS�Ȍ�m2l�}��v��%�"$�9 ���ۭf��Z�{���8ilV�nu���{?Ѿ�Z;��mDG�p�+p^*�n��'Oֺ˔��N�S@
.b���oW��X���%��`L!U�բ��ou�37����o�i����1�J?<�}PB�;�I��Pi@�wWmQ�L~�7���Q��^^�H�3����]�K����j�5�]_^���p���`c$>qA��G�W���8�晆Qx�o�h���e�BM�j8�?���c=0��NB�2G}�ʜá����v��b����K�GR����4����V�
�%�C��iݬ�,7|n>�+� x�����	��O�a�E���j��l�����d�:��tf�C&`ѧ|"k8��*�/�d��Df�ˌX�ֹz![�6	!ۘ�?{��J�Z�Ά��*� �ɵz��	��*[q
�O! �;�g
�T_NY�BUP�p��;��	���jg�(����	��*p~%ؗ��;��M�"�WP��}
ON�Th�ߟH��`F�;^�VK#��bC�1i�G<��<�%ٳ�r0�S���5u�J���Ǖ�)dX.�I�p$E��\ua�?S�"�ny�� 3��vPN����{*궆@"[j��� <cnT�(�z�Hn5=���ݓ�5 A���5+/�u�:b�f$��~���jo�)ˬ!~2i3]UgB���ڞ���QN�3�#7 �>^�7 Sܩ]�B��u��*�ɢ�Gt{�h�fe*��j�=�<iX�P�����y%u1�u���F[}Z!�4�ޫ�B8�0�eY��������|�j;��8Ɓͧ��e�����F��[�#0�K���gn��<Dk!�Ǿ$��FL킞�t�"��&�O�NU���;���7�/�De���cصAl��s�'�r��:�=&��=��+�0P�m��>���V�ʌ����aY|bր�~�^����Ȫh:�hr�tJ�l�>
�Me凊@`�?Dw� �W��S5~��K��X��b�6Ŕ����~��7��ؗOq	c�r�M��'���3�� �f]dF�w�����Yn�H�WZ��.�Z����<mQ.�����K�jDU��.�l� �?o�>$$#,�*g�ƃ�|h�b@�PXlB������.M�!���c�L*�=Xt��༯~P�C�@>��,���cz;F����Nq a�c?a��,e̎�q����1ݫ�kI��B�:٥�}�z�Vb�E]�����1�1A��2ŅSL�*�e�o���z���9>�>����<�`�m��i�X�Q@9�q���X�m!GbyN�uUߒ֋pq�Mƃ	SKc�o-?�?O�"�̏^f#dj�WC7�U��	%�x��p����gv<&^rp�``jء ��l�������X�Va;��$�i��	�= $%�����4 |؈��e	�ys| 26A��+��ڸ��Z׮O�y�ݺ9��dq9�����'��1��cA '�� &�IK����u���=ԔN�ʒ]3>{����9u�	{!$wh��a��WgΕ��.cմ�԰9����%3�/P�Cև�4�Y32��3��d:��[Wh��Eޓ~��OD(zD����'_���U5�HIޟo����Q[��`"{H'��؊�:��CD+�
�<�ݹ���iĸ�G�
3KO��ǝR�4�X�<���3��	����k�[s�G�P�.u�������(��Bbh�?�\�������*v�U/���oEʜZ���~�{4�s��������vm�4�ǀ<&���ݰ��6.��!΂��m��v=���	��1���p�/�5��
C����Q�J��bd�Ps2g͍&�*Q�� ��fP�z�$x*�#~o�¨N�G0[uS���n)��d3.~Kç�SXz]���U��p�)<���$ո�_Sb �+X�0��)�qi¬�ښ�z������-�}qw"�F�l���u]~����Y#3j�%y����lVn�_Z�~�B����d�qTm��61�a���>�4c�RV���p���B�N���Q%���}��߄��5�s��]1�EȀ�_಻K������ �)��E��M��hȯ$��{8��"	RmjA�� ܥ�i���,9�3�e�����k��(�#%c�[�:f��o��"o�{~�}�e��8�P�(��&�u+9��e5�L7�T�e��x1'�u��f�0���3v�)�������*�"��&�n&��0v�����O8�Ɨ/�����Y�2���7��d�*6�1 ۡ9*"�J��\��$y�d� w��*	��q�^ӬU|�k)�6��U"	���`�$����<��6���9y�@l�2�i@ћ��6V�I`�B�0�zw�í�lLI�xk���$0�Ke��[/�~�z �~��~����Nr�.���� +I�Ŵ?D�7�q�}M����Fm�(�k�@��,^���7�t�({* ѧ�Z���£�;��4��7��OE�j����Z3����`�B��'�6���M�y�iYֈ̋KO��/;vx�a�%���*(Mʍ�B� U��{QҺ�A��s�tt�Z�8 �f���/0�7�����6*Z<�k�	�Q�Jd�eS��Ʀsҁ<�z�4�����KFJ��5�=��L�NJ[��g�>FRCW]H/�ii\ڠ�5��E�n�&CA&�Δ-�F���͞GlM,�:>��k\�Wp
/�l�U(�S�Z�ޖ|�3���yr"R�y�˧���nz��7��0'p� ,�$F][��RA#]b`���e,qr����ʵ+!����D�YWD7b����Sw�����m�K��#��5�j�ik	͖���������A��i�H� �]���B)o�W��:Қ3�;P���[D�y��p�I�u���W/�)ɉ��w�gK���ϥ���9�#���B<�R�2���C�`�"r,j���~�>�������x7Sd/�P8~�?�u���$N���V.K��Ί2gEz�zSz�J@����HB�ڲ<������,@�Z���i%�
	���E 9����Ӆch p�H3���6�<�ah�0�Z>�ӳ��W	\�G�̃.��������sCs׼+�g��[1aa���P*]Ԅq���+�g	�bK���6b��ؕ�lǄ��FB6��6SiX�o�䓾+�'�'ü����LOIj1M����;9y5���!�{C���=����y ��%^��,ā�jw�E��2���l��)�����D�E#�߱����H�om�>��D4Q��S�vC����b�C�S�o�/Yq3(�̝_�EF)_�`ȩ�Kle��%�R2�����H�"�F��Lw�X�ut��+y�ߕ;��P�Lӻ,�Vi�<�2D�) �h�c����ք���0�ҡ^lQ���V.i/W1o+���W��S#1��mZ����īP�9���(��l�A�n :���e!�6�"M
%�2̒�	�䐹�7�(��o�æ�:�����B1��>���9��:DX�����Q�S�8�B{e�ܝ�������	�{������*,2Yo�҈^E��/*��A@pE�Kj2�J{X�����Z�Ҙ�>�����[�����o�n��Je9�iı���L�m����]|�sĢ��j?p��a��Y��!c�!=8��J�ԋs�6��F��o��� )�:y�~.�K��������a027yr�*<�=�Y��)�^w��x0"�U�E�'nV6��^�W#��s鴬��\7���jne��<5�K9$�=J�J[�Z�8���� Y���[EXE8qx&��w��g��q�,�@7��u� /����W�w��9��_Ch
$'Z�%���B3{��ܷv�N/����e:dH��uQ���	�/�|���P���u��܃m��N�r2n�@�5q�|���z������M����CJ�"an=�krn�.#�;�}Z*uH�M4��ה��s�4^���r�֒�-�#��3�]@����U��IZ�D{7M��恜�mֺ�I��h�]��;i%PL1�d�D]i��Ϲ���Ԥ�j�;�m�4�D�W)O矿f���&@�����EMTu�2X�J(�I6��h����c(�<X(vsꕑ�i��F��w|o���!��E16T��a-�Gn��u����uAq*C���}N����ug�@Z��O�UaZ�-���D�]�z9������I�pȂ���� 5�U����}ӏ���ڇ�t��I4wnb����}������-�v�c��~Z���v�89?�L?�QI=�n��/I�ǔP:�� %�\�<��ZcDq���mk- �J��Q�~�DP��Ѿ��o�`�3/�~1�Y4�p��G^�$
vW}��|���	��+��n����;H�9ye�x����`���i�4��ᐽ�f�78���c%�SAw�۵<^�I5�kown��	�Y�괁�l�[XY���4�x(�e��9�K�x��cz�vP[+G�ќ�@��'C���C2�Z9ǘ}^}�r�?Ew�	��8����%A��r(?s�z����1U��G�E�F��#{7��_*Y8���  ����7������UƁ���N�V�҇���X���p��}:�&7������<�@�}�I)���ä��l�����Pe�"�^Ѩ�'���'��>��%�p�'���5G4��;%�u_���Զf ���f�0��%<@)ѕ1l9/�U�+� ��|�퇐�	ꓰO9^.�oPT�z?��E}�����#�:O�E�yP���YC���>k2����TS_`�s���`��.������k,)�9��^>�ō��*o�*S�?��� h��)A������Ɵ2J���'�h&����x��?{�@�f<�Ǧl�  P�tuЊ ������I�����]Tx��=>t�]�	���)�0CþR�Y��D�N��C�F{���(�כ�(;�ҳ%2k�K����1���P��eO�(�<%�p���=�*�s�8_m�Mt�6��w☠.�~�zaڡ$	B��� �|���`r��A��΂�xw$�9u��O|t��]�m�|�̛"��9�C�yus�U'K��'-lE�x>�7P͑r�Kz�D�ՍY����n�Q]Y�B� }�(y+�X-�!�מ��Fo�����ŷ��V���c�F��#�h�#��l���rȊ{���t���Z�3P��#�N�q�"_�Љ���Gv:������-�M�$�0y��e6����j�_��"�������|�2[��5�PX��͙d�R,�Dt���%��<���[���k��R�rj�~�R�tA�KM��� tK��!����o�b�Jl��:`D8�^��/%ߋ���/|WM
5-����+��%��өy���c�`����/�(/F�����^?�	7E3q+�PhQ_��7aת#�k+�p��?���JCOf63�����S��~LNVBr����˅Sv�F�;�_g�mH�P