��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~ !�s5���(m���0�=9�n;y����'�O"Qa	���}P��7D�+��ɉv�0��4�N�j���z( �;B�:�6=����h;��p8�n��W��m�?��b�B�]3vN}6z�:�o�3$��;���h�ג�~A�w�Z3.M���ѱB��%��>�ЫT����p-�8z�i!1�I?��ѝ8g�
��-}Oc�bV�ynƃ�[�i�5��o��^g8U�2�P�+���ZZ+���՛y4,M��6O�C�G}ˎ��?G����e㶐dc��-�?M����a�r�e��X ;��Y��<���v�a�ŌU3���laH� ؔY���F�e�lY��Y�KCS���o<�OK��1�<:ox3q]_c/1uj�-fC`+�c���T��Hl��c��L�ъ�0�����M�@-��YT�d��Olu&^m����8��?(^n�.�>����c�=�0�9������4�C��[o���ׇ^*��怨�{�ſ�SϚ�)<�I�u��9�����D� h#�<hu=L�Ϭ��mPr�Y	�T���MW���m ���x���� tR���� )SD��%�y|$�J�mh�Mh3�ؐ��&��<��B�9�ۮ{l���X�ݠ��	�;�_T���ϊn�z�<����7\��D�v����ذ\�9�u�q���\�+��-��7fP��!�u��R���>�\PUIl���N��B�u��W`��H	�r4( p�-�
r����rcSFM��dJb|1��)�[O��|����>

\����ƃ�
�K�'`D����R�R��v��B5�T:�[<J����#��L���VJ@� ح�K#���!Y�0]���e�!��+�Rk�4Q9��[rd�dm/G�$4�~��v����o��=J>�������
56������{-R6������/�$���1��mWgG����&�X���LϞ }:_�⠂�����aa�]W�.JF�xo�oIt���n"��1�D���'�����j�J�x�h����-m�<�Y2h�Kv�j^N���C29;[6��@s�`׵���ޭ���e-����$��(jԅ �����N�����l��p�)~� �2.�Al4��~�1� EiI���vsƾ���C\�������38G�q�.}���و����^  b�Ǔ�[�e�?W��V�����;C0Ѽ�6���D���cN�Â�X�r�V�2��)���[t\�T2�i%�on���<9L��+� y���G���U��b�]==(�Zl��,Z��E�l_�O��+X�ᙚ��K����{�����m�cEƿ�m����<�,4b��r���0d�U��������fA�Z_�X�7D����^"ӣ�@ʍO��G�{c��n��i�k�Ԯ�p̢��X8l^\n�sf��U��X��$b�L'-�Z��UICO <BC���h���Ei�����\�2hxg�S��wh�Η�?Gr~��M��b۾9|�ZЀm��:5���]���~��*�qza�bE-�-�
��J⟕Z��E��zjw
��0ē-��vZ*W�����12dTO�ϟP�`����(3M^�Ok�/�3���$�v�y��n��=A:�1AU������7�/q��>���oq�0_sn���A�"n��S��hM�Z'����.T�1L��^�n��"�)��g��q���G��=�_���Rv�z�B����l�� �,n�G��8ۜ',L؂�K�=�ǽG�q��W�Z�Z�՚�w�Y��d�v#��3�Q|����P��3����cj�����I�*mi�9�	�=H-�)��",%��}��ygc��f&Eʛ�(V@�}�D���j�dŋ���b3��C����>墭;5d����S1f3+��ǂbM�\l-lK2T��DI`T�r�yH9qw�Y��n:JyaA�Z��u$�ь@��S�� �*J��L��Ԩ�,V�㕋�ȉZ���J��U�b0	���1M�,"���.�C���pm,R^u���K|{2����BŰeو*�{x��f�uBs�������jz�9��73bL!�+S��/�s�O뚹k��� 5'�c�)#\T�S�x��Q�si�Xi��ۅ��>�|�]"J^ƍ�Z�/L�1y�����.��@e�(Z�ų��#=����7ҹ�M�A� �����&i��~�rx�'�G�A�L���*���QbQ�2�J�Ӟ��+�?�^��`�p�����c�Ռ�ʥ5�)o[	LV��9���̚�����u^��/�� U�Z���d4/�����&xzp+�G	�r_��D1g�9��$#!������`���L�6��%<	�u(aH�23���9ݑA���J}��a�M��|���T�T��Fr�E����I�j^�{/G��e�F\���U)*7���ձB��Բ]�,5]�xu�R�&M�d�o��2w�N�X��ۿec(��3A
ϸ �x,>�$�hΞ�����޼Ly;K=l���$�����~#��bз]2��a�R���Yt,��?ΌB% �<_nY���L�Rɍ٘;��c���>�,��!mJ7c�ƽ�{�܎(���`[�/�U^��gɿ���`(�B��wՈ���}A�U��V�FxD
<y�����JD��rI���DY���-��[3�>�"<J��d�t�*���:�TBJ𖛉%_��C��qO��d����H��6�K2��]�8p�w
f1�%b�J�T��EݕY��^�\P��.�%����8�n�k_��p��&`
�����V�q��1��]��L�5oT�%@4^ո����EW����ZX@��+B��_�oqg�����{y��ŉ1.����M�v/��m�lW"Ij=Ǎ��wcZ�h�e��z��c^%�l��I�+J�� �r%|I��"!��{ēU���y��G���f��4�"Ȇ_"�����������6�im
���Rp:G�-�H7�Ψ���ؐ*@$q$��z8.�_��A�s3�>�
�(����s���}�Y7�?�`� ��	(
d§�ד�#�u��aP 	��ܚ��X��`�����N��M3���B�����	Vm�, �aE�v���<Pfq��,���T��Q�4m����[{�~�`��:�B���28Do{4>fU�/R��UI[�.u��5  aT��������L�����C��O(}��H���4O�k"}9���T���S�u`vC"^����y�m����`WDn�z-vDq�hʍv���?��F�x�:�Sy��sP��<���w]L���\��v�٣;#e��I�0�������"�z��m�ٯc��B��TP��a�@��������a;�ĕ8Y:Z �V� ��6.أm�>��󤅓��쑕tf��R�8^��fG��r�H���3��*[�4����,��Hd�1��W���e��bJZtߣ���D����m��p<�7x8Q�;�a^��6��^Ѐ0�"u���C'
���}�>,�K�(��_���4�
{��Ė�����>&�i l�	t���X�P� $P�P��0�~|�Y��-���#����� P�ڀ���C�>�:h6]4���ry��xb�gMRDi�ږ"�gY}Nr�)�KJۣR8	ɫz�]dO���,N`�b�����to���}jFɨ����m!R%�FB�ԓ���Bw�� ȸ&�`�	��\�^}�7@&�}���iN"�p�[��H	�s?��%���^L�K� l��@F�I"q�D�/h,�1�e�DGm��|���cBs�Έ!q�����!����t� ��Yx��?��?��rd��D�d:&�"�K�ޞW���-�x	�>�O>E�c����+5�8��[(gDG�C F+G~��dɅ��Ů�y ��-b;�N\I������4_c�S`�%tu��P��*��h����4����y@��VK.�@5RJ�D:I{������\8ė�9TЖ�]O
7G�ᨈ7oz�I9��S�ȫ���+TU)�B?@�=f`�/�qD�tl�A��@�(>k�W�����Ip��XBu_~�ϱc@D���#H�j-2�X�*kAA`��U�b޹}�O�s`��2&��]�3gL������T/ni9��ȭW���5��:��ΜJ8��-��V֞F\a�bz�-����B��E�1g�����*�p>V�K���3�*����].���`y�EɹA�V�>\>qr�g)̾�����ݬ��I�U�^NΩ��I-��/�������b����a۹�	��j�bu�V~⌑0����@H��L�,�Xy���IM����FVÖ�a[��Uu2A<e�X:�a?4�q��Є&�k��&�)N������(+���za+��h��nJ��8�7<�M������\�}O��V�Q園�kzp݄oW@��
�!5�F���h;b-	zޠ@�t��n~��J�j?2<�sWU~�󀿑W�"�xZ+ܘ�[�`�v�������?j���#��:cA�?�F�RU���SU���?d�� ��o�G@l[6rĆe�������2��K:T��g1�DQ*� ��	#R�p����z�*�D�^��:0Zr�G�����DK�vA�ň���ǌG�1߶#���brȬ�5��v����D5Q��W2�0��4·�[�>VӤ�,�`�D�`VQɧY�	�=�Ֆq�c!��e�w�\�;%<-˷��Um�����ױ�P��PID�ݓ��_��4�C�`�����77���w�� IB�)���Y�5�</�E���$�J|[<O�!���d����C��rB�LX�,�� >�j�E|)��:��������a��Yj���b��Og�$����+�mT��{�<8E��4�!�,���t��9:_��ոnQ�Y���H�Q2O]`�R7g���� �0Lk?M}?>���I���BXB����eQp�\%���+��g�e�� t�{�R��-�e�I���}�B�t���Ѯh����ܧ�)���/䂜�����i}[� ������w��-�{�KxM�����S�T3O�l�;��:!��#��`�)H�t���
~I��&�o3o �8|�D|޹7��+c4ګ������VeG�y¶t,E�x��Ϫ7؍8m#�|��`L�_�W)�Y���_�'�ڠ�N'�E��e���4C��S��eLDDQ�C����;��WK4X���nM��x�Y4k�������ꑸ�s�~���ۼt��$�V�x$�b
7�9���v{Z�wTt���k��&���Oy84$$����q!=��u4P�:�.��;.A���U�����]P�i�{�F���I\;��Qf�鄂;�ǆ`���K��.*V4���H7n:�3��4L��oHsE��2������f�Gl�z�aLW�5749����6
ߙ�aA:��x��M��/M�m�-O��(g��{�	ҳ���?�+�cզ7�'~
��a֛?�nA���r{�c|��m�*Og}BiF5���m�Ow�+0���O׶&�0`J��77���Ӝ�����o�##���O�
�o��a�YB�S��[K)�u���Bz�
GUw�x�s/K|B����\fՉ��9<��ª�fk���`����Ξ�D��/C�t�㼘��ꕚ�ݜ#<���b�&���~Fs{��D��i�� ��wO?\����WPJ�f��|0�w8���e�	yI�fb\%��>1I� �f������������f⪌���boc�4�TZ��#,/Y�.�>�OT���S�M![,�"��9ºL\�b�T.��uЩ���:qA��hpEP>����h�e�*��yDo �z`*�*�'|��P*8DeAE^!���j�EaH�ԇ��m��t/�xu��c�F�'E�;�GS��/���&�4�𮺚x� `}=A�)�i¡;ۜ�(���$nU���r)A��O��_�l	앓�"�
��^]���Zu��_��,{)��*�%)-��<����;�ƪ=�5M^^=Ǽ0��S z/J�=P��Fs(#�(��S�҇���Zg�@�?�O���TG�B=�#����V���ء�����w⎽���-�A�q~8Q��<�� -?b����8����s�$��LUz*)�f�-����E����g���6��ث�5��\B��նn��M8�I���$�ei�|ʐT*��@��f���#G�#x�<Fz*��Ӫ�P=^�I�녭���~���^-�{JRD'��(��&�,~�ĉ�0�e�;8���*ǡ�����[���lTI��J8+OE�.��#u�1����gL!pb� �i0o�' #��j^�Թ/ט�&��n?���V�SJ��+_��J٠yDq�QiH�U���Z n}��>��(6�a��"�$0�a�Ng�n�e�ѩ�'��_At_(��ve=�`/��ґ����b��M�cM v��d"��3�̿F+;�,�kh����H�S��6_!�/��W�/f*PD������<	�/
���ぴ��R,/!����Ǽs��mј�q�B��x/�?Ҭ޲J�s�́T�Lv���prz2M���Kg��O�&p{7,Ϯ0�~��X��r� ��㍴w��֓Ce*���i�o����������۲P��"�&�+��'O��1��fv�+�fL�aG�♔��kS��Z�ci�YF��Ax�tp���˕�ԃ�F^�C�l�z�?Za���Lc8�ӎ�s`�=���H�k��|�}p���=�N��i}��a,�Fv�˻��(p���~\��s4%q�(�#���˨򤩐кq쬎J�<�g �U��w填_l�d��*���ƅ�h��w�{���Uw���Z�3.Mg:�
���q��6}�?#�Kzl6���E��1�2�<%�J�������N�n�a�QAf�����$낐 d��Z���,~�2mS4�==�z��oa�4}$�Scdn=&���BU��y��Q�&&yl�!{�4��|�5���a�k��{Ez*H7���X���`�h~INTҋ���s��9PbV�
��Vle��M32��4�?L~(�LƜ�����g�	��d�-��cjE���L@����;k�3���OM�n���!,3�����kS�t��\2�u̇��6���n½�Ry��Mas�f}8�W9�dRk ��xۓΉKI �x�����x��>�d?}�G��yȒ�P�]�Qb,.�����������j�������'�� wJ���S�|ȼ
#��������;sZ0�o2�ƶ����X����¿{��W�Lf:~
@�ŉU����iuS�Tka-�2�}��l.lO�����xw��խN�"�"�Ƴ"tc�O=.P�Z$�ZS��/��K{z��hnX�v����@�N}ʤ�	��N����
���3��|�38��ן�TE�`�F>�g����!	h�U�)g��J�������m����쇕d~�B�^��v��	����I�M�1�?�1k�R�%��$^�\�#p&r4��q���Bb�I�5"Ag�%��rGi��8����#]�e4�y�&j\�jat�aKm.L^�aiχ�j�8Z��G˧�r����4�f����������OY�ǅN2m |⩜F�J
�N�Jѷ��Cr��C�)�YZ���S�CoqnU)�̰Jz���R�ղ	$J����� ��r�u��.y����$r3�S��=N�lD��Bd$�ݪJ�9Rw���&�1Zl6��\Z�t ��³H���k9&
�wp��*������#��>g��^V�2��LNh�'7Ɓ ���W��?�Q1O�M�VE�2���ax�{�QQy�.���z_���-)�%+X;�^�d��EW�m�O�8�zD�;a�08���)�nY�K���Ԕh�J���2]��u��z&����ޕ�<8ٟK�[����s����p�p�:��0e�_�8.qȜ�IU�_�Q���u޴������xR�/d��������K���D�"���V��g����斲)>ԡ��.�hԼΈ.̿3�c�$s��J2�7�UHN0GD�C�Lq��r��8�::H=���﻽�'�7ʎ���E%b�%v\�i��?�&��2K!n�\�Ȃ�lE����Q]>� J��Č�d"rޓ����{YU��!��,d�R87,�.����ҭ�����G������)9��B����e�򈲳m�綝z�����#$qg��c��*7_���	�H��AWtc�Xǡf��j#��M'�L��O�xţ1�5h�G����E
�(�(L,j!�e�zɫ��%�ـ�;t��Oc�?�{���.}{$��txNy�G��i(��n�	��!�ņ����wȞ�����G�FȹGO�_j���νHae����5�6J�f�\��x�A��8��=�����^S�A��>�2
X� ��r�rt����SCK�!�6�s<s�w/��3�#L���*��V
c�4BsW+����C�����a,:&}a��6�9��x��Y�\R��C��w2��.I[R
u�;XX���r��wӫ\�»"8U����g�o`����:(���7�B�q����잦�7�����a���,*���.e��Xh���.?P�>�Wn�4�ҳ
:;�mxo�C�s!oÞ���Rh��R
Z�� �	RCH���|;�t�h�M�H&n�]���m<�_R�C��:˰,���\9���m�!�ojjI�D�)�* �)9T�_�����q�2#䌟�Ͼ nJ6~��= k��Xf���Pl&<k�v�=��T�C?�w����]A�Ac�)�hcr<���2�����/�G�J��;���#mU����Ԧ��m��쳽�;��Rm�~���<��!s�>��q:��[~���j���l�	��y�"��[jJc�%�M�̾���������d
����7-���i��Fj(@��$���u��^?t(�ޗ@|�Wj��9{�EV,�_G�/.����Ļxv�-�Wu}�lSS���"����ޞ����m�"	5���i��C�ȏ��K�%�2��Az�zLZ����_�ψ��Jƴ� n�s�3�y;��������ԯ��g��+�� a�İ�HQ���;8˭0?�'�u1wk3��P�#�q�%7�~\Ne��Q�Y[���0��/��y\-#����{���DJq���;��;'1�O��Ԋ�ݽ���Hp�m��a'dHުi[-�y�G��o�X�j1V,̋W_?i�/�D�.���7kq=�89�6!T{ǥ��	Ϗ���+�j��p��A�1�	A�RnD%�m��u�.<�8Ӧ|�����<��!jQMv����Q��/����F���������[����c0qbJ�ܘ���ia�͹�~�UH;�l��TI��+悯�rTx��8萔���j-��,y]��(����Bf|q:�s�c�7;]t�9��*5��R�G5��P��K��j�-*w/���0�=ķ�y�5���	*��d��N�Ͻ�07�x;u���q{�"�w$�q�J�����@De�Y���U*�"E�q��ɞ�O��Mڰi�V��ާ�H���%&7 wb��7=g��Z�Gdk��>*a7�*Q�1�K�:z�30n�ø/�0A��Z���Q��!�Ŵ	����g���p�TXzK�a���a��"5��+� ���ȡ�y�n~'�mn~�g���]YL��9�?�;R0�@��#�(sU��xX�P��� {_����P?é�s9�x�ċц��rݟY8z�9��x.�IV���
P�G�}M|a�.�vyb�Ԙ@�"Πn1&�HZ��/F=�7OW��"uc!��HW|=��<\ܐ.�x��ć�Ҷ�@vkH�D�Xm���.�7�$ǒqQ�jz%���}W�{�W�b���D\K���/��Om�^�eN��9��e����V�]�9���5�IM����Y9���!ݼ���.hf*ǨF2�,Iӆ�a+�}<��v8���?@Eq�+*���J���������k��Jv~���a|�ʴfrN��U�&���b�N�2<f���kFg���9��a��б�-R���& XILB���J �2�E� �����}� �u���4&Xhj}A��%$�����^��#�T�H��CП�����<�'�����-�(�;����*�x.�� m7~D�5I�wH�az�,��^������nD�r�<���˘�Pk���0�{a��+i�����恘�`B��d<��Ѱ'�dߴ�-7�HZ��= �$6}�0�=9 �dp���K��=��^rw�F�#
5]WP$s��0͌��kM$S��S��X<�@����b���h���6���߼�{���Z�~��Д�������\�̃[�Ƣ���p.�%����K-���H�泻��ݫ��we�� u�A�̩���4�S�����L��T��GR�} ��*ܾY�,Q����1x�3.�i�����S��G_\z��J�,�	���`����g�9�~4��&#�$m�j��)�p{/%2��$2���Q�_����8RB�؋ "��>����i��"S�_+��?�t~�W��[�
./�C
/��c�Ƶ�'۪��=c��h�
�{��Zl)��"��t�90�x)�1�X.=����ŕ��_��|�5}�����1�V�0ȍ֞�T�q׭����`���09�N��°�{þ����(f��v��}�{���:�q��Sdo����/�^�����|��K����^�ų�S�o!�2�3�M���vE���mcU�p@C������!�.�:$&<���"�N��� �-J��T;�	c��\��-��K�Ov�惞4����f�t[��q�a��׎-��o��g(8�7�ņ^8��Q'ٚj
Ħ�`���D�Ǒ��)�	�_�6},nqo��g����"2�h{X.Hᤁ�C�LI�H<�ϝ)�_^N1�$�./���󊚡��6�|�kO�&d
Qz��f=HxwO,�R� yAMe �E�32���F�6�8WNt� ޭ�S���v� d�p�.󥡄�֌��y(HH��\�+�r�ȝ��ƚI-D�����߮~��&���
�>�5��0�--뷤=�ғ=��]���!�8	cy@�b9n�_0��y��A��%$�M���4S�YC�-�p�"�,�S��2fʒIJ%�I�����y��&0T~�>�0�4J��<<�͖2K���n��A�C�W�pf��vF��D&�<��Zj��=������7�U��Uן�Uw��)-z�U8;���&0��z`cFx+@9�VJ/V�gK�=�0�<���w�O�Y�^�u��X��A�8bA�S%�J?N�{��.G&&����Ȋ��[�ȥ�к��`���Ԓ0�EUG)X�C\T�J��G�%��
�{I%mؓ��B��;QZǥ�m[V�"�ρ��n�i�F�E{8 V�[��͛|�4�u�8VC5��_>������fMZ�A���Յ���=�O$OLZ8����}�ˏ�?;yU1�g��˂��\�<�ڈD҇9�S3����HS��Tr*�� ]�+�> ;�����z6���nf�ֳ璳g,��������y���]+���i*L��F�"}���s�^�k�n��%���=���}k��3y	'��L[L�w�֯�s��ZcT���F`�+ƤV����Io7��d��ER���*g��[he���ڼ8�c8\���R��T~e=���Fo�
"��i��,����f�h���:� ��� Y��t}�ѭ�c<2Ǯ;�oin[����J�>k���3~lQA���Lc���Q���@#���Ql�fdǤ�0eް��j�&r�+��wVk;R�.����ص���t�k��ީ�Nsy����la��?,¿%HM�G��ɛ"��p�T�}[ԱH~�A��f��	U�n��Y��;�QA��F���ۂ��\^y�ޝ�������P��!n-D甌=k�!�xՃ#�}��FC���e����Tv٫k�,;�C6g�y�'�QY��S?� ��K���t�|9�ew�0!�:�l�5�-/Z\L~����҆,�K���f���Ŋ��� �a�J>��O���A��Hbt����פAƷ
#+8�Ԛ�,��_���4�dJ��h� �����@	O!Į���ja�+[��p���l�)�Y�{/��X ���kĈ}�09�.�
�$`����2[S98������M)�C݈�=P�:ȶf:{:�Z2|���2���w}��MlZK_Y�ͰA:G�8���G�42y���P*�7P���$w�u�m꒿��`K�݅��T%���x��z���;d*qu#���1���gTuл��(�C{����!������X�r������f�f?�?r�6b��Q��w�:k���>��m�IQi��ڦn]k �גK��}/�B����3�'H|��=�H��Uut��J���#�nbq��W��|�O�2!;�)���r���.��9��i��y'�Z��!q��A�Ց�RQ��|A���꽈�4]�[��%��⨢.Q������	�,##�o]ݲ���[?y��v1�t���oA����"��J�7�%)��Gu�{�S����s@��}>�:Ҡ�!X]�i秇�;��o_�Dw9��"�9��\�}c1�16����_� ^$�i|�4��j�-=��gV�8�)�~R���\T�L�x��{Ȅ ;~������V:�5�����سQ�:�g�+�ޒM��O+��`aF�p��00���W^�?��.t�N0��v��� ;3J�����~�����b���TP��I�1o[�T}�}~�+hu��p���Ew��a�i���&����<�eQ����J���30pxSG:��Q�e�&���0�%�ɫ�j9}au������-�yUc�
;�j�p��8�Ʊ�4Zqj7���|ֿ����ӆh��)�6�x�����{��u
oN���c`�r��ʦH�`pmj�u�sʍ�5|;ǆ��.	2�т���b�1%q�
�N��o9���0ӝ��s���H/�rp�*1K��Y���8��{�����+�풰���-�K����ܼ��G�H����锕҆�t������4%Hs=^�7Wpf���N�#�����9��.�h;��nX��Q���J  Tys�/�gԬ/�I�c���j���:;�xtw���8D;��R�]P��c)�"Bl׬Pe���B8��^2��A��ӄ���LM����e#9-t��Xu/�jT|��l3�����q������	�m�&��� W3��2�����Ww"}� ��z��������>ۻ&XV&����"�cp)� ��с��c5`;�[��y�7]u�j�廥b�7�}�9(��ɦ�}�br)^�pz^ �Aݴx���B���}�t+[tW����s�jg����H���a�N�3v�{���2n63�lLlQxX6�v���.��:;\���_��0�6:ܡZn��Y�.�$��,���O����	�c��/�r>D��մeKI�<��hu�j���L��y�B�pc�9�mhV>����qq�K�%��.�uJ��"`��L��E���O͓u�Vr��,]��[鉹�⠡D�=��~���##���
Y����9���z��R�r�_T��I���?+�������`�ޑ+
����4J�X�"h�;lM~�mN�O�f,NC^��L�KX ��~�V�~k��v��^�hJ% @t��>*�&UJ���{�O�Gv��!��� ���@)�^�Vd�+C����\DL���=c�&�&m�����'R.@������(���>uy:���/�݂I�
8�� Q��D_��C�ƶ�͠F��Fe.C�`��c[ xJ\y���*xQ����:�	�`C��蹶����6O8��V���,#�h%��`~Z�<3��V������?!_}�b�<�M��M� �}�!N@h��4ï�v��-��!TM���^3I�_�q��L����3��^��ɫ����o�jx���Vx���ܭ�M�jʎ	�|g	�f�_�YL��@���(����h�h���'�6ġ�� �kdo@�	�.��Ւe��סT�	/l�/d��R�Z%%"7�K���)1Z��f�Y[Ek�b�W�o2�I�?�$ȗ��3�������ݲ����� e���,�E����߉{�e��JK.��2��c,��>���E�_Ġ��[��3nϦ�"��'���V:�P�6�կK�%"�O�h�A����h����'d�SyK?�P�,�I�i/���$G�2���r��V��8#��Un�1�)j�Jt�:�w"n=�	{�-�r�!mLm��b8��m*�8�t: ���U����_�d��5L@������y���0�?qYT� �s.�bE���C��n�Pz���3�����d���aZ3��z�:)���^��C���k2RqƱO>9�u��c�~c�U"G���Q'�t��>>�}��lq�tE�^�XV�wD~�����.����(�a��M�<�V�w呐N?t7޷���8ȡʓ���Sk $�q� �+#W�T2���@vd�͡�%>���;|�L��@�� �YLͿY��&���x֩&M�/e�X���Rzo� �5{/�0���[$��և���Ec��7xTR�z [V#rVx�%�t�Zo/�>R`F�x�>��޲�dUWFY˞�6�+��"�ĕ#�*Tz�b����q����Mt�"��^������JfcVt����� _�S+��t�I�j���ɀYB�ׁ��G2{~�TCm����W�!U��k9u��Z��D_�����(��0Z��8�;��:���0���1�w�o�'�rv%��\Hm��!�h��l�>�}+H�-�':�[��-N�|�l�8e2��ϳ*�"�NO��w���uә�ڙ{ҩ3��&".�;r��752Σ���v��S��?$���tRv21{��Ó�c\�!��T����sQʹ�|��N��.�V�p�CjRU�ۋ�Z��J w�݄�5}{7�m�����2��2[d����pJE���]�7V��?h�QPRnZ��J%����0���WR�7gl��Ֆ�]ˬ���*�P��ɒX,$%�!c�X���d`.o���6�����"�X?>-���M+J ;�GR���:�\�A�"�6\�G&���Y�Z\��Jʇ��=���Y�n� /��ͦ� �	�O�ט!�p��Y���ˈ���b
2��FwƓ��n��Bk�Ր��%�9������X��5�x�n�3�vY�@90Ĭc��#��^��l`Â�F�.�a^#=�=B��驗S�L�6�%�C��S���|-�o���Ct1F��7p_��Lb�ĵ��:��z�fX�? M �4��3�`SR9�meX%��u}�+%�Kwi��ɿ	�'��٘y�����C��v(���)�\ Ԫ���㋄V*P�Qk��:���9F�y���M���;�,S�d`i���(��m���X�H-Z�S�$���>�q���R4�j��T��11���IA���'7 �հ{BT>O$gʆ�d�*�V�JSm��Ԧ�y?�b��1isP�z�C����������.�U$����C�勩h�u���N�eU��I��5RK�N|���繘d*�/��E�5�1Z��}�k<�Up{7��oc�]�roZ]�aE{�����D�%��Hi�zM3)��$7 ��}2�E� ���w��};V��Ţ��Z����+�﫥��;2q�zK�I�&�%����l�S��Z���u��fHE���gY�g��D��M%�%���u`)��pF�G�Yk��u"d��(]����Y�ҩ�pq*{rV��7��#2�4s<{0eZ��t/S�<�"����Б5�Pw�J�ر���zΚ���i&��:Xu�z�t�s�/;	s��C�BQ
I�D��O(q�P�N�n~���w����s�L�3�l�5�IUmw���IXq��2����M�JYz%���_��+#1��eW&��w�p��١|s'y�k���;ӝN�uD]���G�7�ɿ�	�ߕkA9���jڸhe%��k����ۺ�	��Bz�ZV��u�n���X�{7��@Q'�c"�kS�1���K�����XT8i��n��O�$d��8ΐ����sxVAw��<�p�U!��bU�,���\���n%m�B��)�*����,�9੦�)5O�6?��5�?e�tn�����c仪��40ل��ޡ��R�p�⪛/B
��T^���L�~��bX��[N���	�ڃ������[�R���[��3���qf��3�}N����P�3��Ta��������Z��щ�BQ��|'Ye��Z'���� Tܵ�:�$�_#ɢ��Q�!�����2b|jEe�Zb��q=�~?qR�}z:w���s��ش��"�.�JS�o���X�$�;x+��:x�w���yK��[���pjim���L�OAz5h���?���늨�Ϙ߇2���;�$�B-���?*D�e��5l��4b����:���P��3�2Sf.0��z�}8�,��~�AQ6gD� �����D���_�ٱ�,�j(9\�k�O�G�l��z�{~�p\������f��H0>m�^L���:8���X��z;i�����y�u���g�~sg�(ѨS��{D��.����A��O������<�}�3ݶY����{?N���[��y�4>Z߈����f�o�	w,�xO\��׿*�� U�����6�=�
Z�4p���K���F�`�$����톚��w�3��n�������A-�{��+t\ĳ���4�{�_-Jܘ=)TRGCu�Yx�>���c]~������b%sC���S�W���حgJҼ��\�^N������k�.�44)iA:���r(Bod�W��	)0z�#����C	��ڳ�УFId�4�*y
�������IyP
��і�ð=,�����5n�I P����]^�f�Bbȹ0���{�Y�� �7����U�'� p��IA��$�Zt����DJ��*������GJ;8��R��S)�0�]k�=�ZT bA��%r��.��~M����O��v�/E��4W�:����@G�@�*���A;8�Ո��|II�4o҇�������&�گ'��%
�N���H'}Ka��]��Qp ��zn���n��$��qy�q��yo����*�[��j�UۣF�v�!����ۖl?���2TLJ�umR��%�d�8ڨ��͓�}�'EU�W�^����(��&LB�}P5�Ӄ��!� �j��ɔ�0О))��E��{���j�V`�cV`N��J����}�P�LX����ׄ�f�NXV�[T�2h%Y�<<z2vE^^TP5�b�g&�.���N��l1����Ȁ'�}&uE�U�;�Zl�l�_O���������[����K#6����K��#>S��Z��Cg�؛�y̱�������H��fW��0~;H\0�z�G9
�Y�����5�^}A��C[�������wz�����`%�1|� ��%�����[j^,0J���v*d'Ꝺ���2�h�ċ�����X�Q�k��/�ţÅ؁���n���0$��T�p���3��b�)&
��ʱ�hf\9�ҫ�:�Ğ
V9uȁ�Z��i��g�rC�h�Gօ�],�r#�9�}����PX-����n�#BI͋Ʀ�к#,�0������g�/��n�X{T�y�#�}�7C������.�Ϙ�)qZU*����H�		H�e%,u��.ȋ� �� �	R��'�ƅ�z���xs������6P��w���u1H�~wO4O>��d��Y�+���O�3+��E��O��:2y����uLWr�8c$v�˯��^T��~mʔk20�P�m	z��II҆M���\v��n��L{�ڛ�@���Z�h�X$��_�ber#(q��BT�p+8�*%��|��hC��i�����S};>ũ�NnO���v��E$��ҧ�6�^4 �2!B!�jE�b�sb�>�`ΗN]�~B>�'@)��Q�c �:�ͅT��T\�&�d�'���,v��Z�ގ�,�'̩l�u�r����7���K�89�p�4AL���W�����r����Ry��׎��#���f�=k��g J[�SB�*��6}��a�;���Ŏ��y�pg���
  ��<�5u���p	p7~�W�2��3��\w�D�0RБ�����q�.�	�CՑbC������6dP0�_.M��J7+�YpMm�e���b��3��j�e��9��]����S�|��FT��¥e�㷌C���E+ol�6=ΪLG8�@LOa���O�o��e������}�&~�Yְ��Q�f��l�~�2�V����sk�I��f'�{X�(��t�ñ���:���T�Oܘh�/�K~W�m�����=��,_a��>�c��H���;�4wj����p�WF� �y�����?L�qɭIX}n���x9�0@��}1&(����X�����E�M3��G��M,�Y�1�Lƀ�*��0VB���wQ�{b8O����_O�#*�{�B�/c�f�"5tJޘ	���v+`m�ă��zL����{��H'�����4"��hU��~���r%}�Ś�;��2�Y?�Ğx,�gLl�����L��:sH����L���V:/3��{�n���5��Lu浩T���6H	��214LS����P�������tvu$��+��r�Uʰ�-U>9�{η�@uJ�v�S�Î=C����xz�1�a�X��3��XEzs~��M��[?���{0��D(�$G�'��ڧ���QrF�����-Z��Դ�p쬘��J?f^�d"�|���l��@�I�?L]vÀ���C�b�U���'KO���Vz�oc.��*L6����"Z���X���&r�t�2B�4��2mwP�T���8B�{�2z�N���M 5������B� X6je��:� ��;h7͵d��_��=��u6G��5R�2#�c��"���v2�  sd�0)_�\�q��ϖ-v�<
�����p��3�[1]O�,��3�W"����G�er��r�k�:���xچ0�8��Y9F��u�I�l�l���P�t����p�-(K."7��N����4(d9ΉIr�wR�����|��^������KI��H�9�-�~E�L�������1G��Fk$]z
fD�;<L�����#b%"���`��]��ꡭ,����'�z�F�.7^T�Ƙ�e��*�P�4�N�H����z[4�U�ӨI�1�]M۲��5��1!s�����Z�{�W��)���h�-���8\�a����a��!:�O⺰_��P� ?Q�S�ϴ~�6J�7*��7?���p֘V~�a�ɲ�n��2�T�\�I�}�(}�Y�-��jb3�S��h����$�1��������ƾh[~*V��I �:}������̄ ��r��)��(���Y��#���̒�5��y�_5Š��Iߎ'�����Ц�i��A��vC^�q��Es5)Ŭ��@V˂���4��//_�����*kɕ�5�k���zC�x=���ې%Y�G$��?/^U������s|j�� � Uz����}�z*�;6r�QF�s�����k4Qb�(�1Ȁ�e��ա��Vھ�/ꄺ�t�X��O߱���z9�6���Rq�3���㐁,qk��C`a�䖡�0���Ч���DƊS�����Yg�rLXy���E͚B1<��E�D�ǿ�h�����O�i� ����Vj��Q�S�3F�mhx�#���l=�:�SgP| 9f;�^Z�d!T��<��ٹ�EKy��7l��	Հ2��0�G��yRt���cK� �_�d��hRH�P�4*;I�D:����W~�Ӟ�gD7D+!������Bd�W4)���%1�7�x}&jp�	���KpRM��	��:5򔊂�4�?�8v�C0x��(o���r�8f����G��P�h���2|�D���ff/�C�u��`��W]w�R�
`#�qS�
	5�G���yt��z�V�P<��|�FP�X~��loV��Ǿ�䫔�PW\y
BT��ì�y^ �/q>VȮ�qx8��O{��;xk�S�yJ��˽o���eb�3t��}yr�,nEZ��Ku�:شI� �j�����omo�{�p����/�j�u�����[��а�ȍ�$��M#c+\5Vп�e��LHD�+hDWm1�YS:�k}A W�
�ߧJ�H�
I�Z�e��RA������b%� ]���Y�fTj��i�6�Ñt������X[*��ޫ��HI��XA�//$���m�gA0�1ݽ�N>oJ���c�|�q%2xU�zՈS�OJ�'�r&}��Ng����c�*�aW���	\�C$È��c+����=Bv6�_�A��m��=ty���9�QL]���<�@c���#<���\�T�:�<�5����Z�E ���R`��W�;�ԓ)��מ��
�	��9���<���I\����`���,�h����ݞ�J�'(o��s���i���V�ϫ��0�נ����K�8�%n"�q��S	�τ�k�Xg\�Z�j�����H�@�/F|K���{�m���!�0ޟŹ�-SVy�y�=;���Y	�V'�YƎ��g�_{`G�,եT� ֪����%�ƞ�,{hn���j� 6�����7����Y����\g`b������Lk��#�Σ�+	ERX,�g�� D0�uX?d|�]��v�����S
�M@z�Z�i��lh�2��C����4����Q��pog*��W�酃MM���?�q��+.�?�yZ�^۽�T -���B1��5k[S���
I�E�փy�F�|�xr��'`��?}Bg��${����27���H���D���O�1\��m�f�r�U6��󫂰B�ވh��x��'z@e��d� �^��A���b��e�[0fԩ�e��`vr~��xaK\��,�� ���#�;>�@�}'Y���ފ��P�A�a[$���|��t��~_�i>M=dڼ++�a	 ��	 ?>�[	�)�C�G��'���x��2�P�{�*2���2?���o��dV���_A�V�ݓ� �]��t���Cޔ�y'L�+��7�P<?h��ơ�\֟u2R�fxq����1(�R��U��t�О)�����oi�\�b�iao8���7% N��Ǥ����� kxGS�ל�[���ZQ�U!�|j�+�l�]�AO�2�)�����{0� �^{���C��b���|�~?����\��,:�_�R��?^w�,���׳�*�<&���oqzR���4����
�Pؼ���I'3����G����C�Q�@�$�Q���'T��ׄq�����(NE~�����A��aer!��X�O�=�`�FՋ35�'8���?��t��oL��H�雿��2�v~��x:������b[C�IG��" =	��~���M���� ���H'�,o��d��B��Scx�onl#�w20M7� ǛY��)˦8|��΍��4V*]��q昙��9O�g���J�f�A���ᚕV�o��Y���H��8��QJ/��_F�D]��i)�k�Į"^ U
�åB�B�T���������#�F��O����������1i���X����R䣠����/�wI�DR\�v5��q?�c�$Y���^t'�~����`�WIA��mL���b~�m�L�רu8�&��8��I`��~y�Nwo�Y��O_*br���V�>���:r�q0X��3�+�J��]�H���p�s&3c��%��Ǡ�a��߾������X�+(Iϸ+Q�?՛Z�7���"���7�����XR'!n��^�����^��"B#~AY����侰ޞhBFM��ͳ�\���_��Iz��s�$ ��y�@<5f#�T�{�|_;�A�vﾄL�'C��x);p�_�C���<�)��/�t� vޕk����ˌ��JF���-���!ѲP��?��ٽ����o�&����l5 wg[�,Vx���2÷�c���n�޵�����X�B^��+~�����z����X��U����Dn���܄��",�+ti	���������ܞ�@&1��@���������+������icG��M��b���mИ0%��|��pmC��+#%)|��6�-6aB��F��I�BR��W��p�dk9�Z����n��iTnG�"嶑�7�_�'=wl�IS���;�T��Hp����}��~�Q��?�`�	�W��݁%'J�D����˟[�MO�(��R���c���-��!�� �F�Md:)5���>`��B�z�R����˯����)C!9~�GǷ��m+��B�ԙ>�^a�O������/נs�8te�8O�J�"/��@���;���R��pgH;c!�;����� %�{�y9!����p84�^�_�"s��}�o�uF
Nf�y���Uձ���?ɔ{ �OQn��r��ѡ��.y��3N�A��/��{҆�p�}[���ZG\nЏ���y�H�-ጼ:S&Tǹ�ߏo��ڴ���Wd��^�^�����龯P�� �Bk�1���Y�\	5YL{�� 
�{�bhg�����\�B=9����^�\�t�%�y�n�LX�;�aj��g����H׾�H���|�0�OYaUKV-�ÐC䇯�j8/��Ԗ�Ul@�W�;�L�9�+�⋪��gI��+,S�#���I��3��"��H�>j\�SBV��o��:C5�
	�ޡ�����y�$ZCm�ϰ��^:��yC��D0_T �##��+�� " ~~p��X���l���h���L�Ծ1/G6�gR�,�V0��"�JI ,�喝�M"E�³���j�P&�!���_!mƧb	�O����q`Y_\G� ��b���6����*ay�K+C����z&꫌5|d�Mo'�u�����>�c�>�I�a��J����ju�E�X@���ga�'L[�d�E�٠��HA]'�hf�%F�/�2��}�
Ÿ�{�s�-�����߹ˎ	}
j���
9�A��(�~M�B���φǈ3 ��hD�ܵk�E���!@3��'�s�nDO��wP�͉UGݶe�F@��d������;�iq̄V�V��-,�݋�1�a�ػ�Vo�$�	�XY��ϰ�2_���e\%Z�(��k�Z�\��y��>{n����\��,I��6 ˂7�~�H���R�� ������;��=������ޟ8��_��CL���gSҶ~��?�V V� ��Ż��F��r:)Jv�0K�j�~C{;�&�j���׏i��g�J͎[R���@m��a�ؿ�!RT�z����m��3b�*�
��%�w��\���peuhAMz���\xn�J>j�,! �^~U���+����;+6+���o��7��P K.�_n�,�Gc�å��Ɣ��f�r�����8�"�v[���X����Y��w��O����8���_HH��ˬ�\f�'�8ŹW׬n��&}���"l�����d>���.�v�\�]̷���?:
6O�����sL�d��P��16�0�� NtT]3Ik�0�Vw��ַ��MHBrZA�..�_������G)�ȶ/!U���\Z��`�O�8�5�'����r8>Y�K���q�����������'�n�b�K��Ú�'`�G/�,  ���#|�}��=ڂ��8�!�=,P�L�|Y�1W� ��G8���;Y����Tu����E��� ȋ�~[�5��A�kӢ	��J�`�(������;�H�e��ӡ�V�b�9�d �J�8h�
�y�����EJa~v7���3���DmĄ�im_�,�/�+����u�nf�o,�8ۿ�B���:��uj��nGB}��-ѸRx.���k�ZsS~ٲ����j$VO+���+e���be�\��$y�J�zWs4����m?��1Jpx��$�ɽ:1��:�k�\��,c���I2D�g	n�V)0���_��C�Ud�� �̾՗�M��I�+nK1�[��W~1^��'xb#(�xF@5.;�X����O �ֺԞ{���'A���/�A��[׽���b@$B�t6��Od���"+�-��I��!x�+1
y�$�7FB�j+��d/�[�& L���Y��)[�)�H
d2��;��F��Y���1��
_�����)��-'X�O.����c m¬e�A�Us�!��!9o6��^��pľ��#�	��:��+DhO����2%�2I��%���oj�Cu�Na2�;)���䛂ߦyDm�J*�Ŷ�G?���h�:��3���Ш��mɺ��� �G۪/�`����.c ���C[yf��S�Zf�x�p�s����BJ�]�4��eٺ��1�0��}��`f�P|i�'$�Tf?�S���(/&�Hڼ^�H�#�[�}��>�*��5m�G����Ğ��x@ O�I���*;/�e�ٸ[&E+�j}��0c��U��"rp֚c��q�y�H~�t�Wڞ���O�%9�M[2���_�`�*G��O���μ�炬�U����8=f��|D���5��.fl��}�yà�i�q�w?A	�3��k��8�|Ԃ@���bE�����F�D��V!䤮b%��LY4T{�w�Rm�uB�yQ_?C�.�	F=6H�3��A��<G�1�QK�Z���)���Qϊ�j��~7%��bk�8�ܿw�	��[�-'W��֯�S;; <�鬉O*=�'.���&|^�r^N��c�ᇁN⧕ĕ�AS�ҟ�Q���S��ķQZjGH湷nr_�Y�΂�r�gFp()��Zڴ�V��զ��嗽��h��qư-���;��?�#� 6/5�V�1�h9�;�:}M����Z�F�����8�KS�B��J�}%�&���eIC7��AT͸��;O��^h3�e��ݓ�� ��h��✨a��$%G�A�E�<qۃ����x�&� 0�5�M���4g�[��\)^����@�D�:.��ٔ�&�!|�|{���lOz�E8!���t5�Qc^P֒�d��/&�/c���j
O*2F�o�[�8�-�n�˘RL��V�����9����7Y��2��	�Ϸ���/n�X�ʈiv�Ty������LYV����ԥ*�r��$�ՠ��%�={>��Nty���6��Ɨ-s��`z����P=k�h����w\��v��pX�UR��҇�4�#P�e-j�N
�A�l{��˰��e�[�V���`���7ړ��*�����E�d��q�sq(�S�}n��|\G'���<ߐʂ�������oT��t}IA�������b�pk��Ⓔ=I7?$�7�I�M.��x�n$������P�K#���Jfҷ��G�������C-T�6uh�F�E�,���i0���b������S�:\�ˮ��B�����E��aՆ䠹m\ ��͈�"Лj���;o4ˉ�o:!�N'�h˷:H��)7u���_�"İ:��@����XJ��9�T��B��h���6e23^��,�:���͑�`K:��p�4&Qj�dj���ŏ`8y2Y�����a^R�R�Zb>�G] 3�E���Ϸ8����7:�l��xz��Go�@бO��LA/���`�������01s$�7�u��œ����q��s�_K��ȇ�=��\����u�q��+ld%�<��5�^��,/s� XdK�~��"k��wx\.{R���otq"�;��#G�+��}����x�B@y��$Q��M)�>$�m���N��(w:���6|��R9"����L�BAJ�To�H;�$tJ�m�^��A&�]�:����H!�K�Q��vύ�g0%�;
���&��4�����Y����h�����/Oop��cU�z��L��K��e%�Ȑ�=-Z=@)��s\��R'��~��tT�ֺ.Q��>G�v9�b���HN�^Ԗ����{=3��Ġ�N���K,��>����/Ɓ�)�`+�M>~_Q��k���`- DO��;��f�.���Ӑ��cuF�O[}1�} ̲o^�v1"$�Z���hB�ڳ�$b�/��+�N�{��b�~����8� �̙���iL�-w u3��ׂu b1:@m�W�'G�i��|�w��Bo�1<�ٱp�qӳ{A��[R�;�|;L�)�	\�2�ɤ���������$pJ2�p��>��_h681V�7��S{<L�&F3H�y��w�#����*:&(<E++���˳Ѱ� %���c{�O,5� � 	>�~hȪ�k��zO���+�Y1ڂ���O��T�����x6]=�
�A4C�Ҿ<������*��������8b���m;%��rn,�s��;[z��1�����uG��]���OU�Y�R�}�G눡vZ��ɩ��.���~ G�3��X�K�O��y;��X�Р$3tX�.f{c%�n0��0A��lz�I`@�jA��#���,>�
п1L÷����l�ڌ�&��pfD�A�R��Q�����|�;���B�7T�ܒL24��\(�$[���tLr2)�����%T�(�j◆N#.�0�N�͹�������� 9e�i����w8����b?m�Y�n�[�T�Q�m�&쯁X�p������{��4���������6}j�M|�>t4���~�����]_Mte�E��wI�iS&��k�,�3@"�_��}��(���as�08-5)4��r�ޡ1>"��Z�T�Py���ڠ�w��Z,8I�L�+W����Q��5���a���d��ؿ�q��C@,� /�a��q�S��:;z��ɣLm��6�fO\$D�2��p�)�c���t�pͷkk1I5�g�	�r2ѮFzhR�jA6�E!/ɒ�+��Mg�		J�G��.�~EIa�5�~ˀdvz�6��YP3gn8/��B�o
�K<m$��f�Q��i��\,dZ\����}���i�����A9�S^]4�֓���l�bbq������oV��zI����E�Ӭq������-o�r�d���D���۟�Lr�FXF`@�P�*�j��������>+�ϣނN.��vb�P$��L-b�D�([/xb�\`��F[����@���"қ��G�$:���/[�q�����4nyΈE�h��-/ء��\��,��VvK]C��f.$qD�_�J1ô?R�[�^����&Qs�޷��_5L��~�dU��Ib�G��*�v<����Ȫ6�&�2ksb�sUI��9\�`�:Ѽ���'a�����M�L/'l�ޔfp���hcyp��&̗��el���_���,�VSXʈg
�� �s��f��䁥$��3tX�6������ϯ��n]�d��	8����
]�D�Ht:�I�j7�Z}�����p�_�EO���ʔ��/�:���p��+/Q~�ܲ��R���a~Tm՝i��=��:�k�C��\����u��_F�o���^����}��[Aiw���xӃ�� �f$�-�7mN?M�J=�U��\b�0��Kj����kC�2�N^�%���:�;����'�W�����Uu?R<~��_��#��*�t��ߑ�Qc��R���v坭�����DMC��6�%�5��e(��3�ebLo]~��D�_��%|�̓T&ng��:\� Sv�����?�)��b/s�b���>�3 |��N7���=C8�'��a7b(��c��B	O,��e���d�~�t*6r�q�N�|��Sƾ�����9��gB��le�!
����,�"�;��W���q�Y����׮���c�;x��x=d�$>��Ns�O���m�T��=65��� 3TV��֫�Tų� �"�=+&C�Nڹ���]��?x�ۡ{�W�:�8?O�:K ��V�@?���n�w��v~:���Aᔍ�%���J�ci�P��WHd�j�"������,Q7�����Z}��t����:��܈o}���B{��~/ؗ��vV��>�c�6'�G�8�ƴ )��E�왟.z%ED�2؉��9>�g��'��Bĕ��v#t�L�^,����I�Qv~f�D2$އs2�.�Pwεo&AN��v���\�5<��I,�	W�ּL�/�Y�{�C�R6{�uˀ��b3�S��i=uA�i�3�-<rBtq�O�)��j�:دzּi�<;�E[�V����j������������#����p�+7l�z���������������ݠu��i�n�1fm��㡍��P~)c.��Z7�]Ņ�#�\O�Wu�5ڭ-��S5�PD�eӨ�2�������H�q�ek ��.3J���?f��&����A�#�o�dT�"T���XeV�Wv��0��.��"�I�ahHH��%��*Y3��<��\�eh+`�';�A|A��
)�0xv�"*�RK��G���c�t���zJ�%���B�!em�f��1('@)�E85$~��|6��5�������r�x&�&����D!�ew@��L��d�c9`3'YS�>&Q�d��w�h�Y�{���}�2����-R�ȩ���*���;K�;OѐYy�fD1��B=3K�	��q,�����wT�s@�\-�~Z�oR��A�
���;4.��nU�p�9��U?�:�R��rܑ�y�P�L	5���8����k�L1n�FZ�~��1�Ͽe�PH�V�_�3�O��K���N���3�6<R�Y5� ��a.(��Ec�ӝ��1}K���Jl��oPw����������:ڥ��S�2Ux��Z�$��qAt��$�3z�o������y��-ۜ�$(�/	1X	|㢉<��l�RP�J ���8"	���o���%���#�b�&�B�P�m��eӅ�*�J���������E��<w�i����N<��E�3k5t+4r�h����L�|�yy���I�Iv�R�\�ǖo�I����/QR��zR�z��U`�b:�NܮI툧h=�z�چxJײ��!b�J�?>�R𡚽�JD c��V~cm�igE(�*��X�"ҠB��i\������ ���c(<�������6�&������wW����B:�s�c\;���cEy����"�&��a"��\�Q=~kr���ݥ���oᱨ̱��Aj��({b�J�kť�B,7�W�F�_,�
Ԣ�V3Z��'�y@	  �Kl�(:�]+!��N�j�;Խ p��"��´�;X
�1Ʃ��&6��TM	w��tg)N���qS�o�wn&dg��_��x�!H��"'u�(��?Q�p���Вk����x��j�
3"��9�?k[�0���*���?��8�sc��Dm�8 Ʒ����6��.a�D�g,a&�V�S�8��:�4���IΛ�_R�n�����J"�Ҁ�dɓ������	�*
`�ow+�9��I&%,lųe-���&���{��O@��P,TL�8�&g�������xc,0��Ģ	�;h��lS����Ђ�5<G �F�+1>��i3��U��7��Lm5�(�8cQR�V�=E����n�46��K��Ȱ�c�A��-V~�q�n��|�&�K���n $m�J��4��y���dD߉b$=G
�1�����aO�#������,@^P�sMj���3ױ ��z�C@ș�.�{Ԟ�Ҋa��N삕�~οpI��`�i�ݥ,M��)��Y4�Zz_��uO���-&�$� t�"^��Y��Wd}h��zj�]U_�F�ړ�jW{�5/�!K+8���g2�R�5�%�e&������,��ّ�	��BK��s##�fJƴ~*�� �0K��X������Y$g��YP[ZH����	-����m-���-�i���m�:q�`����yȫ9�;$x.+��f�f;�����*���0�F�Zd��+A�s�e�.XPS3H�8򺏬t^0��	��������9��o�4K����7���A����hϫ�������pi�Z�(��f�j})�q~@-Q��H����E!Q�>��nʂ��zK/�NJJ��8��l�]��9�i�����~Oޅo�^����AcϏ�r���_� Ң��y�8��R�5/���/~��hf���.X4�Fy�½�o3}B�52�뵓��k��4Q�L����	�ZYҥ�P��q�5���a���U܂�j�t��Ä��s>Җ���H��!�����'!!	:tV6'̩�hp+V#��%$��~��|@p��v��x����GE�z/�[����5�j�Z��H)�À!�28K9��{q�R>��}W��dݬ)Z��}�2_�d{�$t�����"r;Z˵E,2>z]d[�,�پ�P;J{�GK̵0{ԭTl@�.�2��ݡ>&��P��	O!�P�R��z`�Ԫ����Ol-�qϙ�wƳ;��#9�,�^N=�=���{s'3��q<'���y��O.�(ₒ�j���6%䋯;��S�Z�ܚqR&�7��sYA"D�j�WظP�I힨/��U� �u|�L�`�[�X�0Q�0,w� �45�K��:oʵ�2I�Y2*I����z��V�f�IJΥ�I��_!����W�
,�Cc�xŇTN��d7w���t-�r�:x�3��"��(�����a����Qvpti��3���5���U#��3'�R�j�܄���Ƅ�!v���{���s�(;�⩆Ɏ1�>�q�ߋi��jީ�j�ȉ��7itH$�QK.;����v�|V�itL�w@��1�r\r}��}q��<��*������kJv]���c ��f�b�/�7O��c�P��[�mLp��35V �>���4TZZP�C�d���e�<�G�5���+�W>QD��*��+��˂��S���_K
V�����B����b���y�U,�q۷~v��8p��������y,�|���%� Wj/�R'�P��t�vX�p&o?9 o3|4v*�jW�_5/�T (W~\G����j�Ϣ�p/���5!A�6qO��K�~��Ap�d[,��K'H�aD
�ak��m1�Lx���$���ӧ���M&�uMU�F�o���<k����
�1��0��G�P��;]yd#x�IZ�34���먏9�C��	"��]�ӱS#=T��;y�5��o���8��y��뽎��;�=!�s�"jiX���%VT"n?ɿj��[���P�7�����8�F(d3:�gK��my���@�H��=�3�#o0�Cӹ���J&G+X�~3�p��z��d�q̕U��a�F����dq����U�b���7)E>7L�w����8���S�t�R@��\��a�dآ�P���M3H��+K��u�+���[���,�	���u�!�Y�rO_3�}J�-����s�i��Z{�t?;����E:� �@������GO���!g��;0"��Q6T���@��]���]�k��Tzemݧ�����)��i+B;����<r�Z�p�E�~�0�Z]�<y� ���7��f�|^X�hYA鯞lh�������:Euc���y�ҽ����6OZq{��������K$V��0��(��LA/���oP�H���Զ����JG��^l��'Y4i��a��v���cw���8�+�@���x�_�~��#C�}�bj���w
�{��2˰$�`K{���OF\+������X��#Wp��z��$Y�Yh�}��֖z}
fq��X�w��]"�>��^���^~׆���Pg�$]�x�Ld�7ֳF8n��H5�rX��F�x�R��fh�*{�Qg��#����؞�e�ѹ��/"ߣ�3��%-��5�T�3�������6|�R�b�k��I!6���9&#JZ����BMXf7J�d���y/륛h �����ar�"�97T^R}Dg���.2YI~��I��� t�0@��� �x�>�ND��e��B
��G��jG��G�C��r_a�h�(k��	KQ��0@�WV�A�d�:rjt�Z��$����ؐ} $3�9�u5v�\W�핑5�`��l��VKr�y� ���hCJ}ZL��˭�3���ePՀ�A�TP��]�!�ҁŅ1�wm玒��p������7�po-6��6q޻���a?I�M��Ff��q�"tP�O"B|��t�R�pFۄA�����GRm:�:�R�kdww��`d:w�L�^�fs���4���kW�z��x'¢�_cPkæ.�#/��mP�b5o�����.�����R5�ۇ��ّ*��F����߸4���7h1����b'E�)�t���F��&Z2��q�5�m�37A�)�2�]�f��GR��m+�hH��v^��9Y��ut{Z��nzq�j�3��w?shK=)dv�M(B@b~j��m�l�K&������7W�_�%�`��uCށgA�2s�~:�x��lv��A+�m~5W����<�-�N�&��3��Ѫq���ʪd�'�X�U�����Ab��zˋM��v͘T�1��M�Qy�=0J��r���n�Wm=|F�j)7bb�s;��eb�py�j�����p�#tY27m����j�}�3�v'>H�����A1��S������I��:�v���� ��6��˪n���/V��27�2�"F�oPB3,#�.�]p�6�k� �̝�;��2��P���9��2�C '��:"Z!e��3� �Q�ґ����e���a���M` uaiTwB p�HV����y��<��z�� �q�I@lL�u��/���7t�������t�+0�<�{��l��Z4R��~n%R#vt�
�����Ѹ��m�f�q^����:��W�tU��m/��Cn4�ԡu�3O��K=���c��^1�,Ci����3~���-�<<���Le�*�v==�KK��~�u��]���a�@PJ�����ˏe���=���$�7qI�⥡*�`	��ۨ*�~x'+�UH�o��C���7�Y�t��b�YW�bC��:9�gڭY��n�30�v���;-�u������}8�Q���0@s:�������5�j�z{Ĥ�+� �刔	Mj��������r5���Іэ���#wzc\�C�0���'R8�m]:K�1d��L���Z|#?�#p����\��"OX]��;���柙E��
�}i�`�F샘�E�~��B[oF���觩i�Z�J��ほ�.�*K�|h4� 
w*�)�@	W�  )J�t>AU�s�(H�A�J�̜�2p)�!R ��:�6g]q+��:gdbp9L:����]�zI�Ȯ慟r5���9c������gz7�+�����vx���$A�"LSl�_FgC~�{�km��������4���M�+R�%A~ezN�>�C�pج��y�����,��\'R>����=�z��ĸ����<Cι��4X�MF���Q/H�ﺫ<�xEI��(I��TaD��zу��cW�C����$�3-���Njt�H��2p�����&[���J�_��}���=/s���d/��S�v͸�w>��Br��'z��
�(�3���Ƙ���������b�2�j ��n����n�Pȥ��xڌ�J���
�7#8�5��й�!:_�3S��O.-��	��ݿ�<�|yh�a�jW�1�gꕴ�D���.������h�;|e��EH6��Q�h�F?�`��m��Y�O��;aY�ϗL;5<��5������A��~
� Mu���6@ժpU,))6�Ȩ.,C2�܏鏜�ж���Ub�X�E���1
ǹ;Ƿe��$�L�m[5�N,B�ݤP���u��_[��Y�����k�yI,�}M����uIv���U1����p�s�:����u�/����mY��?��bW�?�!у	����U
���7�Կ^n�����E����뭺m�@�<Gg[1_���$���?�+cB<}�׊�P����,�HV�9T(�����*�f��&�C�߲	�}85R�54����1���==���Iɿ�s$��EWp6V܃4KZ�}��d�@�r�������^��Ī%��B�^�R�B�RWH�+p��}�N}�b>�r�=��r�6"ة4�ݙ�5��wQm�bS��n��m�X��n��a�J%�T1���R*��mb�<�b�T��ƌ�(Lv���j|�k�E�G��$d}��)�QOtX�|8�<��h��N>��$P@�2�x^�Z�#p�:����&�貏�|%������d�w�����C[�:���[M�X�4�	�r�f������m��e�3����d�^��d�\\���_E����+��e6r���(6Xo�E��3��K�tgL��4b<�z�+\��8�v# ���H����������V��G����Ƀ/eY�