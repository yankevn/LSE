��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�U�|�=���Bk:��;'8�l@���kx�V����&2b	D��t��Z��Ex��v�t�R3+�̊��Ls��]�Wv~��a�MG@g��mVF2�L�޼M_k�oK.fHG'/���Q�9���[�
�����mN�5!\lwL4��(����x��`$�c�0<�,!t
�M����b��*h��9 ��!M���k΂�T�����Z-p����D���G7�t)�ړ��q���3 {e��L�T1���]���l���:q���"w;
РCS؂�&w����7$�D0��@{�qr���y��t�va����ή[�����:ʼ�z�̦����W���`0�M�'�,>!��**�[CC(Z��$(Z%6��BZ#����A�\���g	
|F�ܖ��2�<������T�@�|�E���3�`KH62K���㭾����$L"VTXo��KZ7��m��\�9��GJw[z׷k�{��p��׎�(��C�R���1���Ug���ķ�5i� F�'B�	��%���DjY�}k�,�M?�o���E&)���!��ȱ�LF�����ߩ�ܷ���w�����u�(Z޼l�75���"a���q��� �^K�d�Q�]��K�RԴ2ə�F6�y=�%�&��X�����3����_W��ᶧ!a���7�-�΄3=Vm'[~�iB�Z��y�o}���\$�j���F�ͪ��@g�X]����		T�O�y��`#%��!Ce�Unn}~f�?:���B��Z@Sn�c4��P�1u�ե�d�ogy��d�m�x�~�v3�?f�W*Xe>��%u�Եw��PfJt�����=�]��zg;�G����Z���G��L�E�햋7�� ��L'j1+�x`D3�Ž@�E��=!��ʏ.�D=d'�9���U��������{u̩B�1���^T�r������	�%�l��6蹫
�Z�m��|!��R쫽I6��hf�ni�9���*���E�n޵Н�6�@���n�"B�_�XZ�gc�C}a�٘\�y��~��		����u�''���>Ë����>�-FA����]m+���o��t�=��J��k�H:(=d���V�B�R2��a��=�᭛�1ܾL�IٿZ�<�L�e�\*-P5k;r�:�������h# �)�S��/���X
�hZO���[��|hu��nN+XSW�Ǘq��t@Q p1�ʬ�0��oK6�u�#ԕ��9�Y���F}�-�y6OU&V�r�9��ZC��=�<KսV�;�����M��O��\��Ĩ�;ڒ�R�R@��a���!B��JJͶ�O�������B��RL�]Rֽ&o�U��#-Dn8�6ո�J�MΤ0M=�|��l3?��am���V02us��}t���1���O�m�����U�w��5�MeS�Ì%�!��"�upb~^���[���^�
����m��Ȳ���/�x-Q@�h$-��*8���D 0�eoJ,`��K��s��ʫ<Cp�����E�>n��������=k�^���=���}Uu�0�<^/�7� �5t<p�.q��.��ic��ס�$#m�\ۦBe��v�Z�����D���˜vTd��^�{HF�p��%�r@]�����z�����[�Ĕ���s���
u��i��dUug�=-�� zφ�g��ō�Nm���ٝí�tdȽ��Ǎ&�Κ����F��\�<�_w'�]����+��ԉ�j�r�K5�{�JQ?�e֚#7�:�_;�s������DW��꿹���^DX�uEgF�7��,����֠\z暡�����L0>�~�/^v����Tz�J X�y��f	<�yi��j�&�M�~��* \��V����c�Ⱥ@4�姯�lU�������)<R_nשQ���B���O5;��,{m`K���oXS�P���DÊޒO���9��nc�:K0�h�5���\�]��׸�i��w1������Ӱ��=�]���~4��Ў��>Bq	{���@{
���f��͊;'�6�B<�b܃D��nҍ��)4����va���@��E�M??���W�0�Z�)�ղL{&�c�c��UD�� �޻��*�}^�H��zJt��?鱟L����M�k��}&��<��&�6���"���6BC/]�?p�7�Y���$�D�<�}�_�q��"�q�;�an9����E�}?�=T�e�I|a��p/���?�l ���Z�y��O�d�I����17�h���$� ��f+�q��� �4�IH� c�	�y~����[��ǡÇIjKq�F3}T�ᙅ]����ٜ�
�Q�c�6�ew�T�H���PV���K���׊̋��DQ�[]��W����m�>��~fj#��~��!���u\�HF5��U�z���u%��KL�|��w%���װď��|�˳T�x�"��-Rnp�&2-��k�7Qx��v���B����=*��࡬}X����;{u�
��v�Jc�����/�7	i�ge����<�2885�Fу;��su�mK�*��6��8J�b��[k�Y�iK�/��
-��<�1��{g�\��7�n?%8�V��eU��|'	�,�w��g*h|+��+fZ"H�
�ې��j-LW<��!�o��˹aU�������pf�r#�mHT�Ĉ���T�ޖ�M���,�f�[�S���s�}�Z��� +,ת�gQ���T=�kL���� D��S2;����&n� �6�:� �_
/�4��@kNX����2���T>���	����gd�-'��s��k�G����K�+�%������=#,�i7�j-*��3�Y���C=Y��]C:���{�H���L�Gg5s|�L0,b�z�7߰���.�}h��YG�I�&%h�s;>uh/�T3\y��s3Al�#�3���W��B�5���=	`��0,NL�AmGL';�$`*��ߠB�A�����z	f��7Z���&1
�%R�$ʵѷ��y.����CG�-ڗk�$�F��!�=�IM_3厎R�;�w׆�g�(��Ί��2K��6���4�������W��Ɋ6-U@�H�������,۲𢸖h�.L��D�H)��H旸����ث
�7OS���g���]�ȹ����[�C�)�vρ4�T�KK�U�a��L8l�9b�p���>[8,M{�����w�UIF��� �z��u�+A%}#���%�;,ǲx�Y�%��͡]�χ}=��,�X����$�\��cs��"�0�UmQ�ºVN��Ռhw
@���|�c���R~�_;�Li�2�'�ڡ.�����7p�ymr����v[ئ���2&��5���sP��/����}� ��-v*��e�I�{sq��}#V�2�P!b�w�t�gaD���ɿ���7�� *��b,E��u�7tg*Υl���},_�*\������PD��'S��n~a_��c>�YWb�xu���㧢�I�	Jwyo�������Z���6a�|�{%[M(���xF���C>l�-~�I���9wm��h�'x�^�"��*�.�ק���	����0`ӽUS�X� 轠[�P/4��F�7	��&��r�_����W�-fK5
��9���ChP�p�Փ=���4�����N�������uБ§h��S�"�	1��� ����LLn�ֲ詷Ce_
�Y�U��-I[��kC�4;)"���1���\/e�?K�3�Sںg2��jW�.��DI�J
�롥'�0�Đ�����oI��,P���Ao3��Y*ŞTL+;�Ge�+�J�����o4�cf���Il�H/\M�pL�Ǎŀ �$�{�k)��DD,���)X��d���'���&"��g�i��!�SšM	I�f�ƪ��/�v%�-4�s=��=~�fJ�%lݥ8����d������W��i�&w��d�����n�.��vG�JQ��:�"xzo�y��}h�9�*^�4�'��F�k�h�0��~=r���19��F�MA��QЂyw١�����߱�q+��`-�K�ĈU^1�o�उ)�˪����cy�~Y�ȝ��} ��n��f��Nרּ���I\�P0��-�IX�Y��j�t��Y1v��V��w�0��{��$�=���$�8�p\���<qڭ��Dɞ#yMg��nG��v��ȍ�$ p�� �庐�pyrUSD��,�dýQ�m�Q'���PN��Kp��:x�/�Dj���*Ak�?�����D��RH09�LT�=����Xn�d6��kf^U$V"	�Uzfԗ?P���oƽ�C�	���޺`�D�M�+�Sr$�Y��1\��;��!(���f�0���� 0�o���;�^4��j�3�uv-���w$�������	�Y����l ����F2������0�Z��M\�s
[�����s��s���s
��#���6�������6�u���0eN���w�e�Ѽ��ﱮ�`n�v�5�'��-m��
�Y�"Å<��n�E�!�Q$��ޮE�1^��|��zbO�K�Wʜ_��X�'ڙH[��vG��Z���_]>�z�6P��ɇ�>����jQ!�.N�7s��p�d�=&�W�z�ՙB��R��	S�x�Z�d]#���
[�T~e��3�_�^����LY�����2�� d��!��6<�)�Dy��6�8w��7�ʛ�u���˞�2�D�� ���}'y�$p~�RFa
엶 >�}]��e���p�}�L0��TY��5@�����R���4{���������+������?ftټ&-�A+I�BOc���I�4+@��`���|���6��)�:.ɿ����M3��[��읝K�AL��X��fs����yF�[e�1[�v=�<��~��8Ѣ��O��6[8ڧ��$��>]->c1�]��ΐz��
d���e����P7�~�2�c�>�bs�8�kY<9��][!Z�(��l�ޒ^k����R�q/�hbb<��v�"W��`l��n�p]֟<u���L�m�X���0xY��T��t]��V���]NȆ�1
���}����-��`��3�q���Y�@��(��[�aU�'��:�Yi��i�ubc�+i�����l����,ݼ�K]"��iD��EK�/=+|���W	;{T=�8���4�l���؊_�n�[D13\��G$���;���f/
���P���E:@&�	��'uYq�,E��'c����9��am�]w�~Nq
$9��<W�(��H��o!g�-��1�6��_V�*h)F�Z���E���u�i�EQ��µA��R���> ���:�}E�<<:&��¼�b��U��K��,�I`L�h��}��7�."��8�!� ��#����
b�?-�ZP����V�]̪h���[�Bz����w"X��t��*\����E�i+�����
�G��Xk
���$��s�Q?�y�<�����?X�:�k��D ��h�ؠ?d=��@����&��t�����6k�ŝE�|5�vh���^���Y*�.P�)��v��8�1M�A�y��w�-`�X�7�r�Q�7?��i�?[�Q�"��[�ͣ��+���Z�g17��m�a�)����X@R��X��LH�2���M�!���(���>�Vt�oyƐ�ͫ���$ $�`\;{5��1kk�����b2�^*s!�+sBvx���8}^����{�2����1
ܖ�>/��d�?B(��	��,
��dk��c� �xK��	�®R?���y4^�-�P��P7�8�j�<*9�Q~$ur��rBi�n����N���Ac-8?j��G��חb�'�7}�Լj���S+Tsҝ�����RF�\J57d����E}�.s�q��Sħ%�v�Q���HZ�j|�Bgs� @x�!�U��;�lF�:�u:���)�-`ݗ�_A6�
C%p�Yr�
�L���l2�޹��ܜ�
�'Tyn���� C�)j���<!�c%KI�A��m~ܮ��*x(�ЭѸ�%�/�ٓ�_B.�*"�s�|\�d���Y���3�gl���rT���vB�un������6Ŭ�$�`�����YO�Ϳ|�xK�����7h��@MO�G�����	g����Y{�m&��d�(����j�ݚ�q�����������م91�� ��:U�оp���a'B�#o$Ŀ�F6�����g$�O!o�VoN����湻g���?un�b%#�D�I��$�d��=������W�����O�K����A�-�EJ�QǍ��R��P�����k�9_duqАַ���C�l(_;~�����'���&.��K��P�à�-9}z>i�{��\�<ʰ���od�)-ߕY�~b��ɡ�\����!�5)��dx�8�6�w��C�3�֩��ۭ��$xP=m��QbѢ߱!��>�gS1a}Ա� �j��!��
����֑��yn���7�rjW�� [gB9���dH�`FFO`���k��il�>63zƈG5u�25|z�ǎc�*q!�FV���Q*�x&]�AB�a3��ƘR�F8bf�9�a�-d�%/<���MAG�]ǉ��.Ds�s�[�I�ڋ�i���5�"Q�@�UN�B�{�������]%pU��-���f
�g��N�*����
X~Ǉut�4Ocu�*��:6æ֛2�ߚ|���Q�$�a�2�g�ȈМ�픢@��.���L.��܀mH+�UJqĽԣ"�R1��w�Z�x�mP�WIQ��֫!P!!x´$@H�ɑ ��	�_s+&�!y��rN���ɧH�D���kL�E�5���i6]¨D�@���jZ�-7nn0�~�v/+�����P�γ(�θR�cp�Hu��IAg�4-9y6C��౺�}�9�`s<VS����z)l�/��:y�l$�U��[�;�\���""��I��ѶN�˘X�l���$shy]�6ُ�L"�n���M�T�E��7L�E���cp�+�ǟ���K�H�n�ay�Oi�%*>OH���.�'N$S"��w����.�0L��V���&��v`k�h�S"���F�l�jMe��@3�*�/������p3����������m!��C^�K|��A�#�`�[���s��Rr�u=�DaJbz�uRͶ�[���`E{RKl���VWVuлZQ�7.�NDnE��t�c�qa6�c�!��`�Z�+���?���j�9o�:@7˹µ���}v���.��g����7��)y�q](�vpj�����/Z}>�P����# �/�1��p�Y
Ç4wY����=\'��vo����"SXͲ3�/��HȤ�[���/���3���h�Sb��"�t?嬯�9�'�i��3�q5㉃��_S�x���9���5zN0�5����gna�s��7Ye0@�`h긾��s��k>hlZ{�#����u�A�����-���^t�k����a��P.o�}�����/���1� �`M�_Z�?�4R���{�ٿcـK�or�#�*��G�� ��v(xË�� חy��<_,��R2��8a�!�K��׾h�1��SsX��MB؅���% ���W��G�/g��.a�HǶaD/��(��@}�C7�O�t�Ss3|9wZn�"tѸ`:PAh ��NW+R�w������ǻ������b�I,�[W��3�3��!J9ؤ�a|Z��˨)b�e'��PYf�dT��>�T�;r����8�6�SJ�?�c[P����j��$?r�d���0���!+�r .Φ�v?��c��#,[�D�m����{K�1���L�=��y�0z�Idh��f���^��M>ɝ��t�kN��X-(�Ǭe����L�^�Bd~?�1�?Ag�C2��Y��\�������J�=/�ӌSA��|��Ф���-w^Xz��J��AӃ�[�i^O��+67Z�j�A^��C��cg�R���{����v�z8d\����@��.���i��Qd��n��כɳ����y�[�da��C("�bS!�"yأ ���T��t��7 :�?��� �C���L���Tɴ�ρ����]��a��Q�q펃�J��*G�f�����3��Ęb�c��2IV<�X��J�b2p����
d^ڄ�힏ȬzX$��R�l��t L$L�Fm��{D��(R�;��T�꣋���_4PH�h[�;A�H��9�0D�e��Z��ӧ(tJ�6{��+"�Y�k1��,�s���ǀ��k
�TK�ʟe���>��� �&]l}lp��9m�髉SI���
uт���e��^�ԡ�˂Hv���k�^��ŕ�
 樖���ɽ�
��xӓw^`*$��\זl�4����f�T���ޖ'rX_����2X|��dwY�j����fc�9$`aJ�:�xMgZy`��\4)G���T@[���瞑�i%p�ec�#os�;*h�-��g�@+�qGa͚���r�7�V_c�{3D��0Iʡ���6Y��N7�7�U��ź-8��X=���!�.��Y ���}7��:�_�*�q��"~�t'�{BWN�C��!_��C���\C�E¼W͘�z��G���[���G���BA�> ��T����Xi��lf��|D�*z�WN��$�Ȟ�� |�dg��7ح�Ej�Z5�T��+\(Qʰy����S߳���(vJzYq��a�W�._&=��L(��u��|�M�;�^Ҥ����ts���N����U�u����=F���ދ����OJ��Q�5���X6��Vl�2�2���>�
���.�4R�����d�E�['���f�C�dJ�:����Z����b�Q�aa�����Ӳ��:�@�p,��T1S0��'_l���ѱ�͌@
K|fo��%�
���vJ�)�p5�:$T�V�H�ͼp�yE��aПR�	�(�x��2����c��ب��������;$��m��(�T��Z۸'+��L�ܗ�E�����B�nbOU��sŤ���30����RܹsʆΤ�$�gv���؏�����D6����p��iQ�89\��?��s����?���t�(Hͽ%�:Kv�CP4�HV���BAF<�	Cׯ���(��N���K�$�jc�W1� �/��n'���x��Rc�W.�& �FYt�K#� 8���:���E����~(DÞ!� z}If8�g��$�!g�>-�<т��� �����_8�u-D� �_�ZL�rY�c/@��#�bŃ��µ��+-�du"l�7D�����Eq�[��"��{��M����� )w�Wd8��Oq'Da�)�`�XF�}��f`�1jW�S�7�/%�����i���̂"��!R����.ls(ܖ^2����;RN�� �t�"�� �*Q�hf0��j,V�^bS�?E�+�����z%�X8Aq���N�U�o�!�ޙF]gj�qeN����z���Q0�����:�xLQ2f�'C%�E�ӑ�KmD�5�G<���yk5"�z���yC3���0D��R=��M[ ����-�,�*�Z�h&M~h�2�������`mj�	C �Ir����YX�|G��T�tĹ$��$o�݃J,v_�Dv��Di����"nF���YMs�k�����v�Lݻ�x|�dak�� tL�b���6G�G4	��B\c�j�pKrBƹn,�n��g�aǸ�7��j�48k`��s��z�bz��^����L�1>p`a7RS�n��Ϫ,��6D0�lw�-P1������1Q�Xu��qe�@�_�&1�+�|б����{�L�k�ChL� T��	�$D��B����į� ���2���rV��Q��U3R�{����w�3�I����<h��$���ÌԷ�q��
��l�5��ߟ���wY�����b���A�J�X�� H>�. �n1{IZ����V�5
��#��D�{)��Y� ֫	�XQ'��)�&a��/���.o���x� ���A���mD�杲�P��(3P�Ev�� �mз��s�t��שfdp
"[��l�}Tx�fP�4Q}唐�9�R�T�T3U�6C�����k���~*�OK�N^���Bd!�