��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��� ���/M��ٻ�x~�I�9������E">ر�Pۭ�^ztj�t_˞�x�,�;N$�k_Վ�N1�l��1O����CA�,U���2�8���ಟ���d��M.���p p@ɛ|����$�r�C	������)������|���\�h�@�>����Ѵ��Y�6�պ����o�9O��/u����S^���I�+��L�q�����9�w 	�"����t4O|�v
e	�b`��3(��������ځM~����[�Ą�#Vq�"�� D꛾|�rX$�!��<D�R`� 5��!��"��m�l&����|�Bp��u	�����N_�/���%��7����`j�d}?�PT5*����!����	�b9��XP����;�p�^�6ç"�{)آ��緵�o��M7�8l�;7ջ�֓�iߥ,��^n�ܪB��[2��	�v�!�����iOd�+��> ���f�?-F�8���茘�g��I�/c+�����,��m�`j�� �y 7o�o�GmW���0�U��V5ATwݘ�b8PA�',�D������`Q��Tǽ�U���!��V���s%l5E2���h�FHf�?X��Jy����y���=���朥��G�JG�ZC%�t��K������K�H���y�Đʮ@B����53���^<�=�Z�dU����쁫��u\<�T������P�q:zE+�E�ѷ/�'�E�}���K�.
��r(u�ׯ4�?*ta�zPk��K~_�qo��/�_��X�e��ɢ�%h�!�T��(,� ���^����$_04�s��s�Qj/~d"��S#�$��Ӓ�x�#i+C�q5�׮��x��~;���Oͬ����Y?��I�G9<��G�%M:�`,2��1�2X�	�n&u��0� ���(���"�N�R���&t�@Ϫ�6|݅Q��R"\U������,�\]��>^�F]"��Uf�q<�o�lg���2e����E�]��N$&���m���|���KV��ٱ��״��8?*�pPk�U}�<�3h-�i�xI� �B�Uj+���)oG�H�]]8���O�C"��[$}��G:	�Y�&Zʩ��6��y��=�K&�VDq����w�F��d@�ʓZ����+s�;Z����1#"?5��AT>_���]'��g�^@����ԆY������1�+����b�R������E�8PQ�4���R�Q�0��}9|����(j��jZ��͹�L-����ФK��D�!%Τ�p�M��+t����F19�
Կ�����m��Y��P���a�lI�%cc��!D�j�);��R��K{:%K��U��a��7��N�����hE#���`����e�5G:2^�52ѷ=��1`�w`P}q�����9����O ǜ���>�0/"7���U�A�4��I�kH�l������ˏ��N�;��/�$��v!��G�t���|܈�T.���5^ы"��㸬m�#�Uúk\�n���_�x�`�Ȥ��s1L��5�gV�w�&�K�W�������Bp#b�����|�g�^3�ߜ��u,�4yt�~�[&�4"0�.0.)T\��E������L5�	�N���c��Aـ6qo�^��r�nVG��&�2�Ӎӆ��B�D�$�ܸ�y�]JV�#������L}ڗ�y)W3�P�Uj��Ɩ̗)A��۷{�Z�d(e�I��\����$A��S��;]�hZ��7����Y�v9��**��]z���7�Ǯ�>��( c\z'�KX�LBjw����z"��{	�CPxGTp<쳣
��h�(��W�{"O�9����9�0���*	�m%�7���F�th���"~ㇲG�G+c��z͵ Њ�/�t�H�곒�/)iyYZ;����$�D�
�̪G�����!K=���}�#��J�?�����aΗz:8�ɐ�x��U 9��r�G�zy��_�q4c�����s-�ya&ʐ^�M&E<�vx1��F�sqft��0���4�6�:t���� y�~�ƭ��NӚ���c�n��?��E��K� ;рZ��V�k�P�*�J=au ��L�'0�[�f�^�=��-�V�Dm�^�Օ��$���:12j8�9A��B~^,��i@�Ƌ-��Oۭg4g.j�U���n�B�&()���xNV�PE�fM��G�$�0�̯�.{'V$"�(��!f�9R����Ng�/p>ҍO���&=NS�o>�-f�������O�"�'��^�����FgK������M�����q�֏6�n�o-���N�Aeh7���M����Th���������>mC��9I��K�CTie���LR+�O�Wھ��s���eS���T�}�t����XR���&&�g�a>��h�=nF&���oc���ؚ¼^.�Vk��!P8���ч�[�w��KK7�V3A�*%�R]V<���S�x�.
n6�x1|���P!�k衬Y��U'�Ψ�V`ñ��S*��-J�t��g_%�L8tv�>�A��a��0:3��m�0�Gw���/,�V|;�%��:�M	УdC�.}�2�������u)Qp�V�I�0$��P�a�x�Y�S��5���WJ)�K3��Q
��� PPL��O���y��?v�@d�6T�R����c4�x��A�Z	��w
�<'�M��D��O�&}�H)� UT
��T ��?\�w8·*� �'��r�9���OY�W��r��0<Ul�����ӋI�nq�����a��6�$2����6-k+�&���)ׁ�(t��;>�}�i�fIns��[Y��j6��6�S�ukR��2�Z��T��m��_ւ�|��!H^Ԇ�o���p7b��N�,ɬv���HU�����/�Xy/@f�*~����C���u�0l��v�m��GwNr�í���\	�:��l�ٿm�D����Q�m)2%;E��u���`s����~�������*Mz�Xɺc�I��g�|�io��7UȪ�_ON!�^0)���l��B�c�Xf�6�`M�Ǉ���>�X��[���r��Е��lh����!�����_��ty�Ւ����/9�B.)ڶ�}�h��+/��iN������I���[y�d�"/�,������ZR�M
mp:��{o�󩄢���)l+b���p�VaW�DV�mG
n����m`�\J��=%�&�e��d�T2���hMϞ 2�bz�����
��@q%����iv����n���yc�z$W~��bBb�c���R��R0����v�r5��:�h�&���U4��7��󰅲�l�V�U��M��Y�p��"���ǌ�Q.��FL����j���K��!#0�?����Ď˲
����\��a���pJ	���8ؙ1��&�2�9�<����wV�ڹ�\� `M��NӍ�W�:��4m��e��=����D�f��k�2�Yj��SSB{t-�<�<�mS��Z�2	%���z��F�����;&KU��9�'�b�'��Ȯ2c
�w�v��%�_�����ya��@�d�AX�yV��d����
Yあ{7�w1a�e�SI���kV2~wJh���ͽ�N���ީ����sr��l+���FR����w�|�|.+��i��Z.��x�eɰ�Pg�'�]C�bbN�G;9%� ���@@�Ћӟ;��v��z�ta�C'���)�j]:�K�P3�j\�-���b���jW	b�eJ�*H�r���pX@�v��m#B��� � #=��b�y ��Ў��+�BN�������c�K	fQ�|*�0�Y�j~Q��`���Y����l����N���b�	��GZOеz�IGv.ke�L��Z~��������ń������^�~<G��GgM��5M(�(��ͺ�_�4A�*k�j��2Cɘt��?_Kwvu��L���y0q'(�� c޾��<3CJF>�`��=���'ZN���Þ9�Kg��gï�`�R�-�ڏ�aK�)Wu���0��.(��Hd4-��v�J�\��WJ�JC����rh��$p"��}�5e�����QUV`�l�oJ 5�㵗�6a��SC��=O8z�UL�cD_0�*�#�w �SI���G�%sl�=f��&&��C��u}�~2����Ō��/���i���Y��Wt�(��}�x���������#��|�IU����x~C��(��.MY�Ǎ�"��z p"D�~3+V,�P�k��![Џ�謣���rN26l
 D�b�b�2���{��)m''�&��y��}����$Q�Fgi��l���	"͂X��o+<��w�y�t���2���g+��P�����(Y�p��b��T�^'�p��\{sp��X���_��3b���$Xz�.���	J�_�Kb�q���fh�l�ג�GpLh��Ay�M�D�@���I���ak����� L�c��x�[���v�Ê{
<p+6V��C,���z/��'�>�V��22����^*m��U�zhx@V������!�ԏTk-;'d���3]#(痬�+6ؿu�W����!�����&4�%�p���A����AH|M�m�.f^�U^�]Fjx��Z�Fg���K��s+�6}� �#M���4�$�a�������M��y����3Ew;��Vo�!�}Ga8��8�J�?����=��v�0�� �:�r�a��`��o�d������uTaJRcb�=W��4���%HuCA�#�jh�x[�� ��Z����G��:����;~�\�~>��91�ae���s�ly����(�s�O���-Y�k�� ��IG��5{?�n;�@�O� ^_f[��j�T��S�
����+XO�Y͒�\I���b����[Gȴ�1Q17�Z�'y"a`�������h��� ��k|(;K�H�i����YN����'=ֽ�&�/�W;��u��u�O'�v��
��x�zO0(��lچӳ����#E�>}'u�
�iu�����|� @)q�go֛���3����t*���JI{�Eg h*&����$�`ȝ�xE�]�E1yO'36�G����M��5�^B(��+�L��?����Ǉj�q�P��#^�zbT��ڭBK25��d����=��m~I�X��YL�vt��� ��c�?}�/�Ѿ�Q�6�ކ\����u���D~c�Q�e9���'����s�� 1Κ�v%��*�2`d�f�+�Y<�j+�{kA�!x���d$��*�;*sO�9�K�)ت� $�L�ƿ�;������6����	���8$���-n2��O8j�����z\kƈ`�֓2���7V��{t7���:�W�hO��D���pk<�rM�(�����_�߅>2pM�R�v&�A(�&�p[V�D�5{��V��4YNW�,��� ?��$\�>�֜���� ��F�����|~�Nx�
�P.%��dFh�B5��?)S6	R�  ��\,���.Q�� A��Ϲ���f��6�s<n( a%�;,�&H^C���#��">��%��˫���`{{���J�nE��i2��p����8"ؠ�yd��H�����GQ��}����}�M2�X�.���0��K�(,woAhL�Ak@,y`c��Eh��{'VI_�o�O�7cDP�^��d32�-e)�v���|�AZe�ǜjg��)k�gv{l��6nf*ToCVWW)���M�Et@�����T�lu����5�-c�L�Ŋ":�,�P�����q��5{���&v��l����6e�����$�zŁU(d:S�q��lc9���fTxx������-��'�vك�h��Q�ᵺ҉h=.#��F�L,xd�m73�S�󋬂��и�ej���&���̝���G�;�}!���$
vU�?��Jw*�U��'�<��̖�J"��R��a�ے����7b��"^&���@�An�"j-�y�7p�fs��YÅ�0)A���g��Y������0�j��֩#�L�u&;�?�[�6lK0ū�|��y6o�N����&;z�"]D/��se���=�w�Q�v�%�1��y�	��c�4MK���
G͟��U�ϟ. ��z�@��d��p-b}�|��]6���S|��_�g8ߥ��k6����2z����a��G��A!��R�g��j�\@��$��C �0�4'��bT��I��K�~a*�WYZf lp��H�V�r�"d�D�t}?x7�?��B��߷�itG=j�$��;'ܧ0����!��-0�0����!O������.��ی#�X|!��y�փ�?��c�2������Hh�.0�S[�6.�9&S��ľ��dj$���/�-���Ŗ|%���M���y�o,��u.
KD����Nd�F
y���ۺښ�:T� @�s��Ȥ���J���&b��WΫ�K�?��?cI�w�J�(hh��!{Olu{w��]�@�e�r��3�y�Cr.ta^ҫ��X��ߒJb�@A�0	b^����34�Z֪uf��nh޶׷�lWa�{@6@� ot��t��@�=	�������a���6G��� ����&e?��o������i 	&^a�Mƈ��b8����0S�����N�sɚ��{0<�����w
�c��Q���9��k�h �RԆ��a�0��q���C�;�֏�|l��u��VR�=���	�B�!� _�bl��J�nz��M��a����<�_J f�\�t��?[��>>oݻ_dHi�EV9�WMxBa�i�#�딴���ZΝ�����K���5���6X)�j_:���U�U"�J�j�jM���*�htFF���5/!�L����̀�n?�{��\���B���A)ñr(�N̙5"��6�<��kǿ�����?i�d�F���Y���g��ۦ�rI��#m�&ܚ9/�堟�ق(��V� p��oR�ѵ�EB4�]��w�蜾*�T>1TD]<�od3��f^����3��[���BGo�%6�+Gx)���47�z"�	��z�\`��hd�ֺqȿ j�
͂�tks6K�Q��ǅ�
p^5�_tJ��W��6Гk�z#ż+���u�#��I��)J�9[n<��d�{e��bJL'&���@���E�[.��#�)���R2����vm��^b>`}a��~
�pڣ�K�=��G>��������(�n����ul%5wӪ�4�B}��%�u���l��Zu���͏�P(7c�?�?�+�����o�M�������y1�{�D	!s����%�U����G�9�[����!�4�t����T����0��;8��.�C�Y�D��k�Yu��o�ϵ-��mh���Yf,��Į,�Cr�9�r|�v}�@�ō�Oq�huFuפ�:(p��v6�(�gԵ���q�2Y�����jFuA��9�|�ħ��������`J�zy4[�.8�5hd��
Gi�զsM�~�H���2s6P�;2�f��iA�����N��9R�O���֭B�J�����N�\�1�g��A�wpqD�
U)�B�a��~�@������P�'g�WX藁+���ɑ�s��aG�&��wM3�x��%�
�B/�Y ՞y]����u�.{Y�
Ls�k^�mֿ�tFh-�Z?��5I8�3�:y
�'>q㺨�bs�)��?�l辅	hi�\���
�n�[K	�]j�k��ɱ�&7w�}��L>���K�
�:��Y�@���2���(ٕ�oj��n�I*�u�%]�ժ]X9�Bp-�|�ة#�gOWy*����L���$v�W�^>�4�6rɧ1��6��0�)����5a��m�}v�?Z��<9g����YU_I����1��m @�?�����ሸI��l|v5#��̪D8�,����D�i<hi��Cio"�wpݜ$/���9���nP�E<bq����7�I
�`�!�M�©�jlܾ7�F"!u��C6%����<T=o����^R�S��^�f�Mi:Y�wa��m' �=�z�C�W�0��)�h �i��o�پ�_ԷPCE�P�i�Ւg<���'�'�m��� �N�x+�v�h�Q��m���|v��9[R��2c׌�Ȫ��9�+���q߯SLP�9^L/� ��e��٠��pxu{�+��~��%&���v �쳗�`�K�����Y4�mx�~���"p�Ap�^~�On��X^������lY�n�6����Q҃W������qM_���n�����-0�'�8νx��c� D�7�k�7a��FC<q�
�&�qN"k��#�_���v���W�9r?G��I�������>a*���A&��K�!��%k i�I�O>�R!�9*�S�N�9��`�¡�I�J��y*�n���K}�˫�7x 	G��"BTK�0P��ۑt3���r���!ǥ}��n�W`v���(�c�U�>�c0D���ܓq��TE�_cƓY?��V�=i2.��l�v�U$6�fM��]����A)DJ�N����J=�q�s��7I�N�QP��n��[m�����s�H^Y��0�SQ�L�>��~����w����[�A�������<�"��`��,����d#A�8��'�+c�kdO^ K�(	��ROӀ��f:�я�X��IĳD�L����5���0��@�A )�a�7�u<��G'�W?0�.iƞo�% o�ճj]��5�zX,��g&�ŲJەJC���{��0���.ܱ�����n!�*��R�#�<݆P����㖖!�|@����}�c���Uv?���`@�Ko�e7��X���(
����$3\�Ex�b��v�	��O���>quh�b��ǮC�������C�@�?�-|}�ĭ,�=��`"WQ��A
���}�,�U�M��ݯVĿ ��ϐ����I��'xK����)���Ym� ՟�k��q����j�(�]�n(T~���`5,��ݴ@���v0#���e�G.MT� y�àR��'��!�Io���e�D��o�`���D�s�,�1���1+ 6�D=΁�n�6��!^:X;&���_
�S��'�+żD�*�%��&�H%�]�}Ү���e����qq���7������� ��c�b,��풞���bDp��6�� ���b&������L�߿�ݎ�h�c\�x����P�k��S@A&��4�6�����x��v�ef�eb�ΝGK]�"�A<*9���6��C�,��_N\�M��%|���>ͩ綊��"�޸�)D?�f��@�~д%J���=��>���^9����IK��1��Hґ�7�B��|�ش���,��	�0.G-[�]�lҝz��	k���`��������(��ዧl=6�-`O�)qs~�_��	z�FU�
}��=��<�p��� �u_+n�Vf�,���6��9;���Ec��>}ް�h���`��$��Ks���Y��{��挡 �548H�jB�"#�|�������+|w�l��j|�*=���H�U~����}�
o��Y�#�&�4�p�cxF㸜\D5��s�w��K����{B�S�O;�A�@���տ�&h�>���E)8WS�==�en��RV�Ҫ�KcLw���7s?�/A{��S�o�D�`� 6G�Et x"�w���
g�,��>�`�r�~Y�ʲ�o�?�z*���%(�,�q���˗�a�(�u�����]k��}���ys+���q`����	��F$� �����ff�o�B��߄Њ�|j}9�����0H����M���=X:�2��YP9
�� D:��s�;����9��~�����z�<��~Eg����\��+GA�����ҝ')�Oğ�1q�(��J��&��N����r%�nR5�P*��A�%�}�8s�,��78��0Ы]�]�PN$���@�鉢�9�#2 1"Ȭ�^#��d��&��T9ް]4~�}HSjm$�;��*xmv��>���B�_���b�ث���`�3���Uc�/|���ITդ���wPo#2��DBh�Z�.�8_u��i���#�誌[9�cq��l���w�U�C��i������c�k�+��q���Q��;�]H5$��d��������X�ч�jU^qF&g}�m����3�آ`���G1w���='[���*o���d?��$��U6�,`UUAU
�FP�������!�ɹ��ȼl�Þ��%5H���]��Py�;�=(��
��Y�����Q+CA` y�2���5�[�ŉѳ$q@��5�n,+�\h�u�CNI�/t��YfoQ�i4Z'�ˎ{����σz5��t�����L:�Wط}ݕ�W�^8��Ŋ{�V��Պ�IÈ�kiѢ�I�pE�:�a� �֭��ـ���÷֩�M"�`�����4%�M�hѿ��P���%F˷�s��*>�	(�'j��<p7g>^�ne`�b�R�R��B�1�^:~<p���M���Cp�'��X��'	��G��}�@���k3uw.O�V[ƺD'��$T�\p�:�K��P ,N���P�U��Z˷11��K�m]!
ʼ[�5�w�拪Xc�����?XV.��!�9*xk��Q����^���Z�5�u�#��U�����D�^��خ0h��.��8F�\�`ݼ u>I�}��i�_ٶ�1 l���������j�@�%������/��:V���J�D�sK����9�$���� �B����8LaǳG�la]�K��z��E��g��.��w#��CTN��W[X��̤J>cQ�+�?߇��z.s['Q�IM�7���ba�X�� ��[ߝ�KbH[�w���dM6,��ќ��$	�Y�F^�$Џ�A�^���I��@����;�J��5����x�oޘP*������;@Z�t�JN| �\���O����M��Y�b�dv�CE� </�F	+�(	k�m�d[��T��7�A�q��Q��L77��σ Dx��t�࿉=�@��r�~