��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�7�Kۺ~�۪��������	�SL��e=o&3������]v<�1�,9�]�u�sH��<��K� �(05ۥ=[3�Ul���M�%�w�W'�'y��/�(��6�2u�����I٢1<��jqt��%��E�a��ҁ=�����u���3M�{c��co Hw��=V�|w[��e[����L#�yz�ߒ�el���t�̨�Q3��9�l�4�b�<�p��MnG)���T��Н���ٵHEBL1�ޠn����\��,��A��
����ZX~�C������A9C0@�"1ٿ��%2����N��)�£O�ք/D��
��rx�<�v;� �w�aO�Fc*���q��YX��s���ർ�2h�X
�]�� ��݈����Pw+�A������q��Rl9�*�e;�=��6s �'օ��Ho8���.;�83�4Ȳ�
g���Z߽&J}��;ެ� �_Ne5�Z���e�Zɼ>�|T���u��#P�a;�$/�Q!�CI�m������7�(�jz%EN��&����w��zik �v�_\�I_���TJM���1��ZP�1�$QT��Ey�R0��2k����29��?��^3$V�\��Wt�e�cTx��Aj�Sb�f)�X��/*����d]��-��JI�2N�E�W�.��P
4���.��X����cj,;G +�a�������S��8C�� U{$�N����PY�����%�,�i�ʱ��V�o��g+�)�R	����!��Yg�~���X�)$��1I2���{����zV��!r�ʹ*��;3�N��T�U���Q��P�x_���F�p�
C���F�������Vc%J��؁�X<-j�����DW_Y?����m�6
�f"\՗�ʅ��`r��O��yt�9�Ϯe��Q��s�_������Q$ϙ�Q�S�I�@��=6-��CT���I*���I���PR�Ұh�w�F<�8�u6��t]_�< �F�߽^ �D���|�}�߀�e��%l�H:��5�)�5<��c�%:Ac�ެ� ͧ�F���rQ����y� l���v�u����c������! �'9��~�B^mӇ�=����ʀB��Y�
�>�њ_uIv���=�v�b�,��`ߺ琮P��8�����Z4eKvip�{m=�ⲧM��&�N�Too�x9IP���#�}<��Q�s�&���������hЫ}��ՉE�1�D�m�u�#	>B$�����u����~���^ˍ�G}$Ϝ����y�V��z{��&��M����m��BH�XO�M@������؀����G\@!�E���G�aL�&0IY2]&1e��R��&�*�8k��3Jΐ� ]~�y��,��{�7�d�Q>�Ԟ!�'�M�$��yˋ�ɔ���E?*W�~(�h�V�@s����VDJ�� �c ���tY�w~(�o�{(�����|���^H�5���NҾ|$�\k�e�5�ddz�f������+Q;�]umw�v��>8����n�"�,�����ԎYї4w��U\�����Z��E F���`_,�B'J�T��C-+�X}��*���%��2�������\� _�RgkY��[�2tϟ#�;w�����}����� ���n������neٲ��,�`6�^oWf�ąS�8�x�dؚ�S�~�Vs�q�gA�WN[碊BwN!�,�!8]�/j:,��p�^([����wV+�@������,�b�\@��>3_�$|�2�fD�9�9'�.8B8�>�J:��x?�?j�������8G�C��g�s��C*w���)%�9���k�'y4ܐ<�8�5������~d&��/���I3�S_�E�@Q�x���e��X��fy�l�O[��Mu���:��������=KT`���2[1$��D�Y�RG명��j�TnX�鰁��+̗D��l�Hk�ݝ�]T��o?�'/c�&H�f��3Ζ����#L[�I&�P�qT�ꐾ�!��n'�>	C�K$pV�+zQ��Ѣ��c���%D�t4�N�wKV�B��e�=��{���|�"A-IAB��N84�F��1���L�(7Ks�T��I�!�+���+���Z�`C��l���/���>r����dg����-|�r��8�f���ǑF���6��2���ҏ:���X�8'����X�9��r~�����2��Y`�X�h���?욲o�)��T~g�,8 ���瓅/�OԞz3�{٦n���ھ.i?�<˳��H�;�k���ѧ]T�����c1�����6��Z@��㣞�?Ӽ���=Tp��N�=n���ex��B=M���<���>R���u��Ȟ��su��{z%6�z_�j�^Lx�qq>p���dX7��c�^:��@���#��AпՕo�BB-�s �F�a�Gd P�#rB���TWg�m �#�Ga�xw9k+>y�eK��(���vj�5�7}��H��ժӃ�Sx��^����W\v�(�7�.�`�6�A�MG{p#����{��F��F�!"e2��県�|[kA *�����a�1���jf�[�>/Y��������ֆg�e�M���#�.��o�2D朡*��#ʡn�ZOp�ME>FS��N�(,.��v���6o������ +ȥ���3ǁ���Y%�U����x� �3_�T,�����x�>��9ܲD�G	R�4ե�$�
Ы7�9N\6l���fګ�e-��}���HB�h�
��wx��al�$NP�68����uɐ ����� ɴ�%��Iq�6��Ǜ���kӫ3�\����+HY(L��j< ,�N/��{_�7��9��O<�|��Ve=O����Ö�x��@|o��B!���,���/�mN<�[�^wJ8t�� �}�NE�Q,;��rg�t�>D"�k;!�=Ǖ��VW������i�L�80{·�K?3�82���?36��Y^4�iX*+��.�-�l�Ьw���a��c~�S�*a�#��e��x�n��sg,����.�_['[��[$R��/���<	�[B��Ӣܻ�&[�z�A�tƅ��rO�@	m��!��iW��9��4Ƿ�o�pw7ġ�k<������D���U�D�IǎΘX[ţGំ�cY6��W�R�v���p�K���}+�����U��d�mz�u�_D����f�oճ�5�����*�����.!l ��n翌����aklHs`�*
�c�ɏcɘ�����NQ� �±�k.7���0�(R�[�c��l~J@�꿻ź(UR��%�1c@����to�L�#��&������}CWڋ:����v��1�q���Ig��J�vI\���0V�oT���:���sJCD���'�;Y���(2��!q�HI�e�ó�J�^V�	�:��G��l�E�"�0e����b&���U�"���2����7� ��op�Ӓ=9"MՌ��*
�^^P��b�YF�Ǜ�;&��ٞ};��ў�%V�"%�K�("�Ƶ<8�:�`E���t��L�E�3��q6/���
x�����܌�i�:�IAk<��8�_���h :zi7��	%�� ��!�nf��:U��N�6���� �X.C�2�m�dI2��mWG��n�D���|{�P9�)W� �u(��\�hc T��P�>9�Ʒ��5ܐ]�9�?��\͒�|�(
#5g'̹�s���B |1L�
��룒K�km�߯F��� Ž��.�:e+�fk��Ff��cm�[��5��R�e���31�})�k�������^,-�.�WlW���@ӟ)�܆7C`��
���"P<B�A�/aK�Y,�bs,�8��Y�������><q��1S�O�J���m:$ܤ<��U��0c�[��)����h�P颱.Z�M�K�1E�\yt[aF)ce��+�L2L��_t�3I�>^�b���۲�J }"Ğ�$��B��M�%�Cރ��d%ot�<JA��%𮮵 �}���iD�LY�b|�;��Z��+�F7d��d�ԺE�N�����'G����L�h 
.��_-<7wr롫���:��ld�W!��U���"Vp���g-��~�s�W�y<���ur���p)�3uK�#�M�KW{$���N�����U���#�tW�냒iilvɈ��iv������3"�����UKC��Q��fZd���E]٭÷n���8`�#��b�^⳨�⋆3?'i��l����V�[8���붺�wd�s����Z.�0ʠ�؄^E��ܿc�d����=K�y d=P�?:f��>�zb�iG���(X(o�	��&�2a��-��=��<)u�*[L�L���9�n�M&����'8o����3}Z�W<d_^ 6��)�-{�FVvz,��h���<o;�ߑ��ꙧ��O)W�:�O2�*;oYA�u��e�~�q�Ə��aYao}�'�R4w�J������K?��l�:�]U(P��W`2���1�@�KG�j���67��q|�y)AE�[��uW��"k�BŘ�~����/ )�y� ��Q��ཷJ���ɱ�[� ��z�6�4y��[N֧K�*ff��ɒ�HC2�$}�~=�	OȈ�sQ�ss�D]�u4���"u a�y�fL���O~�G$f�ȯUi��&��t|@�C���U��rJJ��u�Qaޕz0��dE�_Y�{[f�s�&h!^l����q�ue��Ncĝ��hI&IOK����^u�8��M�h��v��k��jcJCyN��bp8}J;��(�R�2po*(e�)�B�Ґ���V>nk���6�ۋP>j���QQ���)nw{/��P��[m��c�C��~��0>E��)����i�|U�{c�Nۃ9(Cy�a�nr*��ųx�ԁ	��V>��;�G�0���Z� D������` �X w]�7��T8��&��_A����o��0h0*]�{Z;�K��V��2[TJv2���&�1�g���)ȋ^W�+�r����F�	{w�d���?+�풄��C5��=���,{��;6����bݑ��f���{�|.�Qʅ�B����Su���F����]!u�˘���͒&�Lx�0[?����S��y�;��ۃ������GP�za����D`�Yޯ�f��M� 3e��6�]��hE���-0����a(�l��h���E������"��ސ��/Q�Jb��#r��U��)
V��׺guW�*�����9���{��&g|��ҳ�Oɜ�pNZ��/$��+��߈d����,�0�����]ݲ�S�O(�Rt�'�`��L���m�f�j��ɟ�exP�[��P���EލD��c�J߰��ߝw!�!T�n�(f�^�P"������?)��������"��T��Wj������������+i{��	O�y�_�8af�1�L��\J�`��Y�8�1�b�xF�(-�84�?��%�̳x0���L���D@Ӡ��)kW-����N���Q( U���N	�;&�h�QU��$�B��;l )�$H��h�s+�����zm ��.�����a�ׇ7_����y`\B��
IV�'ا3/M�H���x��֊���?�<���i�=�TK߿����c�de�n�7������tm�瑖"�����M�>�L��Gݷ��h���w�'J{Eu����O!�P/�C��򤗆�x����%
���V�'S`{��S���K!�HOI��a7���ഁ
V��E�����n�Ej���F��"�&%�~{�R�!�Ԁ@���$��(E�h���6�I�����Y���/���0^R�{���뿏�e��\x�6 ��l��ktA`bi�����HB�K{j��˾��Z��C����/�T;�e�ʪ�d,5+\4�LL� �U_�*�jbA�0-.�k|Qy�	���]�Ė�A�a�*������8=	O� �Q�ιq��{VȾ|*��zJsK0�P�*۵�O R^���ڔ����0��b�!�4�/K����zA"���.n�hb��8f4�����u��p�Uy*
\���ٷ�H���A�����0ք��f
_��%����Ճ�a}��[V������Ki�;����@��p$��� ȩ�m�$%Q>d~i�R�P/���ԙ�~��F������W���e���V�8o�_�2{c�]��9�PV��[�����R �b/�9�J�9QL%�$����T�i��ʹ/s����]���)��ԮSn�r�Q;{��ɛ9_��M��������p��'ބ��o�[�\%�N&�����L�s�����i��@�,�u�vITC��~.�?��%���y@�y^6����i�����L�ej'��@\�J��vO�,n_�g�>H����=*��Ǽ���tvf�S�QVL��{|�8)����D{�D׾�����X/ye��Z�&��ʕ�����:�0��㮒�c/��BE�����=��!7,ڀ�y`�M����^���}PR�.ʙz�D%���pnja�O�	�p�d0��2/E���EQc��H�z����r�c��$2���_�JHȚvYH7m*U�Е�8�_�ՙ�x����e"�ѩ��ր�l�0�P�J}���)F=u��.�y�6$2}���U����A]�.�Tu|��k��|�ۭ�������4; P'K�y�=Ξ�,����e�0Ъb���
A
^�~"��������=��
�r|���.���:�-��,<�k!��dұ
�E25��f�}�X�(��,A1M����\V�8��Zl�T+�RcyOV�����m�1n��h�`b�G�^�g�(�`�ܙ�T��U��IY���C'��-7$��-T�M�2s0W.�FZq�I:P������5�:#D��
��ۋz�gJC]��8�6�9 6��ʧ;o"w1�  ��4
@����Ө��MQ��i;S �|�/����M�N8/\��I5)��Z�(vѝ:l6Hf������K�&c��g�5t����ŧX��7X�	nT:l�c<�k�R��(A5�۝r��5�����`(=�O�����.Lp)���fG�ݹT�넍[%L���z�g���$���G^���5��3�nc�f���	�*^��ੱ4o�����X��(
^��=[���Gb> R�9��8�O����o@{�/H�φB���<��O~o���'���j5���kX��5���ֈ_��F�|�����籙
��E��i�x�$[���?�A��j�t�o���q�|���.��a1�:<wc��EP'5lQ��h��	;i���y�e�$jH��u�t�2ğqGN���Gh�8��9�%���M6������u���m��8��eMDx��K0�`���l@�ͷ�;f]����,Ҟ�\+�{!5_�JU������&��<����y�$�ΰ�iԓ���e0���[ )Hx����;J@�	ƾYXT��8�]븹{/�t����_������zm�,r����L��p��lb�џ�Ծ�3�k����S��*T?Sz>W/r��1ݩ�KV)I�e�.�+|γ���i��ؐW
\.�+���q�"z�/��o�E�Җ�>��^�<����%� �=�MWJk�a�����<��p!�� 7�V�Yʐ�E�_�r�"��eGn��\������.��(iu��Gmϻh�i*+
�L,xی��M�RR _/H��)�	+�����������y��^l�����4H�|�I���J9R�t`I�L���5�-)��"����{���TB@`Ϳ�����ueJ�[�S%�%2�����8b1�Q��w\W�֐���ʿ$J��ժ��4b�]����%c�)��"+���!�e�^��KE�J������_'�l��L}Y�����7��Ӱ�=u\�ޥ�[q��E{�K)��/¾'�˫|~�a��~�,�1�b�7J1�=&��B�Z�
�YDic��^G؍���A��QJ4�M���&,�
H��`f��3���\f|t�v�/�E�؈ds��ђU�&��:D_꤫�9�`���0�ki�L��.bQ��Voݗv�GTb����傘&'5��w�Sq���R��Ȓ��2����R�!��Hx�����a�ׇTG&"'�O>##����Z�m���~^{ZD�����h�LHRr>A��Ȗ����#;����	�Sv56X�
 ���@
����x�;��mN�����h�K�p* e]	���.Mi"8��OW��:�b'����� ܝ�����F� �R3���Hx�1�ǋ��>�i�hb���D�j����]]܍r���u�Wo~�95�%$�]r���p�bv�v~ZN@5.�N��ͮ�6�.��_9����UT���x�5c�ծ�܉Z悠� �z(�w�{c�ǯ2x,M,�KV���%�{$w�XE�7*;Y��^���a�,�ȗM����;^���ԗc�˺hE���f��F�C�?�w3�͜U����i��~}Dh�gTA�����:�ᲩS�Uo繩�~�?,�g��/)�wާO�'L�Tƹɝ�����V2L�[ٞ�������Xb�/���0%�����Q�a��.�򥢮M���#K���y���w�5J��V͞B�C<v̄<�\��9�D��v2����^��򠱂r7��!u�(�X�XLگ�x
�
�(�@�����-�a������h&��ٻ�͸�����{���l�@�0b�������#��`̛�Ozb����ʇ%���0yڡ�j�-N�>�&u���w2��b��Zwz�_��ˍ,C�hŅ��\e%X#�D���7��[��)ķ����'�J��(�H+�f'��R����˻k�7�|݇�O�:WwA\�0�0�O��{�C�r5v�������z2s1)��ތV3�+�O�~����~�e��Џ��4�	�J�xĈ�.��%<��v�9��K�=fЯ�٫î:�'�x��k]�油M	/�9�k�ˎ)��9��{�|$Y�%�)7+�!N�C}4yZ�ZlƯ�m��0.�RCt�la=�0J�ݨ�['�{	����T���5�ө�k��S�J�s� �x���jdz��]�	E��]<��H�Û��t1}P�r�:@��/ӕ��?����]-T$7)���:�dNz�&c	�qf�:ev9*���:�>wե�\����,1�o�l�g�,a�?�axz����B�lH1qu�y��D��H��Fn�s���ܺ�g��a��dy3v�� z��l׫�=��*I1���~h��b~�b�v��#��l���6�K������U���¶39B�����v��/|S��h�)y�ڠ��qZ��M����!�Z.���%���)��|����$@iB���q3v���\���$dR�i�Q�i�|���I
�w�~!dG���Dt�𠩵͌�`���
�@�.�S2�a��D�������S�����|_U�v���6=�)/�t܌t��������jZ5l����3���u
 1o�9�_�cI��Y�S�4����X��'�^1�8����&&q� xC��CprE��PovQ@�ȝ�Ǆ?��9�<����L�,<�<������VH+��m*��������I�%-Y�c�5d�8T�^�̟f!6��i���peQ���/W�ǧf���``d��]�#6�K֡�hk|r(k�?}*	�rEe���r�~��!Q�����Yp�h�IE��!����K�^�x� [�{�\�u��b{�z�6$�����ӡ>��_y�IP��.V�3,���T�'V����́�ۊ�L?����2���6��h_�a�C6�dOɍ9Т��dv���n��Ac/ٟ6u>?�[L�����mw�fb�C�.��((]#n�*j�6&�,C~�O�P6�ގy��%�M��vJ&F<g`������1�g/�f�}�=ԯ��~�9�*�^���ޓ��Җ��X^�ɱh-�bZF�ݮ���k|���PX�����nqEi��`�dP�ψp�p����/U�$���wЍ`�@�3b>�k��P�\���ݕ�����0�|h�W�J��+����gP�?����w0Q�ȼ����d��=�}����X\�K�w�pi��"�"�����dJ�)�;)�j��}���"�+���s����>�q�����V��R	 bܥ��酼,r�J�.��ya�s�~*��+�3�h�8i�n�&z4�Pb2��襮$��ڃ�j�س7Se�:�/B�k�ړ��'�q���&.�ߢ[�R묫�+�o��>-�>�8�a��
�0[�ڹ�OA7�z|�y�I���L����Q��S��J��*��!�}��T�#�,o�0���}��{�K��o;M@����5ԷOQ��'�����l��0%Ȉ�I�����1$�C*I����ؔ�r����	w��R���6;��9�⢲��{bs�]�������M���+ҥ��aP�䋚ĸ��Z�_�#Q��@z\;*���2�7��3�G�K�ߟBK��˷y�-vK����"�޼����ZD ��ð�i�n,Ǜ����M���2�B� ���'��v5�}eW�B�羹պ�)�$�)"�uJT��2��e���j�`9�Am~�$����A��ɻ|�������w"�;u��6�'��d���3ܖg(+�xRۺ���u�q���-�R.(Oԑ?�����፜���<�m��>>V=٣Lh󼡷˺�*������\�GEz��ˀ;�(%؀��z��\YLH�
I6)ZR�r��e���L� �̈��M�9R����E�u+%b��9�|�/�ZgE�"f �I��Y��e)���� ������|fD`@�&�~�.6 LO16�v���nX%+��0�8��H��NGf�p�j@���`�i��~���s����W��#0�ǙDDs�-��ZC��D|1����]id1���}p�9�W
���w��ԱU� 4z��]9��v(�?&_��!Q��O��Ͱ���K���h�
}�K�i+�ZJ#�=�B��Z����$�UC[�����P������%��o5��y��r��IO��e�7b�:wv��5d��j
��t"i��f���B�xC�5�tU�~��﹜�<yl�f�Dս�q��6f�{ؙ���ȴuJ�g8�_eo���޹��%��gʚ08�l�FsO�����q0*<�Z�����3��Z�ϐ�ƈ
�Fn�|W.v6���7�Ha~N�a.������gх���풆i��nI��2�T�6��!U	��S?�*��̅99/w8~A�QY�����u�:�=dSV�9�#/>`QX�����bE�1\D��90��U���Is�k,�T���0�n΅�B;?#^j�Yv��-�T��ȡ�c�zv��߳<��i'�d`�'�U��~
5nd�$����)h���p��(��T�����q���s��V��91����?�`C�~؃Yt�����eE���1x��h��=S���0Zc5�ج���I���8���g8�:fAh�>�m�ᗔSM.% |��R���'��vėay�������<spF�M�w~��D�Hǥ����#y^�o��hP`?_z�3��	щYKn�f�ȴ?Tɉ�K�*���j! �ّ�Dq;�s^
�IAqƃV�k��ˁ�}�!D�UQ:>$�]�gՔ3�'�ã��F\��,����?���}�C�+�}�d�4�B#|��V~uW�s��g�\e,�N���L1�O��9���f1 ��֯v�;�H6Qs�g�=�k&6b�z�	?uFҤ3.���ʃ�j?�L�_��HO�<؋����(U?�c�,a�_&��YqB�.�ROKp�)D���~��N�Օ��[���Z�Y�[��0����}ΐuoX�	����@9����5�k�k�*� '�V������Ě�b�$����$`v~_
�^�R���}�&�`U�@\����w�[�ٟ1�.���x�Ds���H�e�	�q�d54���Jj����1^���6�d+��Mÿ�����3!��C�����d(�r���N�PN�=��B>rGV��+T�{�>��Ýi�$�6�g���R�ݓ����T�Oc�Sh5�w��E����S���Mh
���2^V���Ğ�b��q��D�]~�e�P{�-��c�}e�G�I���e!ߧ�P� ���Z{��^#�o��f/�:N���m�Y�%F ����4��=��[��G��Ǽ�x��[����t��l��,��u�%
9�{���-0 �'#L�)�ڪ䞍O�l��fH�@]���O1C�(s�l����vg�q߮�$�o��;���UZ1"e=[t��>\A}$������=eqe�r���/~{3��[�u��p����p�����-�U@.�x2�	�5ĀuEߗ 75��`����=�		J�G�����+3�x���E� �k>�Ga �����v���[~o�}>jJ�'q������0h��{}�niբ[є
��JPz$~+K��Re߱���:�3��LҠ9�+o��y����ڱ����5pp�QJ�+���Jc��1�L6J�o�� �������	�s�H/�"Ζs��QF�n�������$�xUn�I+2�8��v�����{* E��j+m