��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���ڿ����à!����; H.,�j�gN6�<���( �78"�����MO+P��e3�X��_�qz���R��/�MU�z�O7��q�
�J�<���eK}�_>Y*,fӃ�!m��S32R�V�6g�R��Io�6R�nVF����]"���ț�L�݄K��0xe��f|��!�I�m��-�����s=�|���F S+*���W�a�b�;��?]�,~[ʡ����dy��)*\��O��t�2�0�q��i��ã\U�:��E����ޙ��hM/�hsC)�һ�H�7}��Ec����|��WrR�9q|�рf�8uƊ [Q�?]֕�=���<�#!������.�D)�)�r6��UM�4Wm4�(�B>����̯�֝QQ�ᛶ//K���Ff�#�_]w F��MI���_�X��D�
����w����x\�� �V�h�=�:LJ�I\�iKũ��x�5�p��n>3�T�)��n9	���a����E������~���;�}���#��ԛ4�q�4�Г�1BB��KgJ�.Lޢ\f�@��2+C�`	�Ñ���s!�0�Li����`<�r���L�P�Ć��J�QmaUS6�t78�N�%)+�3�|�������;��d$Ni-lɴ��B��_�<�D,��t�F�B�byM��c�ֆ�#��CU��A�7ꬲ06 x㛮��0�>j��Qթ�t@�Q�t�w�ܚ���/@����qߢ?(Lp�z�Z�R_-�M.�i��{e�J���ձݺ'���i�w��Z�z��͢��ߒ,�n��&~VL��>bst�7���c���L�\|�5m��ȄUT�0���=�o���\�)֤ر8�/v;����*w���'�
�{��>Ƈ��"�YL�Zv���g�pY��o��\����N������F� 0�ڄPj�8Q'��V�(���lZ
������ϯ[�,Ut�������I�u�\�	��~܋4��{(���6�V�3ַ>���@�q�օ.r�xq��j�W�;S���:G��O~�BIn�H�?1��� 6 /�X��̀e��y:��ַ4ed�X|��״����$-u�@�'ohJ�V%���e���fN��~�d�0�М��Q��-"2:�T�c�cP�ª�0Tz�8���"�KX�k5r��J�2L���3$MbBK���	+1�c伉�氝ے�m��/�}��mwf\1�'�Ȁy4��>���k4�L���	'<��;GW!�:�
,)�s�dI�LU+�=�XiCl��p��PNEXZ�Tt*_97��Ղ!?�]�N.�>��ݜ"-9j�Hx�t��(P��]��Z��mc��<��y�
dTYɲ@�'��O9��_� =�g�B�Ȇ��Ya�d���#&>��F3*���d���R`7�ՠ������>������Lv��Ĵ4@߮yW�(��N�X�ޭ�7D�-�Iv��i,�Mͱ ���hh���)��64'�Ί��Xg^�����E��v�h11+���zd������ȯ�D�y��d�2�ҕ�V1\%%2��}���F��)����*i{��ԉ�g5Gf��Iv����k��%�f_��h���gjh�ε<��K�]}e,�y[�)(SWK�=���*��s�� ���~��蛙ꥵ5�-��Pc�	�_�Ҩ�W}�]G��u��٬1�_��f��#:�"b^G��	��A�WxU1�˚�'A?;�hSW�~�T�mVx�I��y}�2Dqt��C�:ػC��� ���QS�����1\��O���f�[v��U�o�큂�)��������˵n�iB+/2�$1������1����K�� A����~M�y�fdO�>A,��B��7�
����W0N�����"iL%�B`���4�d���T/A�]��c��y�����еBT~Tp�	S^t=qk5^���E4�-�;Biu����Ԇ�NP���O,��8}E6�4[@�ϪOQ�l���	HU6s��:?�^\%�%�"2����\��	��D��$N2*��A.�B�X;���荢�8�G��$>'�d����6�B$�#�{�Q���>�K6b���1���^	�����֪>�l ; �t�d��mF����?N�x\�$lQ��(�W�?hD�Ԝ��z��w�%z�ebЬ�]DT;TN>���H�c�*�;>�MZ�fv�:�&'ʸU����h>��H.Z�]���G�E2Y͈!|�"{�z�{ Ḙj9�ۓ�s��zȍ4����Z\V���R�]���3�s9���	W�y�p������T��K�\]��fH����jǈ4Z���z���2Ir��b۟�����Z�
��Ա�@6V2���ĜƧ�����\G�"G�������OUVB���"�Zo��*�c�� u�17��w�lD̎�+�t��C5�a��0�� z4Ȃ:�%����H���&�>�3���.Ī��!�k�0��pz6��l� ��L�30������$(���d�0�$�$r�N	�4����X� c�ۻ�ȺU�����!��UG��x��m�뽼,�	���n�t0�7�&�b�8�~[����߾V�HD��q�p���F*��*��ʒ=�FL*w���s�;Jj���?�,�6�]�	��z%��՟n�0=�M�,���.����;�#����OZb���r*�=j�N�d�� ,����-����N����%�}U.Z{w ��$�r��L�.yF�'��|T�p���ОW�W߮�`�8�&�>^G�!+�i����efȆ}:���fk-�Dl�9G��(�����"芨>«��s�D��Ks���e�������N���C���ڸ�j�>m"�H7��K�q*��t&���-�%�[q`�����P�Z|��#���kǥ��AΘ����ޞ�F5&%g����!��;�� z�Sa�f�M�� u�2�k��ӂ�73`�v�aW�n,@�D��*�F�S$O����+[r����{�����6���it�V�?E� RM��juCH)�r� �NI�6vIm6,*��N�,h�ui8;�S��2�@?�S�~ߙx%`
D�����n��N,�챴�EO�k�%a�j����p6$�B�Y-Y�t����n�4;}Px4�Jp�7�=l�wq���3⣾�)�����qT�{[2����~6��X[$0��d�t�6E��ϡ~1if9���	w̌��S��G��m4QC��W3�
�i��n|����n���b�&5�c?�0��b8ԯBO6m��R��r��c�X�	/b�m�Ym�R���~��a��]�[��J��*��R�=�㹿P�b���xcX�SI[(IҚK��c�N�b���2�vA��:g����ڥ��
2���`Dw��Te�*�.�pvl�I�fu6A9�f��]I,~7Ơ���JqF��n�tu�����S�g��#3{/�2�k��aHfd��n����]���%ك��怾Ԉ�V/�̝�^1�����C��!z�6��Ei�=��׺���(\ �O[2*�r�C*��^�j5�U*>җ���T�q�=�Pq��_� ����3�K7_�~ ��+�k��#��t�V d8�Je�B���>���W�3/�Z�$�s��к6���21�ɚV%:<M�`=@��m���2�'/XgT�����%���ĭ�J5A�Eed�	��.�+��O�rT����������®?7��N��q�ݐ��������\{����v��s���z�ﺗ�J�ƨ��3��92o�PV<i�+��]٨�4__��1s\\�Y%�D��/��./ì�H�q��.��H��|lI�%�dR�q#I��	��nN�$��6�VZ�9;o�%�O����B�t�H3'1��!��6l�|0>�{e`����a�9z������b\2 �تT�y.el<�ە��*����3��"�EH�]Z��`�= �qm�@�/���Ә� 7;�G'��U`�{(m�Wѧ�s��y��Y
/d�z��1X�0/x &a�FNz�w5��7ᯁu�kw������Ȟ��)f!��I��op�e��K9�;F����I��W=�����)t�D��g�ṘPB�͋�f�!�$����>�B�����89p���P"$�ע�VE�^o��n�Q�mih�4�!��nf��B�t��BlH\����I�S,�{�������i`�!d�����5�c�O�.��B	�t:��b6k�R3w{����sU� Y%t8��
"Lc�C'���Z߱G��r &$��(��\���M�B|��{ie�i#�@�|~�>�6�F�IShV�i����c,�w�z"�R��ܪ�"�##JL*��f��_蚏����ߟ!�tt�I"�O�L4�9(C`e\��fq)*����?j#���Գ$�^B%�y!{c�#I^}~7-	^���r�Z���d5/��$o,L�Ay���Dď���[�����f���P7[�.������-�z������_ñ�U���F�wN�(>�}�φr����]\��ǁ��AI�+��@��I���=3�o+q+��&X0�Ԙ�=�����3
Ө�
.+UqT�4���S��8���GQ�L�cK}���2�=�����Թ�v�	���ZȯݞЙ�j�@{i��`;��̅����(��m8#��&���8g��0�9B$�]P>Z�ޑ#�d�)�����~Gjg�<�۷����qR#��S��4I��p��G��3�nn���e�Ze
���R)jF�����zgI��0y�
�[@�V��P���|��iVMĬ��8H�b
�ga�i{b���fin��Xd2+�i�����w/��fӁ�c߈���Ao*�,�,yʂ�����+(9Ƒ^cޝJ���^�[{��6,��c&�?�x;,P�^36j�p�dk}5lؗ�(5�����4���Z�lg\��H-7,��'�,��jr�A��B�O�]ە,�F�t��sE~���h2
���֟��k��D��-x t#t��(XF�kw�R�=�^��!��Ʒ�.�2
+p
�՞�����?����֜������·}u�K���-z�8]@զ�M��'ۿ�K@y;�:�R��GsC~$Ʃ�������׶]�̓9B���5��>�,v"M�SS,Sr>�D֛] .[���0P|�V�-`�[��jIq�ނ7�8t��Vx�v���9��#qE�b9`k�//�za}�!��<���j���5��͠g���x�}l�Ob���x�nuT�hI���%���i�*��$��G���	"3"%�����8Z���:��َimfx,������:vT_�S�E��nw~D��F�{�Zf�vK�3��	t,��x��W{BY�b��S��'�xc���s����[;:� +z��
�6�O�St�6��pܛ��v�)=Qv���R�����W�	R�k����8y�d�!?��ưᨄf�<kY�D�~s\��?*gV���)b��m��C�zd��B(U���9��e�ʬ�WsEn��9}êl����ϯ|��n̶���yt[-s@J̾�@@����o��o�\��OC�mM�$�/tMhK
�W�4��q�!�����K���M�S��bFZ����݋��Ԙ���Hv��i_��h:1�.i��ϹQŶ.�O@���Ls�����O/�]���?-�ßIZ9!#�b�%�<�<�.b��j�����ȗ���9.ƞ�/�'�]�4��<�)��#{��5�i�kT��x���k��c�5Z`�=�e�n�� 7�V��bT��$i.��`w$�JN��d�a2�؄1-dB+�.�2�e�pdxG���6=���d��8��SpV�4!�4��-4xY�t[���A��w����{^�r�Q���6L�F.d]�t���@b�����/��n2�n"�Gы���h������������>�)���rs��lƇR_G����	��ʐ�e�?�.��3x������Y3���V/�lwجy]���Â�E��M�>�ޕq� �h��{��I�!'"蔹�oe�Z��#��l� 告�30=*��%�,ʡ��(�q���Sl�95������8��
y�r$Nޮ�Ss�x[�����$��'�Qc�t�Z^���?��Zu)lG���� g��i|� ;��3�-���S��F���P/`T�K�_��o�����}c�j �O���#,(�À�PǶ-J��W�n�_rc)�%�ym��UȒO@��&XƓ��&�P֏�(�)]4�vͫ9D�*���jb�x�xL��eZO��]�誌h.��4���ڽmm�J�0A&��K(��"蕺���b�����4�'|�â�3�sQ��(h�N��/��1�
~J�ʯT��W��q�}й8�o��WXg�x�wq���''��U��#'!�˛YI^�v�9�(8v@�6����N�7��ow��AqLGsn���PTo�b����1^>�#?c�EOa���#����������H��+ox����Jyl�(~݆ކ��${dD]�N�%*�W� ��h��	$�_Rsߦ��5��9T<�%�W�z2�k�W��bܔhԱ�_��(V� �B3�ӗ�����u��4@Eֲ�8���0��E���k·��!�,9ɵ�/Ng4����0VNzu�:؞򏆉�>�},��������p��E`7�hyo=LSC��vjAzc3�mY��is�䯶���'JO ����M�F���@��#���6��C�Gv�/"����@ܽ@�������o�M�M ʑ�Z(��1��ED��l鲞�����	$���y�C�_�e��וX�(�[��lt�?4Y|�6q����Ri"R�,t���X���g�ǡd���+���B�,��;�:�
������`I��og�7m����h?��!gcp�A6$`8��i4A����>&����$�*_Isrl�J8��%��j���bF�����2��*�LB�d=˥�̓=@M��dH!|��d�:݋�u����`ڬ[��� �0�9ET�T�lٰ�s8���^�׍o�{�L�)������q�aZ�+�{� C2��#�HQ�@ຘ��a%-`�j]`m�Bƞd ��2��/�.�ȫ�٠�20����O��GY;�Э*��NU��%���˗�� �]�Bl�H~����:Y��*�N��4xaƆ��5������-!��г�>6�D��w����;J��2�؅]Eq�_=��6R��nN�nQc*����O���>�ޗ���Hх �R�)�cPpZ�3�BV�ڰ	ݘC�a�ᖷI�U,���g��c����nd��8��
N�O�~�f@����Hh�����6�b�5�����\,l�����h�.a&�������PtF�x�;���뙦2���
�Is�^�	��ɳ_���V��3Vm=R�GY}���&I�	�)Қ�Ї�2�1F���8�k�aHv���E��OS������uq�\|:��o�{�Ng�C�Ҍ��?١�l3
g���Z�G��w���3DM-�軽��t���R��s�;�����[ �k��y%��m���a:}3B*i�������"�����>U8��[A��P	U�����2b���$�ཽ�����$�1W\�R�'�mr�?��}s�Kq q��I�n]������ASs�]vEX
���z��{U\���fD�$�;� �ǚAt�g\�W���:��	�e���HY�",�V���=)��#����=}� �.L�[?��71�^�V�����[��㱙�!�A�{�{�.��܊1�e\�1S��/���[�.-w��3��`�U����x�PQ0��z �q��͐�$�%R����.�TGw�5�+��~�5�[Wdƶl���ǎ�°p��ޟ�z�|Sh��̮k����EՇ'|�,Y^0��zd;�k���7	���pڥ�@�P�_lҠr��嬥df+F }2�	s�;	��0ت.4��dȡ��v5j<� �I��~�l����.���T�������m�,���*��('TJ�	��uVr1��\UX7��ʌ��+!qU����7��O�N��>Vƌ��B9����0� +��y�6_t��	�����H؝
șt��N>il|ATG��FO�h�q[�y���O�p��W����h=R��{��˨<-�|<�u>��mt�'jK*����G�ۉٵ�7�����S�>��T
HO<�i�0];�7�_ �������-ڹ[ߞ�=Uɴ  z��o�c\LPЃ4+N*�
�m�ih'��3Q���g�Z0<����e>Զ�˞ڈ�Z����|�cQ�61w��X�(�ʰ�~����h]��0� ���#m�sM`����
;�����p4��݉AP�7�42�2���1�6W$�񶔂���������`.�A�X�ʣM��_�z/�����P"��*"h�@"[���ەW7�Ѻ��*u�����N�����vIk�-���"�4�uz!�����\��t8�88��'����q�D�xS���� {�}�s�!�c68��c�Y���ֶh�c��䚓:ti�6�@
�fI����㦖�����Q�5M�ER�
��,�b�6�E����F����h�+���z��b&����7��Exx��5�������V4��wf��B96��T��ƭv.V>��B�\������y���}�cW<�#=�`�u^�Å(�](�Z�˓���g2��o��>��R��\��!��ug$��XAc6�V>8M�w~�
'�\¼p�L������w��h� M�kÙ3� |cn�e�^���E�������,���F��.>��d@N��=ً�P�g@�`���~��>��XP@��`���]�s."����4��2IK,#�Vt���[r����ѳ�ϱB[:�П*膛_*,N'��ee�L�*2F<s�z�QS��p9���P5��>��(�Փ�<�����%}=�wN�Lia������x��@��fI�i�1��V�1m)�͐X��<C��%E�E
��?V���(�܀Ť/�]M	�;�`�}�i=m�0=67�
L�8�1�.Fx�7���T�� �y59槪._��k2y+�P��KS�#�Zq�6�C�19�� VJ��o8�����N���:�{mɁ$�=�,�^]��a`n�a;�LSn٬���=_/�{��$Ö*��tʓ�B)�q# �LU�C�6���������or�5R��d8{��J]B�zP1������S&ؿ���pp!m�o�ȚL���*fW���/��%f6{`%4ou��G�bX�djtg�z��׏uu���F~��"�Rn�e?V>��ne��В���#�댟�Y��Dâ�Ȇ��]��/���������s)�\|r�]�r�b"�1��>˓�r"�6��
�����ۇ�^������"��њˆ�x�Z\z�P�o��Q�S�$KQ*�C��WJ,���)g�p�Iä�&�'���1�b�
*���=�,y��*��W�x+���+t�MC�4��t�_�`�2S���eU'y�{���,�'b�,d��eݳ�$�$��1�LIfxO�G{�uM�#B������A :�.�@�F��}����޵�;]�π��Q8lcF�H��svs	�������`\E�w��wG%tI�~��N4o�Ÿ��p�EЬ�� Ƹ!�p�wW����|�J�4����b2�e���Te���`zˢ��xр�����և�b�T0DS&bť�j������ި�h�צ�L�ܟ�w�AP��ōj$�y����Ee��[I��7����c<�(IZ<�_�!�P-�矌���z�}�y�N`(;1�N2���H�&�!JƨU7���n�#�X�"a��j���֓m1D���h	LZ�+���	u]~'�K�\i}ߔs�'0�iJv:���,l��WQ+�>��
�i7b�Dh��qJd�BJ��OA�)��8�������Z��1w̼��qew���]�/n��YB6mSG�1�r�/КZ)}�!��JH�5{�q:�!�1�c�)+,��4ZN��A7�Y8���D,g~�9KC�}G�s�ϓ�A��\(1��-
�kUT��Te#�Xo��5ɆP�Kn������m[Z��/���QDl;hB۰V�f{x-1L��t9������_žL������C��d�5A��T�4z����6t8���׸Y�4��D[Q��`-�3��\L5��LaF��;��W�b��[ս��:Dl�����^����$.ÿ�gM�ִ�a}Vڭ��I[���\aXY_)��h��tem���rSq�|��Y�v��N�β3@����ɲ�"e�8v��8?�Z؈K�8��<����ǜ��	�6R��aiB�L�ڜ~b<\�}��3���?���T�.p���I������|E��$��̔�C��Э�Ŭ��}-�J
�V8���G�VF>lFVM�Zk��z��P�5X�N��$�����(�87�#�Kk&8u#@���}��ėQ_�`�Ӳ�5�=��͞ �B���=�����3H�[�#!ur6�q��S#w�O$���=DTG}~ō9��_?���h �q�\� �4v�k��}��?�$�7��Lӆ��`b�ե�(�;�ͽ�e����T�9�=Y���=�gu��cxۈYS��Ze-T^-���ïaTG�C�פ�f(^��$��P�z��sTބ����w�)�/�ĭ̆gc��c��k��4Ft={����:� 7��Rc��к��9��ːv(����KJ�e�A�]<������%3%~�m��A�q���QEZ��B���O�yX�sP�N��!PnM׃d��6����P��c����s��3�|�\'*�jY�LI�|�;���Qp��=�5p�u\#�ۄ#���C/������Y�ΰ����]�ʾ�#�	_�׮3���0�El�����Bu�u�\�}�j��?iP��x�韜_5�D���K�@��q�&�Jڝ����P|ϣ�f�g`l.����,̬K#:2��U9�_����Mĵ:i��2���F����T��zD�4��j$X�e�%Mk�Z��٤e�����ۇw����G@����Fq��4��8���D�i>t��{�=E\��[�k4z�x|ޞ�|#����?����s��g�� ���u�I1�VɁV��u�u�.�b�Sdb6͵ap�Zlӈ?���j�"�ff35f	��?�����ϟ��$�U�i����ԣ���yc��^���0�'g͵w`3�.�P�-[�A�2Ydb,N}]_h��J�z�&����pS
َ������ �V�C1�В��s�e�Bnߥ��\=d&;dz��!�G\��5#��ʻ!�ǽ٫lS�"����3ew����o�9_�.�K?�t{֝�#�YT�Q�H�LF̫&f2ì��F	_@�|��e�����6:��CV"���e�4�g�e��7���F�ϝ��j�
ߛ�� �-�e�.����cǓ���X:'9��F���:�Q���'?���g �k:u^Y�b���Mۤt ������\�D�]�0�1Y,��8i�Wߧ5����,-f�@f����g~�����c�<���}D�Aj�G��3���|g�&f�;���GՖڟ���������e�O�k��c�K=~�r���:����K%���s���*���1wz�.6i�9^���I�����U&�ɳ�t<��6�.�|��Y��5<K{|�灭���Z�}H�T�/�Q���������p��-��@2#y�`�6'{�s�?2���FJ5i��m'$.ّ��bihīԥR��������-�M�E��45�G	�fYQa��t3rM�N��A��F��#E~�vq&.�Uct��%F�/�����'&�����LП��~���p#��Ѣ_:���B/]�Ì�"u5%�\��@as/8����hfޠ��;X�A�2��Gp��.�I����?���_�/J9Rlך|��n�ٻ
n���L�&,8���wңt�
�#Up5�P쮤���a[�
l�ө4�/Ң�6�؄�%���,.����!֊Y-q��;w	���xG�����Nj���l*�7#�55#�j����'��Y�Ɲ�9��#)@5��}�'��N{��i����)�>�_�:E��n�P�!�z�T^Mv0�Ph_�su\֗�����Nf���.�I
��'��J��#��� �2E�oQkf�"��G��bA}.�p�����Ap�L\X����.Ɛ[���_n�sܦ^�=(� �3D��0�y�
��gJ���/�:***�9���;]���wM5 ��/"��S����eȁ�=Tg��Cp�*��F��d�Yy5���Rx A�℔Irl�һLC���٠8��w���~�l=�c��kPK�<�O�^b��)��3@4ŎQf�*ײ�.3�$~��Q�'�}p���w�73�0|�26Qb�)V��7sb���D���;@?��G��RО`��+.�q��_�R�)����ZY� ��v��v5����A\�}M����;����ͳ�mŌ������H�H��1:x���9�E˲+k���&p����S�y��\�%���d ?�D��6��N�\��5�8���0�{Gcg��\vx�`���yY�:�ٱ�2@f�!��e>mds>8 ��͑�p�G�~� ��\���KӤ�bqퟮ"�(��%���lD4�JfW��0b���=gZZ ��v�k�9h�*o�}!��r#+�0V����2�޺RE�Uv��=��i��J7a���3�U��E���,y�ӯum��6�MQ0~�����6ͫ����|�8�����q�)�/*Uu'�f: �m�W�L#L8ԩM��F&��i�8����v-�����d6���{O�J������ f��~��N��r�J� �r�m�;h�c�]�X�uW��y 4?{$+Ӯ������t�s}YP�Y��n�a~ֽz$�e��0["t���z�-ɧi�r0�ek7�5vT�H|K�-��,�l�;����o��M�{�@{�N�����` 8lk�1p-U.�{S�,��7LF���`f��k�[����L�Yvmr�4��(���cZ����?�W"k���^��2B����U���sg���`푹���{WF�����2�v/Ϋu�~��lC�-:�SA��i�d�O-��G��<�0�%6���#�~'�C��Z��ʓ�������z��Ԙ���军3d�0�(k�(�t�8�Y�D�:�|�G7*��<\e]h֍�*�Ɨ�D͢=&���ˠ.5I����&��ƌ������V@@�G6(��1���#���Wq=TyĭEs�����\��U_��}EPw��_�|h��[	�
�r���������f�����"p���y$+њ��#�8^��=�����X�1�'��A9�󊮦�Nh�5�Zu����0>���`�b��]1c4�Y���η��>�#���Th���������T4ֿ��t�[5�~�4n���o �o�g'������)��g�ձ��ܲذ=�����~�1xY)���S#�� F>��9~���!�F)��c����()����2h֞�}i���a�-S��m`I��3}�p?g���G�����j �^�Gu|�KP\ Zw:�9����&E�:~��_��-,x�	��:���Y�S��
�j���l�r�� �t�����7��2�:4�q���1��I��v|��IM�����'ʔ�P��N����uC�0(����I}^l�U�G�@>���p�)��M�|&�Eh�\OAX��\VmH�
�����
 o���d~���}x��̷���7�i�yq�ٺ�d?4�
;1Xt�N5,'&�&���3CҜ���"���܅��KH����f��s�É��/l�yi���5�B�O�������ݺT�o��6]̐��w��yP	���Jǿ���>"A��oԡ8l��"�[M�ޝ����Y%�d(��-�x{Z�V"WN�xv.-�F�����_�o��pIyZ�ݵb�y�\�Dn_�-f��Dtךgh�y��.zx\cx?��R��#̺�*|B�S�NՒ�d63����Ǘ�-O��H�iDRK�(]�����刎�b5P|�،�Ǽ�)���񜡎�Բ�׻�Tڬ���6G�oy��J)ɺ��D���0x8�lD$���u�P�v
Q�<����S8�����J���80�HÅMBQDX���qgq9�:�����T��4		]����= �D򠽼Ug�ȵ��]�Q9�EK�^���7Y6%n������U���L�g=756L,�/�1��z�Y�ÿ��@�"��� ��S���bW�T�����ٺ�#�8'"�|��o���#?����� �'2����������b�B�w��^\�.�VќPİ�ٸ�}/���a��!�>Kk�W�A�T��g6kP�X�ca{w���F�2g��Z�Z7�G����V����ըbR�ʢD��7�$C~"J*�}f=6��D&|�-�8�@��Nױ��>;�g�#e�T;�~J$L*�T��E�f�Χ�e�G|X1��k�I�	p���� �T$�����`-̰��.�,x,��i�U �E?3��6�pWoJ�W�"�����ߎ�����Ek>�W�{]R��u�;��>��y9�I�'���~�Pbǝ�'U�R!f>8�ȣ����ƿPb��lV���8lE%�-s�%Y���K"��0]�D(�BHaC��e��
&�<3�x�<k�ӧ��W�� b=6���P���丅RUm��-LsH6�)��h�*��[Dж'�����A�7,,f{Y�'ˁ8;Me��s ���[�&Q���,�HށQ�6�s��|��@#;��?���M��<N����W�u�S��xu�f������֬('冀��Kk�kglCT��1/��`|'IY��K?�/^��0��]QU(z�h#v��A�}>��j=͗X����$�����T
&9��u-K��L
{l��y���>��o�LϾ�c�V6�aҟ�T�A�����`���u��"NY�tVyF���*�l�1��?��[��J.#��ף��A�a��#�F�`�o�H'���"e��Rk֊p]Q}��l8Cg9��N�<ed����Q9�J�P'�a��Swv���*(3�	��%��0���PٲE�S��hWhs}a�mع�3�X&���lY���7�b��AӢ�'����:�ص�����Jd.�����.O��I%{:����"�zp�?ܙk����oKY��Q;yiC65@9���[�iC�����^�[�o�K0��F,��ƨ)k;C(>�!_J=+�A+���_���ug<?�s�>������U�: N(��8�D�� ҁ�|'	Ky^o fVP	��G'ʒb�7ǒ������������i�㪚���6"$�e}����/��I����{��[y��!�ݻ!��ʋ�'��M!�]�>�.u��/l��V(��7lD7|��Ě�u���Z�@�ι��]���P���<��p&5}����ًm8 G��7ق9��RUKhL��&q_�36(��A�aI����K@���ˁ3}Υߗ�X�z!�+`�����ͦ�}�P~sU�hhf��	Ѣ����B�/k�U���t�Ed#Y��135B�(kA"�b�@g�b��oa�LY�CYNK�uQ,�{�\�󁵂\�����sj�b�H��H�_���U���7��D.���ɖZ�}'�as	����ir�DP�w��\B��|:�]�F�|	�yxrR���Y�AK�J���i)T�+�W�RJ)���\��l�7-�	��Dk�Y���x�/������3��~1	ߊI�3�bes*�Կ�ᰵ�R��0�L����Dxa�YMy���w����`�o�x��U���5\�Y:ŧNGH	h�g��^2)M���F�b|;��rB�{8�C���f�Z�?�eE��.�z�3�<VXy:z|�{8ґ��񉹙Z��ȿ�H�����ш�$q�؞t����>Me�Q������ú̧ z���k�ǲ�qv�ӯJ�m�����"��6�RD0�"��%�l�2&j�XN`��Q�mUlE@�:T�Lw�G�>!-�T�ˣ����#�Y���$�� ���	�#R�!�=��g���q]+"��'��;� ^�qkE��1�
L�:r	��ߐ�+���2.��9��b�0�����sXuէ��(p��c�PE��H�9y��f���#!Y>Y�u�F�f+�i��X�*����{�.��>#u��/u0��|YNr�o0vpj�;铱�����t�)e��oA
_����8���Zi^D�@@F��Gٜf�ų^�'��_\1A�q_Nd�`IK�~��`s��>~��Im]o���hw�������:[���pD������"Ԙ5v��@,�B��O�'�����j���a���V_w����?4�,(oM�v1	3[�c+w4���߂Z�ĂѯMr�TX������T)r%�H�o��@��ڻۗ�ػ_5�TBC:�D+A%����v�Ĭ�ؘ�a�P�Ơ�E�s�R	�ѝh�UD	����T)K\�����3�4��(�
r��"���l������:&��$����;�	�����.��� Vt�ͷ��5s�S������lU|7��?:�[Pw��ѧ ��I�IL(�;��p����ҋ�y�XZ4M0��t�E���-du�8twyI�ߩ'�M�����������yD�KB|p�	�ۤ�%�1hE������OC)R��e���%�X���%]�E�ڠvw.�w��4�_&���P[�>�N���ɐV��v%�׏�B����So���Vw�F�A�iB�ĕ�Y��k�u�5�`�?��#�B���*�o��&�,�4A`����[��Q�˜q���,h,�����Q��0bA}�@^�f�1�>�aOg'��%�߭��\��}Ԣ�z��?ⳤ6��?����^2�OG ��}�ߗ��<�GJ�	@rN	����F�D�Q�HwE�v@^�=y�1Cu���ij�`�#M�Oz��kV��oD�I	�[��u"s��c8��S�-�#�i[]���h<
�ra�T5R����(���48j��JUB��t.�a�	s�D��r�m r�߈��������:˛���5��5%ۖ�Ϫ��6��f�&ZMКO�+L����~������>K�x ����az������D�A~�ߚ	�f�����1�m���9+/�D�T�9�S��F$]`����A��������l�SC�[�@�~?>��ea�C=._�R$���	�#(*���J�9�(~羁s���6�L;躹$�8��N�Ih�������	�o�n�&~���ʠ�V�mqlR1�$=�TB���t�֐��La��M��U���H[�,3��TM?d-_ƻ�w�$h4�K���� C�4��k��������!�V�@�D�a��u�1�MZc��na���Ke��Y4�[��l�k(��_(3/�^��T��3���,G�Hdĵ�5m5#�+d]�(7F��<�F�!겱�vy�b|��q]�n��Ǉ	XR�F�j�W�0&ukO\<6��m ��n����3D6�c��4�$2"ߢ���	�[
T:����c�8�b�ƾ9�}��fΔ|���V��N��y��7���\���O�r��!��xk0�a�%������(���d�����rLT�����	s�?��΅�fd(��'�?SqX�-m�0�DB_'����[��#��� ��3���G�c�Ė3ڿu2A�7�v�y9�^���^��x���P��5Q���&�U9#����z��*r��0񧊵�_��2zt�X`��/��z�'���2l��OƱ��𚽈��]`j�g�CwG��U�گ�6�b�,!�k*�C��'�����UǗ
��X�Ħ+�Qy��*۹���bkU�ڗ`��И!��8�i����>�-�͌h��#�h��L�z��{xk	��^&���,j�$�Y�uD�N7s-!
�A�G#r""�2�n����A���5�����RR���	�5��M��Wd���2�P�����ƌ~B$;�IEh�.BY�ʙ�I��[����J�ȑ�,���q�29���]��ń�D��`�q��Q�	������.�{h~7�#N�=���l�6��	q��H�m�{<^ ��k^ǩ,<�V�e)��a,u���7I$�gT���hD�����wz��4ӜB����$�cغ~�/��p�L�+��Y��~�K2��w���[U�\���ԑ�<�.��Xt_^!�:E��O1%�H)�:���r�bT�2ޝч�$�����ع�^��MDS�"Q� �o"�Q�IX�Ӿb�����!���E��WT���:��b�6�w�A�ۦi]�0��V���X��_v?��4���I��N���z�/�]��/�������Kt�X�<J��H��m� J8���` 	h��»֨��ti?t'M����w��NW�-9]�}�����L������:��aA8V����e�k�X�h�x��5���t|a��8Sc��Y+�m� o�Ӡ���s��b����3 o���C�M=��Ny�PҖ$6�oư�3�+7�_�h�tO��`��99�&���{�v��XsWb��.�=�� ����`S�,Imp�l�Q��@yb�-���R�8��,Moe'})c�/-q9���1
�T��ҖK�C�$v뜻_%�����l5z*���F���6���HJ��U�P%�u�IE�E1P�v_8��¶�+�/�^��TwJ��3]L���D�7fI��N��������%�J"���Cl��y"*�]C��3��P4�5�8�W�ϸ.~(��9�q�4���ᓙ,'��趠m�5OH�,�:>u������n�� $J���k�Bq��P�_s��5��<]7��U#�^��){��Q��csI�?�����!	�Z��ڶ�]�;+.���=��a�:ܧ��# N���x�~�)CL�L}m�m�@��:���<��+�V��;��W�_�Gg��m�h��Z�MV�%#x�|^������]9�;b�6+����׍�� U7������Z��OhY�
>j�#{�ά�ax���vU�+4��v����cQI|;w�c��;"��
��TVBÚ)�ޓ_���fROzȅ8�F%֍�ɳ�/�yP�z~��)���g��j2���Nde���6�}J׃^qw�3�:�K�G7$u_�#�b����ƴ�
FG���뮄~�j�D�ЪV�e)�L��9��r�H���O��E�-c�U�D!�!r����R���|�������L��M�"�7o'��nE���r5�ڳS@�y�s�\���u��뇳+�Jna;i�w�*^�>2?�K����;�Z���ݓ��WO�F�LE�㒐�u���&��5����%��r00���o�'��P����q��n������
ѱ�1��0K���x��;�MZޏ�∢6�����x��/Gn�t��1\����E�������y;��7�|�H�F��.�������*�b��mn5�O<�}��A�	�.��[>yb����6j�B�̳��QH��j�yN̖���ۏ7c�E�
����G�<�I�a{�,�o�ըDu���A�K�U8y.�|dDޭ�F �����Ĝ�PP)	�?��I��m_r|GP��UJ��</�� ��?Wҫ9\:�!6�g��P?�G#S�O��x#�3%������KA ~���pP~�b,9 N��k�p�|t'c�A��ʋ�� �^y�3�6�i�Z�����c���=���
%r.�]�I�y�=q�|�����-�4������`�6�`�� �n�TH���I�Đ|AW>�j*0��X�s� 2��o�����C甖� s^a&����lɰ\�$nsy�UW��En���0L+sÖ.���Z��9��6�[f��<@Gˍ���?D�ڶA�z���硷J��E����F�1ӆ�DD���=k���Ԃ����ᦜ��9}��G�wO�"5^�G��s#����Q	�	��Ɲ��\���ʗ�x���~�-ێA���vާ�T͍�+	y6�b�\M����-J�zb@b;J��� �m�h�}�\w攒L ���i9vc��� ^[�9����s�ס8�t���P��Q8���gMl�{�"l����=T����d!L��%��-,k�
&H����lE�)� 0R�1ˎ{7D��kf$��î'�s��,Y��pٟ�.(=:��T�q�}�b���S��v�Tbq��K̻L��]�A�[AG��[4@��)�:tmeo\u�	]�������M�_�ӫ����/k�v`NIb�����&�|Zҥ�n:��$%R��HF8��R'?�1�A�����_M!��a}�w}��@���pfD����խr�(pD T��D�/��Qw�J��<0�{A��W�����o��?�0�Sk%z���kw����C��4<�@6��f3�Y��rF�Q"��&:Q�j-�C~��!��J{��j���cɘ]2�%l�|����̵~u�G���������5�

.�u��sf�a<��ܤh�ǝےկ�1d��f�̺���=���g����X��	v��u��/�ǋ��з�\���xw�(�7�KDڅU͟�̨���o �,���u�aT�l<6;�Ŕd�A��kceD��D�����+��׺z��:�yEk�P�X���<�z}������Nv7��W
B�I\���"�Z%=�X���pL�zd���LA�*%l{]�mqK_u9�� Qᛀ�Q�ݤ�
�-d�1	N��� �IO�2$Wax�bT۴>`� ̝�b!f�{���jSx����B�1�l}�8/% �Pɾ����v9ex�&��}Q���)��0)���#m��!q8_~l��^��W��F�T$5�6$Ug/lw2Y�����wчh8<׫a �:;����ok��~�AN/����Pr1]��p��z��NtO�uа1�O 
_�I8���\ϴ(�]�i��[�.
vp�޵5N��F�� �&7qO��8e�W� ��E��7��LF���O�Pl�Lڔ�]9�Ԁ��9r2d/>L�
�2�%�����m�c%��~9YTmZ�b>j-�"9��ө6+\�kl� i�p���j��͛�D́����!e��C��ٱ[k���ԋ3�����}yqQ�R`�Bf�?^"9��(����w��,k�]�^k*"�i���ӂS��ܚ����A��ɥ����@b1Y}��<����3F`u+�J�0�y��a.)�
�J�A�f�Z�}D����1˷�/�h�?�5:4��:���"܍�7R�^x���;��!r�6E����%J���0������k��(�}�Q��,�+2�n$L�J�P��D%�l|��\��Cj�+
<�w��	��ظNEQ߭T�Ka�Gk|Vl/F�x)�ā�-譒�9u[���az;�a�7��=��4�Pg�6�mB*O;��bƆ]�*�gWr�ݯ>�ҘL�(�~ۍ��ܗ�H��'S\ֻ
�� �?3}�n<P���N�'Z�[��{a�����_����b���"_rVt:k����x�D@����j�p��;O�J�>�-.2�������O�����Ap��v(�B��z��V��!J4�Ŀty@��挸��ӡ��ܫI,�xB�`"]/4���d
h34ű.!���!�-6�"h8�s7 ���Ē	)a�3R�K�-�4F)���-M�O�<-�� �>�U�m�&��z�:z�������(JF1�]t�K`�ˁW�sNpbY�0�k)�H�[*�p7pnY�*��9��8s�wc:fk�e��.8��d��Q�F��� �uJ%���w�����X ��W�1=(ogp�Pyw��;ۄ˨�j�(eq�j�� A���
F����=�'����u������N�=�z����i@����;*�Xۺf��m�Y��;���#v��������E�f��"6�5����:t���D��W������+x�$ kȺO/(��F8Do[�&���b�g����ߒ���3'cC���gϞ�O�m�،�p�
�"�Q���z�����1X�4��N\�2 
;�������8���
8��}���u	`���mw+1
h��BlA}]Û�1깊�6^��<S�'��S�{���f�K�0֧���ͳ�fr���j�?��H>E	�i��6�T71��ѐ���5Fh�Vڢ?��V�ؐa�B3.����z[c^&k|�-��EɞВ����*��,��hP�$�ޞt��#�¯l��j@�RR�ƤUL@���?���������l�T5I��Q#>F�2"/9ͻ �nhH��T2x�!!8��GU�9űȔ��7dC򆚨n�=�P¦lX�t2螌������[���i[:�%��f ��_U�W��5����S���/5� ��sʽ��3�e`,>Z�V��K��2��=�J<S��
o�����&t��]%���$!Ib�~6���].��S���e
9���ɣ�C<��pŋA�����w@��풡�
��1�j�hV��*��a,�|�E/���bQ��	�NZ��k._�P��\���af��3(J�:F ��D�F�&����os��K�8��Wg�>K�J��_k�n��W7�f��f����*n`.��g���B��m����X.r�Ev���oֺՁ!��b�&,��Uꫠ��I(橞�:�0��2�X#��ݦE��T(Wuh`�� P�(���<�l�EO��WU�'e$x�����]�(>����5x���l�/T:�
��g�f�ޚ��j�����r���LU�8�\[ry�]3�"tձ>�CӮ������-m�"$�U�<V�P��"��C['96�g��&F�WGnH]��w�i�. ��=�u��(~�ÿ�~̃�]�ꇊ�V���ma�H�f�d8�oO��c��s� |yZdH�̍���Ȣa�\y��5��/V�P���^�.��q���V�+h{љI?&���\j�d�>��]W�����%B}�_R]�"�*G������{��0 G/?~a���\��饋q!S��o�N�
�G�)�E���@��Cf�t�����*8g
�ƃ#e�9vX�X�f��ѭ�Å9��^��6䟆u�o����|�c���ڼKk숔�+���qb�+w�}�����Qaۡ�/x��@2�vt&����<o�/`0����%S�	e�0}�`&�!��_��ԉ�ش�B�z���x�ܘgH�"]9��{����kS²�*��=~�3.�l��ت TD�5]I��h�o]�sY~�A�<�"�Vq�9����*7���`?G;N�M��0�|��`6���ʖͣO��e�H��N]����h��eM���5��D �J��Ֆ~Pe��C�)MxZ�@]n�2���Ču��w9[["Pv�C��0	�wE�8.��)S�!�l���Y�m�lb1\�4��iT�.�'����OY��z�3�؁��0��w��Z�g`fp^-�a|m��������Z���f��H����a&��-]z����TNV����5kr/���%,�Z��M���Û`�eľ���jyU:|Na��A���Ǝ��Ӎy,~�W)��$��"�<
�������B鸗sP�#�nl9��z��W�A�׌�l�Y��?��^�GR+P=ϯ��)1�"ya�Z[A"n�/qǑy!�h�x��t[�x>S�O�d-/�S�q���t^e��-���L����p�1��ǪDro����<efۋ��Խ�r	=��=�I_�K6zؽ+�։�YxX�zyx�^M�FUSGQ�u��C�Ԉ]��L���/Q�
/����A�M�Ac4Z�[����&�
�L!�k�3ˋ��Y.���G��D��jS?�)gDW~w4�W��o��ޘ���l�09�6BO�W�sh�[1��A)����aU�fZ{�׍³ �{��P�Y$��KaLN����J^���>E���`W�d ����X��րi�9���q�HJ��Q�a�@��t��fV�a>r�i��ʅ�qs��i�lgsr؉���}�[Y�� G��5]�W9��rW��'���2����P���!��"z쯤$\���* ������%��Q���M&�d���,_�
G��v�eQBw!�|��6ٛH��Nݭ�=�#/I}�6�.�+Wܪ>���m�"�D��C��q ��B�c������%8SՍB��	�_P�7;8�Z�:/��xP����%E��:>�D|��@�K��c$�ȱ}�ɍ�J�}Z=���M53kH2�dD�J�w@G�\|L���N��4�R����Fk=�h�%��WӟL�^�-}ƣfP��yi��X� �i/-g��I��Ў����P%��	Y��� �F@ٻ4�6U����:#�����m�uPpr[�UQ*WȜ��$��n��=��q�˳8f%����r�!6���M�Ym�����k�2��G���
��P��oE�a�R�H��_R����#���ҵZ�$�&�,�	tu�{h��6�Y"-�>C{�N��/����]nj" �JsI� �R�B�K
���o=v?�1����o�aH�O94��7Ȯ��>��+.�.7�P3��kسm�|��e]K�`�?��`�tǭ]�ͼ���XuGd쎀�
8�P@$�8�mdm��߭��d�m�whc��Rw!"z�llnuf{�%B��}�S1�����8{j�t:��h�0��|�Dz�Ƕ�ʅ�@����h2g74%#�C?��۠;Q��#K���#��H��"�>�vl(-aE���ɔ9�du$�k�Ԉ��A�t�n��C�c��t}|��g
��S��)�Vf
lq��/VǄ.���J�I0W����J�\�~��x���\�4^?��Z;9q=g�،�� dv6a0YAW�9A6���18}y�RE��r�_�A| �6s{.���L{H����=�s�4��P�x��u��^2��M��N�����f
�Dy���@9��I���E%�fh0��0%�Ǚ>�8�KD���x��i}6x�%>7pp�p\��h�l��p\T��8p���������\9����6l
����]w� �m�z[F,����		H\�@���3{��Q�đ,?]R��y(V1r$�����Ny��Q䃬�}i��!x�R+v[|aː�tX. ��=�L��`���(�_���_�asS/d��W�����J���7C�+��q�	D�޿z��.	<k-��増2���|֏�Z�P�)���c�)V�0�H�2��w}�`��.0)��N.��yrK���>�*Kl��R�1'��h��舼.�A1	����f��!��8a~��5�P�W���=֭�S0��#�*J7'��p���d�$�&�D+�cc���ׅ�_�������z�:����-�9x~��N
����/z$1uD<�e'�*dВ�j�xF�,,J�vJ�*Z�&?�p��/��,?��f2���ԓ���U���	�,�H=�ʡ�`�ɨ��nٰ�f6���Ko���
�JO��"��7�6���"�j�v�'�s�5+9��%��7�?�(~��[���*ۍ�t'_�<�7w���w�Ti�|`���q P�;P�ć����oֈ�N؛�s��!�B^#�ˍO���j^jC�Giv�&}_��2�h��zG���悷x���Fh�e���)�������t�v��[��%���ɴFů�&��ϭc�g���fx�n��Vf�MED������Jb��ĸ�@җC ��ˆ��婲h���܇c���Hh�+f��)����(0��p��Alf*W~.)�`s�f�r�$,�ꍸk��볠�.^g��K����rHG"�4U�-�+5��N�(����U�k����
����ٿ�?�%��<�a�ثSC�d�F�7"��6���Ga"�o?�>��B��_9�3��8k�o���e����NoZ��#����cp֧�xB�_�;TK��8���k]hY{��OE���dE� X��|"W�-�#�냥���2���/���H�I��o���\]Z�����8��[2�&�_���7��&�W�E*���9�x������<��$Z!w��&�I�\�44�� p�z��S��>�J�0/��t������ܯ�s�87�5��п��5?W'{�l� �솼�m�"�j65��.,��FD9v)����L`L�&�=|2�0j-���E'��t�*H�>�۝�0��r:ԝO��nEl��_gTv&C���bT�?��Twhfg7�3%J�h!��d�Q�#�-lQ8����5:��'��uk��%.*�P�:xRX���4����
+AY�M�9���m��Xqu`�E�W�ER�G���v��<B<B��v(ع����Uu��W�-��.}����r�^��׭x�/!�%z�Q����Y?�z��f�᷉�A5U�[��=эEeQ�ӿ���=*oї����wM���/-�J�S��kÍ���A��8��8�������<=���!�5SZ�?�An�o�K4��7$V�Q^���Gp���i�B6ꋆ?�K'e�����մ��D��[=��<A�-��B��3�r}��{�� l4 y��͂IEgO����Z
�X�^���$����wD$@��u����,�T���l�n���q�'m���%%!�io�����C�'�p�Q�](D�ĸ�5�6u��k��1�E�Y�k�$/f�1T�+v5:�0fॉ�X{����S^�?嶨�T��:͸k|���g�qF4�̗;C
�{��e�Q�?4� �F*��h�z7=�3�[�`V-��W��Y!�J%�����ptN�9ZW��r>�����h�B$2+Ao�`�:�Qp���1ɂ'��z���af�o�S�#��c��8>m���1�L�J���ܢCy����Ix�S�>r^���6�a�#�K`��s��_�O9��K�g�o�W�6KP鄠�r8����[!)�$�/��!�ͽ,}mB�+���^&`�6UM��a�P�h��6���Ѿa6lC����A��yU��
n!ZT��I3T�+N�r�j��ڑI���&30��;߆����w턥~v���j���#��3�B
�?(�
l5���al�5:�-f�l�M�������Q3�R�q���y%I|�Ԍ7N�O�Y��Nc|���`xs<`/�f1� ���2ݨ�־wEC�� 6�|�(r h��q���b���t�Ժ@[�$	���I�ό� Fg�P��/E���Q��+���������߳���^D)�}܊������^�e�UpjkdX�4Ə�׬�Md�m��A��inz� ,e���.���fTڵ �?�7Țs|���`燣��E���@�S�6ZS5��/�~z;`�f.�z��}�AY��-�Z�&�lk��]��cDǗ���ؓ+I��%�ڎ{U�La�z�J*&�5R�� �~I��	�
,��w���Z�2\����z�6����R���[���=ac��:7�z\��E�wPύ�y ���Ni��: o�2�Ж�Ԣ~�*�03�*$y �A�Fj.]�^>r��a�̢f����5,��o����"^��k�4d/-l_$�H��a�(���ˈ����2p����%x_Y����l!�� K���8��Z��`U#:�WCm�z?�[�i0�N$�� ��}�H_DGSk޸��KL0�n�N��o����Ƃ��p��+	�I�{)���'�%$F�BV�C(o'dF7�(�n�4ܢ|���kxM������e!jO+x��|	���c|�G�C� "Y����/ ��s���&������f�-L_�+�RU�aeP^U#k+����ˎ�l�K�ǹV�I�B�7���YQ)ֆ�v^��
�S�,�u�?�|�.}�U�c�(��+f��ϝ�`��|���{®I�135��$J=��oUj�$�[���:�VH;ʜ!��F$:|�[{���[���鵊w�}�#����9{�J�*�|� ��l<���%c��R�n&�������x��G�����9=k��M��e�&�$%̮:�T�ܫ]=�����lVFC�$���9ȶl�@��_h�]إ ܤp\�K\W3{p	���g����Ёx����h�ެ�P���������5|0���K�ꉡ`��{ˇ9�z�4��l$p?e�����IC���V��X�Cs�]�5a��t�% x��o���JeZN�OY�]�?�CYR:��G%с(� um��������t�͛�����gIG�YDm���'I���8ew�Y*��}���%A���*��?����2��QJ���yL��kGE��2�S��L#a\�֪g�o��S0��L:��{z'�%��ek������o����+����@`M�>Ù�����iT:��4�ȝ�QE<ӘYVŁ=q�6NHp��B�z��!s9�u8��$W!`�k)p�����j/<줴! �ݱf�_�<��=�6�����P��_m�VfTX��:S��fT�?��0θ�C��ƂN�����j�~�I�zR��j����[�������I�6�N��� h���ŌO�\C���ݽ��������<`l(
��*��ˬ-4�T%Y�;|S$��%aޣfzY20�*Ղ��C�Y�bR��I�� fD��F&�U�M�4�O|i�]v1��3K{���d�K`"l�V�S�:�O���R��:L���c}�QՐ-x��Χ�bk�<Y�lܡ0o9$���w�"���U������0�kB�����+l	v��ջ�d���i֠�b/���A�͂���9�3�[���/�jb,2n���v8���n���o��/a�XF��Q?	�5q�ÐݭYLeD"� vO<W�G�`��+a��)j��;/#�����y����� ��?�*�grD��lP_�g�>q<���f���p!��1���B�����D�w�
|��$F2Ԡ}tD��f7�05͠�m>��k�/��Y�x
�Y���C��n�/B*�`� P!	�'#	�5��	���!Gr ;���~��ʸ-ƞZ �`���٥�������H��QB�+Q$���25ױ�\�4ƈ�,P�?s�b��q��+� sg��M
������Œ_,R|Ğ�;��%��@P�X�������`q���>�}�3\�M;Js���c�`9LC�H������rh�M�G�ۑIEW��<��@����mG��v� �r�6������^�`8f�j��<�!�d�\;���9%H&bC��\���B/�CO��/���v{�_�[{��
�8�D$������:}
"��Ph�x���vd�H ��,%�4��I*�B�$_�S�Xc �i�V�J���ݠ�q#!RF'�ڻ��y��wPs�hdS�!/�QBӔ5��a�kF���Z�Fk&83��g�	jW��1�>��)���B�&�e�As�/�T'�,Lq�C�N�N�h���كakw�6�6�Z֩E�}���3��*�m(��'<��m?
כG��U!9(�������>��d}G���)�q;9^o�gM�*à�C�q�a:_Z-oW}ٰu�0�V}|{w��i,=~I/nz_�a���<��Qvғ~�����7�F�ºh����.9-�z�H���8�C��I����$��O��bv��"=Ng�u��>�;e��
l*;�^��RL�_ P�t��U&����ʮm�q��c�����@/e������C�������
��o�~�塲� 1F�/�Ԭ���j�/s+�[tʔ,%�h�i	|��*Ii����W�Ef�����9\Z7 9������z�PHyRĳ��|��Yy�,���4S`���&`�����ĉΠB�!�����ã�}�����3��R�vG��1�����o��pz�a� V���P�敋��;!���,>%����ڄ�!n��Ej_ȍ6pHX�b\�,m��}�_�����$�l3���zՄ���k���w���Gc|�ň�?��c �)6%������PA����K�^ƙ�.��<�!��"�W%�*����ߓ�]e���1��URxz���o6y�����0�}�5[���P�P�K���i��X�s��	?�1<%�Õ��:Dv�����������	{�-���jɲ�3�j/�4#t&⦻ON�K�SQ��̡��r�TŃE51,�&b��[ک�O�F{����,*�38�b��W���8�	K��#�����CWn3[}AFs�N�;�5�v����.���e����R�)��7I�vqv��d+y����ʊ#Р�Fz�x��ݕƃ�S����������o����-����&jS"H,l���xy4\��{�I2�U�u��\W�q��������S�8�y9lL�颣D���Sv7s[+nt��T�Pd
R�x��[P:r.�L�k����l�)�ֹC�&�82���S��}E\�3��t�J�tE��vZ�ɇ�1��9l�c;`�1�I��n6�p�(Ұ�e�BP� (RH�������`�8��ŉ� /M��_��	��3��`5�G�BBD>'���� ���Ou����̊��y��d�I!i�������b�WhMvM\l���T��9�X���.%2�����GG\��$Y��#a�v�C_���'�h̔��Zkx��,�t�e ��B�	p�FIЭz&Ҙ�K�%�k�����`�����\���|�X,t��u�\�;��}�P�$wK=��]��X	� ��X�#�{
�����6=����g�{�[\�Ƈ��^w }��R@����ŋe$T�q\�txS4mDL��<n������v��*
z*��Uw|s�����s	'�Xz��fH%��A�����e����{��.�R5��"}����k��S��F���d$�-������P��B�YeSC�mPbI����+R���Վ.�q,?�ծ��{ʠ�*�6=��'�eg���ĕ׺e��T6o�W�[�@U�������2�9�F�b�pR��E�w�\��S;������,q���h5<̀N��S�T�b̼�pS1����l��uCx��Lb"����`J��	���/Ԁ�Ye�R���N�v"�#Fk��?-rw��p���2�������3L��<�1 }����=[n}���.I�j�S� FyB��8��(�4���+�ƻ��?} �!E����/� �2C�Eu�����bHQe��8�I����^�tV�P2EޑIZ�!�(!�3��к@o�̊�]�����An�M+���mޔ��Dh׶v$:�a�&����+�Zl�*e��N�>#l��;�A-[�3.�n#���Z���'D�YwѰ��U_�7�lD���y��}@�F(M®�����?��B#a�։��2UDR���<W�F�&�Kl,b��M|��S�֮�e��G B�uT�]�Y��s���B���Ҟq���>P�V�����L7�@뢍����+��!������&����Ȟ=d�Z���V�q��o�J�lH�N/�H��A�� �����ꚉ3�%�߃�	�D���DI9����[*�:U_� 9��I���^I|<OJ��F�7���c�Ye���e>et`�&z��%��]�$��8����_��z �ZR�q	� \m-*���0�jL�o%>tUQ�;� ��b���`�\WC�U�e+��:K�pYq��8a�>����Y����@EFf���m�a��V�b@�RP�q����t�x��ى�hn�|hN�(���-Y�ΨPT���\}�����J���_�J�yuS�o��v��𫌰�.�6X�����~���B�hP�)��ݝ)z� Է1��#5\�b��{���y�q���v}�u+\""!ػU���h�V��u{+���V��H��"�@e����ő �u[ս��������|e�#���R�-5�T.N -�e� �E���S��A��8���cy9�e}vU�@'Ρ;Y *�>��N�;��`h���t�����(�4�X������ �&�K�j$�=���i�|���>��:"�QރM��,����m�IO�/C�-�I��8#+9�d�d�Vb�/�ؔOI��+��f�}U�v_�P��Ռ�F�,�JL5H�#̣��C�x3+�ˑ�{�㙌����nT��4<��$G>���ok5����ʹl�S���H��t�?R��O[��R��K�kcᱳ��w�Q9(�ܘ�%�![��8��~Eo)��-�Ec��<d����.]eB#�G=ݻ�����h1����gxB�_�������ׂ���w͸�M�`�B��T��U�x�QG�r�;�2�$/����r�KE�	G�󜑦�y}7�P�}*���h�i<��'&�ʉ�Rn�
G$���=�^����� k�v��i�1�ѭ����5\j'�@m����fC���#y?���Xx�>���v�+�3��5.�g;i�5蔼;����]�ޚ����Ȟ �����k*�(Q�����3t�o[KZǧ�Q�����|�a���`ՌXw��r��}���U��>0{��V���c��B(6���ݣ��c���5�f���S�b�8�Y4T6�x�o�B�T��R������R^G��o����i�j܇ѣ��>H��,��絇M߼��&�6dnI��l���,��"�f�k��cO�h_��)��WK�Q��r��B��:`��zeX��iJ��ELpi��v���^ �8�G��B��b
����r�͊���ќ���z����j
����9�0g�fC��f�aI?@�SH<�I�'ً\$��Ղs2޻��{Ʈ�t�Z+w�~@G�{ �NB��P�x��l�*\�ZY(e��M�D������n_��]̀Lr/��PR
K� u���n�d��_c#P��\^�޵Sa�8q��䷅���s���1���P�cQ�cR��X�eNR=<�P>^P�9 1�D��7e��@�1��5��V:/��? w��|�ۅR�r�>���+�o��=6~E���!����:����$zA���by�z��>�9L�B�j*���}��\�u��$C�c ��9���u��$����p*�r�aF�R�L}��У�_�9�ؕ���'"ݮ2w>�1����;ڵ|�{ҕ^��F�eQ[|F���0�C�Wo�#�K�F�^S�Uj���Nҭ0j�y=��:�����Z��D%�f�ď�
�������j�]�<6���p�$�2[~[�1�5��p�K��Cr����e�P�Í�mr?E�q!�C�\�"��E g�����>�g0����{�@�`q���9o���]�X�G-��E���8#9�zqR4?+Jq�g�ݎ�*�b[[��e�<Ż��TBWnsh>}�ܾ���i�Y/�t.["�py�Ck��q����L�|�	Zd7�����\B�˨C�m$$�Ui�M��
^#o+��)�a�.��9����	�>�!U��\�;�#zA&.�fY=��U�J���Bĝd��7��nq�������9k��j1KL�W;��%�\�2%mJ.g�e!+��k
�2�5X�G��rk�P"ǂƆٮ��O�����b��4L��1����N]{��|�E�^�l��j�Q��T�|�G�СuJE��,y{�ʕ��u3����B:�9\��N�	���%[	��؄,���)~YS�h4M���:�sOC��Oc95ޥ�'m!)�P�\�E�C9JU�5H���h���Y��6���	j�;����!�Ț]0}��性��5ДBx����a�M�Lx��
*���t���R��oYp�?�;�Q�E�p�ֳ��	v;L���dIx$D���1TMy�]������rcf2:%�k���ܟ[bv��掷�'��.Vvj�X���m�61�D�sd{��?rZ߀�����<KD��G��#@,��e��$��S�.s�46D�m����䔽쥼����i,�<ݿ' u�E��S���̺��t�HV9��i��v3��� ��U�S��r�2���dX������6t�c��w.ro����C��M��E�ot�j���5�)�,�/�В��ǠƮ��K*��֊��u[(d��v_��~�a���3o?m壈�[����ċ�:��������K<ez�]ۃdq&^E$��nw�٫��C^�sEh�*o�H�r%�(�~��س����,O�;�5�V����G�`!| LNu��٧A���s�ք�?�����N��A���N���#"%ȅ^"��,-��1"��� ���|3c�kfh�s�y �/��䂤k.����p�l5���2~���H����m� &� �{�JDV�/�K̑X�z�f��#Z�8ׯU8b�ska���2V�X��r �H��6֯Kz����_Zq�x��(�OY�~7J�	�������u�MI�%n���b�c�c4q)�c�ݡ|F�ɕߖ����٢>����V`�?v�=9�Hq�1,3X8��v��KT	]$�}�x��|k��dR̿ �9�~����8J@�#�-m噱�tl��M�1�����+{��.��ֳ��|�"-��7ە5�T���j��Bc�Pn�K�x3lE�Y
 � �־*lB�?�[�6;�:�t�m��~昘bS����k^J�s<��5%h��RclX��q���y;�5�YbTQYe�����_%��1��D�^?���K��R1�2�-��â�P�	F�@�vÌ--� ��kd���3,r�Vܫ��i@����gh*�Z��L��])���L��g�B� ���!`���1�+��c������k��^v���6��Ck�B��C�n*����3{�I(Z�}|s�`����Ko*�r���B�6BnWѬB��f���F����Kľ~u\K���QZ��ipAȠ!Y�
<l?�����LBȼ@���IQ����dѸ����B��� ��l�����疇��Ю�9�n�>����ꩉ��V�_ΡS����u|�r$������ʲ���a7$װ#�F��ur���Q�b�:�D���X3J�����Z4��挔enԕ>��{�*�Xf�TcuެW��Ƙ�3G�Q�"?�N%��O�,�a�O�&xb�4N��MZ<�i��&Bb���h2�+d�C��1��y���ʯ"�'}?�52���<����ż8V��ے墚��5x9aK1�.<���D��C��1�
���6F�ފ�x��{�(!b�I�[0�]^
��V�L��Ç�S��x�AH�m�FF�d�8	�"-6�x\�Iu���6�J��L�0'p�o��8&�Eӫ��
�yI�/���5~�� ^?CyJ8Gu��x�2{e����3�[gVV�u�&�|�:�w7��15GD�]�<��n�x�6���ٰ��S����6�`K����0���e����H���'Tf��a���
i�n�#��p�Q���[���<��ȑ�^\��s0xm�w��p��� �!�I�n�cdA��ָ���a���A�-��a�;a�c���0"��E;�-$�0���[d|��˒�%;�>�Tm�!��e��F_��{��_�*&��r^]�­�����v�G�i����F}&M�PJ�1 ��\�%��B��/^��q��ku͕[x��$LKMP��zx86�,�] x(�Yaub�w�)2��	Ԗ�1mw=�,�9���V��oSd2#��#�ڬ��I-���d`��1�"�ctj�٫"�O!f��?b犥=r~Sj��S�1L�,דAb�!y��E�^M��O��}	JX$�ޅ�If�Mk�5V������WQa�} �9v����y��P�.��N3pq�����x�I������6�?�>�$Y�^D@�ك�HVOo!��t
�������6�tL�f@���7Qq?pYT�B]V�C����}F��C9� #VT}�\H's�g�����}�H�&`�t]\��sX���R_���P�a_U_��đ\ef��*0��cU��a)�Xs�i:�*ɕ���,�r�/���U�ar�0U%ٱK��M��Dfz��$���m;�}Ȼ��H��B�,���P<�9k?g�p����T�$W�x��-w��A�;���t�v��91�[1�}�Z2�4�_4�W��>�_����:J�B�0��v�$t-Ƨ���~`ϛ9I�������Iy2D����ԝR)�b����{F[i�A�RZ�LtXߟ՝y�J����5�y�ό�\�c^y�d"Tn�5*�:oZX-���Q7#Ցy�� ���^�Xh���Mx�x��;,�����5N�@(���Һ@b�*��k����m�4&�6�ͺ�������G���2��2��.�_'r_$��:prgv��Hg֧����\l
�4�I�)��p؃�p:y�8R�Y�DL��l?/t�:�`�<��A5RO�r����2f�W!.ڸ�۫�����R�O����g�&J�z�;n��5��G߳f�jm�,������O��m�C�������{���Z���9G��U��?�Y^����[�^0 �����@?6�����@�S#>�L��zn
O�ߪ�ӄ������ ���jw�좹��׻�Pl�s����F�"љ���{�����Sh�MUz�c��
,�w1����=쬰�(��u�:v�Q�e�=X�X�x�C�.^�R9�v-� �N(�j��|�u�����ű�$�CPEP�V�Hޯ�'1Z=�E9�݌�����1�P�4{{��hS�9�@B��poK��@2�1)��G��f*v(.��~������~b [�����<����IONkù�U��p�༥s�^�'��^S.�>�����X���]�C%��a��� �;��NV��Dd{]f�v���.��/BpOɨ��TD=s��s8���_����iAE���E�*�Kz��+j�OnN��$���OAqJ�|���b�wU�OPH�n>F0�OȂ	s��� ��{^�I0>z�⯝��]��e8�ʷ!Z֝H�Z�p��W���$�z}�S8��'�ͤ��=k�F&�(V��e��z�j9{���g����<qᨱ7��`�<��t��1��/�!G@)��5�:�u�I!��pG�a�E������Oț'47�,j��bY>��S9�v�7�t&��Q����u�M��E�|ۥ=Q�=@�/@aS/��ŏ̧%?5i��!�L�c���i��Mo�Na��5�@��P�9�m�[҆���%#��y�b8^�D�<�������Lʫw��ǎ��_�b��d�[�ݨ+��8�tr�y!JȾY��!Z�t�T���K:��񑯄��44Z+q�������B�Ƿ5��"_��gK��X��{�Մ�w=�,٪WlZ�H�v-��'�>�a� ���(��]��ն9�7�/�N@�k��H�>��e�i*�3�����ߪ"��3��f`�-癁M��Uꨑ܏�U���}�f���X��C�j�݋eo�~RS~<u03�_h[?g���J}���d�u����Щu>�ǉ/`o�D��	=P�����Y�����(�%3��RW	$h�
Kǳ��)z�-�WAR�=ی��'焒M��;^k�֊V�cS�j� ��޲��@,��_ˣ�W���U~q������@&��6���i�h.x�ҋ�|�:�L�J%�~������>��X�_/c	�v�����G8�ʅ�D��z�*����_��BD&����?7���o�ۚ�C2��X��{�xJ�%?C-��q%�
�
�I8s1�����4N���ק��J*��On�(4��1�Sઓ��p�gN��J�i�+_���=/��hC�s�L����
�$�}�z�N$��p@��G�V��=���&Kj�j���CY)(��5�(���R{<tȝ��%��C�NE�e)�P�6t𵊺.�s�W�����J�E<�0X�z�Ќ�(�����s��Յɥ�s�:�|՚�05�5-��?Y�s��1�j��j��cѲ�UC=���\��􆛕/���i�2�I������w9��o�Vs���"&�O�aȊ�f1���G��r�J���������݉H��̂E�@�=~J�j��K��w��VEgZ�Q\&�9J�=���h'�X�tsV�+#��y�p	�XA�G^�9�:$3�^-	^��$ɽrT����F Ox#B�ea
p�r����۸R���)�����04��6')����z�[xjmUY11D�)Uݪ���Yi��}� �?�&�
n;3��eW§d��j�=�Iy̓�x�I�T����ӫ[��Ig��aV�z��G��E����6�-�GZ��+�l+���0P��ؐ@�b��^��;����m�#����Ӎ�ݙe3��Q��"��w?-@�˝�����ʟj�2�Á%x(���
�TŐ��e��3e�u�%���P}K�*�ψ-5�6|�L�'�A��"��@�g�"v�<���Bb77m����t��n�ݔ�����<@[y5	�^BO���S�4�Gf���~�U��[#(hb#p��۸f,gA�.�� ~N%����G�S��D&;���Y1_��bV�d �hh��{���hY6\�Iav���/�^H̜��S�贱�|\iM��/1��~t�����z�,�e"V��7�c�	���F�� �/n?�/��3f��lÛ0�g "���*o^OZ�kmEx�RV�W�V��"Tb�pׅV�"�\�=�.���,L4�w�.9&���]a�l@7A,C�?H���ɛS �j�.T�U�: �.���~��I)�Ɍ���|�k0M�1na��S��O�כ����H�y϶��L���o6�4T�H���G�\:#?���7�Ty?D�T�H��J��|����'phJ�w��P�\b�
�r����ǳ.F��y]�Clr�#s�T2{C���&��H`��w&���kyfX��R�7y����6}�Jٷ9�$�����.tQB�e'��uRF&��̐�7y��$��?�PQ����*�ty4Ekټ�Å.uq=������R}����L�����vG�.\��Hh�����sr}�,ROPz<�]b`��
BJRu$eɌ���`��|푝��+^Y}�Reb"�S��o��Y�t�.6�sQ{O��-ٯ�A�}�B���7��ÿu1�n��~=,p5m+���IW��NZ��6~)�_:Q�Z��v�F	YGU#W�n��bΐr��hjM��l��I�ˤ���|�K����s�{�I��}:B���b^�?���FR��!�SȖ�W;�V��(%+ß�݆���hn5�K����xh�*�1|�y�=1��lI�}�j��J��2���l�t�d�Y��W	�z�3�kP��˝n2�X��n!�t�-(��c Ѓ�s��k�Oz��=��>��[�C��a���?-���q)Q0Bf�R� ���Ҡ��&���'o���ݧ�'��5pf��Ϻ������Bp�����&��tH�'�2�8�G��8��5C��s�"0W.*�w�$�2Q"A��<�.@i¶��e��U�����Ux�7��l��Sk嗬���7�K"�+��}��f�����G�1	��ɱ�l�Z}g��>�T��8�|�_���8�K�[	�|G��K���Op�y~�� yM���ٖ]�"!�*�BMGO���S�My�I�"��Xs��;^�|�t�(@SQu�,F� �,�4�%�Y,�goIC_�;�ê?�Ⱦ]��t�H��İ��dN99��c�T�WRKfh
��&`ƶ�UG+b@�^t b�Hr�	w�o+�j`n���v 6�������%p-_��I|q�g2�b�D2��|�2}�^Pm�#�����;&ʕ5p�5������Z	-���Lے��bK�v�L֗���UQ��;�E,�G��1�x=o��Eч7����L�0�c!ٌvH4#M(�`\B�fU����_�,de�����D�.\޼--��(�����8-ާ�ғ]@�yZ&�=!�7���0��o=��jc�a��o��SH���%&*�P��0�E_�ү��T�vX�䉯cXkԓ--��-�m�jp�ۇ��2��$G����[�j<��q�U��%�/JW��gU���������|�����:�ƶ�
�6��[������������eSl��Z@��3P$����\57��� ��QL�������H<���>sS3s�.a��8'�,��)@��i���F�up��{��n���R�/s�u���xr���L�o�	�v�_�QL|ۜ�	Y:9����d�`)G����YU�W���t#Q�T��)�W����8�Ns�2�*�\�s"�=���#�H� 6*��f���=��_ƃW��J"�n\-�׌���t��ų�NL��� c��T�8T{OI�r���Ԓ��P[�?�\ɋwܶأ ����5'�)7����m�I��i��!
+u"�a}CC����3)�DbJIՎ�j#�޳�:nC�4�:��I�@�C&l"6�f���m~���GĄ[�#|�5d�	vfl
���7�ʑb��`��C!=����ݷi�.!��6)�¸�W-�*�)�3M��&�ՙ����n�Ғ��P�%v�	"�����t�p(�0���@��SP��d�gt���s���>�a��v����i%�hd*�����s%-�J�&-C7hi\�J�˰��VV=��p�5
������Z`^Փ�
 �Tc�E�f,�oV3a��(�A��M��qA���:�J�}f��/����P�}�H����s���.0����n��Y�D��?@���y�%d�*.�D�)�h���<U��i�Ʉ��������LR������Ф��6(�ۘ�L�#� �����Շ*._����2EH�0��v��&Kj��0 ��{[�㹋����%��d3�q��wB\A�8Ը�r��VU8�����yiz'��v�)�tץ��'�8TY�_k6~fY�(M�_G��E3�˰��H�>��'J�^�Iy]�¸Q�	U���x_�"���~�� �f�� =���q��ԻA����R���kޑ�����_D{,2IH�.l�a��BL}��ʹq��#�Oċ`� ��j�pr����WfB&u�e�=�<��	�kA�`o�'sO�Nb���S-��y�����}��EK�[��!�L(��-}*�Q�x��~p�������o�H<��J��Ix4�:���+p��m���}����`�/�D�W[����?��	����jq�H��G�2�<׭	�Ͱ��
F��@��_,���i��:��*���l�j0FBwї���(Ѭ642��a�G�����h�矗 ��m�g~�����c�x��`�!qb�B�O_XR��Lr�t+K,$%(t?{І��T�V7/8꛼�#��d�W]��BϺ �����4 ��p`�k�yg�����u?�O�.�
����|�d8�Á�A��OwY@>VO�}g�q�U���Gw}dx�%2f�GzW�M)�3W���uѪ�]�\د��t�>�c�f_�e�I��4W�s��qz1�A����r��KV�"%�8o?�9u4�f��Ɔ^�?�&R�ˮ���Җl�j����$�:��W���3Lr����J�;���k���~���͐(�ɐ�jh�,���ZPm��)��vE��C�=��bp>�/���P��[��i[R����H�܄����MQ�ypʒ��yØ"jH2�+��YY��r��+S6ı�D�*'���W�-�����(i'4�r)���M����hG��F*@�Ӿi���h��3`�����G�7V����op ��k�N,�TIm��<�+�K��h�=l��^�5M�h|y5��^Ѽ��Cʧߚ��[��^H��1����|`�����Y�Gh��z�-�$��BT)G{p�R��v�kj�h��>�M�d�1�Y��xKJ�$Ht͕=���7�K���>9�� ���j�sz��;&4ث������ʇBt�L'��,��Ȳg��JJ��%hW����� ���]�K��E]��+�=��J�R�����w���(5�3p=QGi[�Xk��V,ǒjJ?HNyM��8��WN�-u�uO�f	�G̈�g_�>T�"�Pϐ<1���l{V� z��s���
�f��;��"�k�P[1�r�o���m�^��eo@«d��p|��n ����$����|q�Sv�Ol��N7)b4qG��s\�����[.\����@aPZپ����o���Li5��P\��
�a����!P}ʇ)�k)�����S�K�n˥�g.�#t^AV���ΥsUƟ���ȥ�a֯�j;���{gh�����)��!�K�0a�7M	����{����^ND?��Qi�5��"·���a�Òw7Ϊ�|R�����Ap�eߦ��I��t��J����<��:YZ���ڔp��!��>Z<�,��@��������eHQ�i�_kk-���;�	��/f(aU���,����g6�!�������}�႔j�p2HQ��v%�|.��*������m�L���ͥ�b����	����ң���ap���0���HjL'����K�%��Ez�,���������8(Q���/Yf�=����(����!���3�]m��*�&2~\ 0�	?�#��<u�"5K0�f�ge*W��t�Nr�4�?I���7s�%Ev��!w�{���[�od@	G�N���#:L����� �����=*�dN�\ L��Ȓ
����t��Hc���ӟa�	�X�#L;e��S�>밼�۶�5�.|%-Oh�
!����):��]��b�0����9t)I4���e�U�̏K��`f� ��qL\%t�/�Q�n���s�����ɉ#�3v[&�}�\��eX�Fj�.?�ӂ]�[W�O8j�O�+uP$K�1�X��\�j�.�j�ڔ�<Ad��RH�)'��m���Q�?߻O�.���֔��B3�x�?\[���v�g�wZwi� 4#��
{�{��W�<*%���Zt�a��2r�S���6�}r%w)�(P�֜(B�G(��狴����|���'�`�z�8@k�B�tB��Ո�M�1�\�M��k��q�a���hF���D��蜆��,�>�n�Tr��p��9��WP�ؕ�9�R�������T-Z���&s8u&'��g$%���;ߛ\�o��*��Sr(�l䵾��$�����e�xvć�l%���dAea�uU��&v��$�ٽ��+�$i��-G�p���D�fl⾄���D�$�Ӈ��~Sj��C�_�樍v��k���ɏ���y�U�� ������ԟ�Xg�g��ľ�~�"ֻ|��/�Ұ'�M��'�q22��E o~8y�0x8��k:x�#����|c���K���[F�U��7��N'm��"��_����6�`g����Z�C�*���4�,Sޥ[[�:|��7��Wx�u��F\��ri�N�(�
�����1o9#��a|!H����wxo!�)���2
D�$���*Q��sI���?F�_5��|(`Y�E��L��&��7KH�u��_hM5�u� ��Ë8�]���Rڝ1��q�LU}�n �	��#�Pvi`U��/��k+�ARl��;l�W��d���'�B�s�� ��Ӛ?E��o��u"8�!ˆ�u������p�چY�/<Mz|�����2��^�u^��"�r:S6Ѵ-��Fei��J7�\�'Ñ�a�9T�N�3�#�VV,��$�㇘��>F�L[��ԝ����s7��&����c�q"Ո�I\?VB���r"T�;���-Ekݹ;2+ʔ#� "�o"���6Iρ���ˊYdtk:���l0�O���,��B���ݩ\���ꦆ8u��^w^��-�m��w�����x�ݑ�|G�`a�����9�b�j=���z��kTg��t���Ip�S��|�����*���/Ĺ͡vl����E�9e��0���ʮk.��b@�$|í�!��\�p������v��&9:4�4�Hl^H���)��e��8j�]��i��5i�`�P�m�X�4�#�D|�rD�W�s��ڿ�5#FJu�o��j�nR%{q�	��hNl�����۵&�z�P�K@��y�m��N����$�,��<�i��E���*|������z���og$�������ѽ.H׎�5�\������z��f*}�ɀvg`���s����[�W�oؿ��>�@Fń�c{ͮ�ǎ7Y5 A�N�R��ʍ��!�D�������G�)��ه�2���9�%Nv"8߀|bWD�����]��>q�̸�笑p���\ڏU��yi��)����O���L�T�PU0�r��j�*�ļ{�X�ᥳ�����3�|�X1=��� t�,M�r×&�� 	��[�oFŊ�
Ƚ����VLJ�b^��vo�q����"o�*h|�gO�z K��������x�W��G�-5�U��g� J�M=c^9
b|��s<�]�I4e�NZV Ҷ�����SR�0j�Q��N�P���C�)7������#;��[:'gU)�C��S��x�se;��ځ��A���b!(�N9��b�|�=򑫻�ݑ���ۃ�<er$�������i|h_�0ӕ�'���CׅY��橯����D �k����� �sj���$�����K��Ȅ�W����0����3�"D*"5�7Mn��X��X�e:n�}Lh8��B���m�8�4hKQH?���e�ά��o:q� �0���i[UT{��
��n�4������Ґ�n���Oz��#;�}���pmT�, 3��wc-���h��Qz`�#��?�̅���ww�N�D��T��U�39]m���Cq`M��`s�LqB�0�r��㪨ү�.V.mx1�q^JZDYZ�x(��,�_bO%j���3ܒ+�\g������S/��V�r_�9 ��2������
Ax�Hmtn��1Â'XQ��х�w;E,����snm�+�
��?���Nl�2���uӴ'o_)�Z�R>	���ՄK/��3hK�w�]�x|�Xzŋb� ���.�|�*��{�u
�ڒ��:�p��D�r�����Q�&j�8�L������\���݂1/[Α0C��h]����������@Q�tA���g[N���lG�f�u���nj��kp��9����u�f2$c���Y������+�8fF\#����K�X6��,�̄u>���vٽj�ԎW��Ēua���T.�Y�������#3)|j�s��1@
;�s���޿<;"ߋ�<�#a�Yh��K���aI� �oz����p��ݼ%.�Q@AÅaQ�,�;/^�|r߆�r���F�zb�-��>����=:�h<^��/���8��R#gOol�Uغ_�C^���9j�߄3ʏk���&�v�P6G��U��jG��F�wC)߇���iЪ�L�1*t>��#�OSNCP�F52m��}^YѳYyeԽ�iO��Y
�9A�����8��qϘ��[k���V�[n�s�%�AjXk�~ ֊!�8:�=�vWyƂn�mC���=�����ypWJ��D80L�m��ؒ1�I�l�:���	xO��=�l}:<�,o�d��Z� 5��QU��}98�[����́dU��c`-kA�-/�Iv�H�7Bח{���"\ୖ�9R��o�J�e} �/���V"��'�˕)�8F�AY���,{�*sqz⮵�9�Np�멷�f;��U���X��ZQ� ǜ�N!� 7�;�NAug!�!��Mi�
�Sf��JR�����Y
���Dp�Y^�bH5\9�X1ӝH����vNF{}�$�I�-}3�4����B;Ϋ§Q���K���s-D�/����  x��t�N�c�'�7T|q���G���9����y��z�ӃD���������dg6�ˮ�-Z��Y��f��u�I�1үۜ�O�L5}��)�q�^��2̱��U�tO!����7��1��;͍��QL7��_O��9��V[׈|�݁���)y7�������S�#xV)]�e��?�c'G?Fڳ���6̶0ZG���]���='�L��B���������]��1�/�`���f���H��:vdu���"ws�0DH�忆\-D���,��t2iF�s����Py!qP��4�'��Di�i�o���%Γ�7s$�<-���^+��F�����
�Y|*�N����;�8I�%<�L;�Ef-���q]�h~!������OX��9�����ZS�SI]ݔ �o��� p�O��W�\p�����+q��"P��s����}%��R����(��ӏ��ȊJ���x��o��a- �q��<����`&P�=85`9\{Q�a�9�:��%��W������*�����3x| e��C�S�H�p�{�����Hq�ґ<�@�9".Xm�OdcUR��Rs���DA�r�E��l9�`�x�|{��ۗ� � ��I���	�א��U�-6�Վ�bc�!p"�hr{�h�=��ָ.�<�z�4���2��|��2�P��9�6r�秵��v7Dw�a�b�RP8���u:���3|�'׎�`F���,�d��A�t�!��Y�m��^����B��r 󣽘�	�j��c���Ѕ�R»���v�@r1I���$'$b�[A�of�W���f���ZSi��Q�V\�����iҿ��5��V�
q�.�����z
i>!&�t	0�����.�n�~X��PՑ����w��x8^s���yPj�>9�ZM*3����^?36�`m���\�u8�f_'q5�������P�%W@��dp�	V}����#��Ud�K��9e�i`��9��^K?�?���Ԭ�M���cg�{s�ArJ�}�'h�$+�XB?Q�7R8�rh��7��̕#�?�Q�Ə˨�K�}�_�*����W�����h"���Q!��jZT qw��f����P~��O�sm���=����>䤮�����95X]5ѧ���y��b�R5�,��˪�;�QO�©E��`�M�`�:��8+v���/�?Tڸ-��?� ��1;�{*�]�'VH���l\�|=
�����@�ϣ�!�M����Ț�v=�=@���Q#����Y��i�Užv����-|1�9��~J#�O|����NU���'�O��	��k���Jތ��:=�[������_�m��GngA�vnK��u�L�a�xy�v�^��+�Qd~7cEߺ(n�Q�{�7����w���qćC�P}��8����˲�/x��W�7VF)0��kӉ�)��1a����;!��!$e\�$�0������z�D�[;��R��� ��P��@�]��sDO.N:�#��xL����q�����R�^��͓�@��{��FW
�n�zP��w��T��� |g�Y>S����~��|�bY`B���-Z�3`W�Q	�}̻�lb����G�V��[��v6��]I��|�>����'Z�t��^�5N"�Q6�ƕn��35CiS�my��PJ)f^�Sw����������^�+���M�N�h_�c�So���@���<�`�u���R8/�Yp�ֹ>�x��`�H맫�56�w�.,*D�㋓�P��K��o�%�!���+Џ��ʮ�u��4���^�)ꆕ%L�������z�:�a�9iQ��T���������2u�_�ɘd	���nL�[�c���Xqt{�����>l�L��	kѤ�p:�BT���$���T1 {	�C�S7�Q�=+k7�ڱ��#^����D���	������VpN���H�pM�K��~����9�A�/�*�+3��l(�3^;����x͝M��V]��4W2X�r�I�7,�[�L�ښ8A>V���C6P���!���~$2�z�
th��3� �\�/�Z��"D�{>�cj�y��ʎ�b>o�������n�G	�wy{���{@�Ӷ�~b�5����gg�?����ra?�E�'ح.�I"W{�3�lǉ/��?eH�2�=";��R��W`�ɰ��s�p�V˳\�-�GE�6�!Jj�z��>3�B~��'&����Ƒ|/�ġ^(�>�ˍ�"�Ǣb�(W�0T]˓�l���i�
�-���3��1�g)��k��*��&����я{�E�}g4\��i�W����
�%�J�ڔBm���~��vL7��=	�y�":�7�w�T8	~Kz�.�w��/ql�;�v`fU��#���b�ʤp��P��a�����5�� �o�]8t��O썙&��7���Ŋ�����vt��z��'���c�pT����e2}��o�i~M�b+��*�{�>X[f(�Ht�_�pU�h�g�d鍍�M��
�q�z�w��uEsl0!&��t���j�{�:^]|�j�9�MrqD�~��i��6չ'C�2�"��T��>M��i�#N=���&��������ߵ���c6*D]�B�*�6�����Q�k
9_;`�g�JM������)0{S�Nݲ�&S����_��!��V��խJ�����f�ULnV5����s˥ �I�N�!9:������(�����?Z��[S��o�8��e��Z��9 Tj*�����H��r��5��ND�rR���ĳ���r��2��[Q�bԏ]C��(Y�s�ʚ�dbMI3����2�8����Kv��W��/�kg�%��>J $P��
i[	3�=�Uep�6�؂z��@�"�E�k� B� #����&3\&�`-4��U��U��S	(��ș`^Yu�<�7�����=����@��Kw]U�0!�f��@CWGA�YN��k��T*(����P�����,����&��&\��ה}U��Īz�t��/
�X �̻գOF:������;�7/�:�>�>�uO+�o�鬾m0�c�m�u��џ��?��h�NR�I���M`7���_�*Sk�i]�bk�`@��J�ۑ�`|Դ��9D}a�����r$��G�^D���Z�OP�i�hK�
��>�&Y�18c�"�B�`n�)k�{���ݹ��x�{��@��ԅ��}�=�u9�Q���%U)�p��<oG�nN�v�2 
�1�a��f�"!��^�=.�;�����`m��2?]�(��䁔D�.�g����N�3"[:��6�+�r) 8�ף�ה�Ȋ�f���=�2�(v����j�k�in�v2Q�U�zϿ�~��/��b�^�L������j�w��+埓��)����¡�"#R�,��P9A�ϯC *��&���@`�L��M���79�!ϫd�8d��l%��o�xJ;��1h}��]?��(@3>��al<��L!Ƃ�"K���SsAo�h�+]����Ox�`L�'�-���CcF��t�Do� ���!�j�_��r��R�b5e�'~VԼs��h�{{�[;UZPY x�p��P����7�|�G���M�q��}�>�ղ<�}�a\:y!�kG���Qm�E
1��و笏��w���C���
v0&�zwp�2V�����q��J}+$�5��r)���y�a�g\L�k��T�����ֵ=o�/`�U,��ޤ��G�S����pJ��X��&`X�S����D���`NJ�9��[�n����!n8���^������Ŭ	�2P���#tz����@t��֘N>�K�͍��C;. b�r��6'�/wB�in@T	�2����z���?�����H������WE;�B��Ttf�k判�s��W�Y���m�T�d)�	e��mG�w�)��L��)�^���C�t!��,�f�����X����@�ŧJ�|#볙�)�(�\��x��a�R�W2mj2 36pr��|���H͈U�W9��q��d���l?b +!¤N�3������4\EG�u��� l&��%��\fm���Y�~<�ZF��+��ڭ�k��&��n�e#>����ҤM1� �pN�ęxR��(K�{�DMv3k�(�ƕ6�k>|�jKӮq��!�*�R�/R�UA�EW'�n3k�V���;j�zx/Ln��^n9������5A��xb,p0��c	=���AzP�	���dc��~ڬ�F�"I�L<�T�ӏ�&�����7n8�)����omM_8���:�.�HanAI?�Д����`�Sy
�8�>�'��X��e@�镛��NS�~�{}�aߦ��mq�p��Fe���V�\����Tv��
��L���U�j�r/]��Ī':nX][Ĵ_���
|E=ɼ���5mn[vЀ�8Χ9YR�j�V-O��A5fӢ�l�` �X/�� �M��V�>"ph�����*�Y�@s�}K<���ؗ�_��K��e]Wp���.�ݰ�> r+8���Ng���^�� ��22û����%�9�I�r[�tkk"w�+�g}��끯M�t[B�B֞���-�F7��m���j~�#��=�*����E�T�<����"��4&�����x���v���o!_�4��@R�@̣��]�=���t��kj�p�\r�
��+NմP����<Y��S��%@�` D"�v���]���6ͺǲ�;$�4�uNK-˭i�̱���I�|SQ�I�k-(�h��R)9ۊ���	nO!�4� ���f|�r�yQ��\:�p��
Vdʸ'<��sZ���u�`0)��<�9 ��v_T�Ngw�Z��|<�'���l�S���8����ȎV=Rh Ԟ����w_u���d�@���v-���Æ�V���ivܲi��O�����x0@m���+�B����_�D"X`�J'�TT7�
tWV0�m`�[�4	�
�,Z ���[�K�t��?�s	��UZ$�L��@�sG;��b����lb�	&XT��o]�t�����@�R���#w�c)�-�@�e[��wb�6c�!�`����6���ܠ�Em��ĆY�WZ������	��X�#������h�W�G{��qosi��rwAVҞ�ZE�#�m��|O[�����y
WI�*��0���_!@�S���37j�����-�>z�>IZ�j?烘��y&ߧN����^z��>�S+Ԫs�A뙉_��S�u4dq��#-ʞ3�o�}>K�:=��?l���0T*Bv�۫1�MK�) ��,v�H���:�a�a.�Zo0'�riP��]�E���BG��HQf��S�?:�\ܱ&76�CU�]�d�$������kx�Ta(j,n�x��[�«��q��"�a\&ʝ4�x��(�9��� �e�*dk��]b�w�U��g2i���+��e�㙢	�##h���o���NU!��\I�;�@���F��l�w���독Ev��0��mI�k5�C�"���R'��潵�����h��r_IX0ѭ@��#ܓ8��$������nɊ�tF^7=�%����;�.�-u`�@����j5�v_���z�*4��D��*jRnʓ�j�G�Cץm��A��r	���8�sh��'��Rݘ�<�m�A=f�g@��'�{�Ա�� bt��f��v�+�a��B�l��^��bb2���ⶈ��M�,*ſ��������Ƃ�=��/�B�%O�ae�=ifjpE\K]7(w��/�b�92�7$��m���6�ԝ؄��^�
[�D`=ЀX/9���4�-����ɤ�����/�Ԥf��F2U�� -]d�y�Q(�m������l�-A�b?�I����:ly1��o�gWX��Ē�_�o'x(�^�D���FX�˨y��.�|�aӆ�\�\)�Uc��Rȁ;36ѦCo�o�gVX�;"&Da��� ���Vy�Ε���&��R�'�4S��h�>�Z7�D��3u�,bHq�9���i�	����b��V��V�l�4M��MH�qُ~sQ�/A�5 �U�\	A�����蔤i:Y�-�R��n�B���bZ֫�
\����T\�<C��Y^N�SQ���%�8G��$�d=���l$�u+ZwŖ��y�����`�T��]�(/��}g��(�Fɷa�f�o+�t�6�u$�����+�-���O!K�zc�k@c����8C��$S���Ҵ�vCT,�9�?��:��bQk�q=�u�c����M"����{��]�y�>�pu� ̧.�����zܚ�i�' G&�����L˲��|��<�GX��q�"<Cb����C�C�HhXϥ�*��f"^-N�l���pgҲ�߼ou��9�Q��[�y����t0z_f��>ӑ0�x�䗶��@S����ǘ]!4uO}#�u���J��_��H�G�-jդKhu�v�,�����גH�a)nFox��ĩ,��Q�8��cEVN��_��;�(��=���]�O�T����n���\!�z�ՀC*t4����AH�-��a�*U�^@����O���o�n�E�������]�!��&�_C�:_����d�.:<.Aq��qOm<��N(�E�ガYBo�:����ҵ~� ��ʠ"�\_�&�;����w%m�\5�� ��8��^�>1έ����9����� ���O�7	��9Y��i���q�[��p&��������}v�Ȋ��="��v��<�d�p9a�<�G��@
�����XU�4JǍ�bG���i��*j�{Qf�k-U���"|+�4:�;-���,AL��I�a����U;��iL��r��<5�p��~�5�H6���5�G�� �������h�:�0Ǡ
�� [�U2��M0����,>w�� �Yq����|���l���זR;f��b�CZ��l�7�N6���b�5'(�;��L{X�ϑ/��3 ��:�N�m:��sG�}l|���7YfB��d��ka+��0s���Cc��$ɣ�0S���
��3=S9�'p�	\������"� �
ع�!]D�����C<W~��F�+E��$��LK<{�6��G���-�zK�k�9	��Ջ/LW�F�L�=A
%|ntl2�W��_�Aչ	�>I�q�B��!�u���l�H��K?�f���=�I4�
�Do�D~<�&�nE�'��H9k]d���ve|vߌ�W����$N����q�R�b��(L!˨�ĊXM�W}�����eA�s,Ă#��_3Y���K�,Q�3��2 �)��Z����% �?�����-���:evT��d8�z��/�s�\�y�]�0�D78Tr��XO��zn�~�jw�Xwi�px����S����!����O��C l%���iͥk��ܰ~�ל��un:'�h�@���ݓ�;�n��yIm����"c�FL���t{�xˠ;��\K�Ed]Z��B%�ZL Ϝ�n*��G�ԍ8��}:z�o��`[Tf�%I�+R�N��SC��@�j�n�%U�8�����o�g	*eȑv �(rA> w�N�^�\r����H��*,_�t��z�W�6Ɂ�I���g`C|�- �KvK8N��`	Nzl���RTJ��G\��Πpgg/���Z�d���`
	�
�Q�k>���͇3BĎ�߹ү�"J2�?P�_N"JԣVF�/r�칤�9��h_KTT�N�Ң>u�9��Ʒ0Yv9���ga�l}���em�KvǞy� �����
��t~���y�W��1��8T�f* Gː㛫$u�j���c��ˇ�02|\>��8�D�5�2�m'Tz�Y]H-���Tۋ��_�,@N}��p�]0�+;C�Q����yL��Y�+8|y��[e�UɌUBk��/���[g�JIi}���'!�I0�˄y��)� `RG���܍�F�pZ�U��sO���ʹd�8�4c��+^/ۼ�t���&�����'4n�t�߰�+��ځ��sL��t!F����LF��g?����7w���(�}k:�pb���L:	K�@�{�k�5o�nTP���ĦYr].�A/,U��S3�je�_k��u*��44'*��TV�s�;�������Y���LA5}CG��Q�39$}�P`��<Z��^%��a�ky�ՏE6�����[3�7�����_���jU2x���Pn���Қ��l�~��s��t��Q"��X��R��ՎJX�XY��u&��Z׼Ǥ~W��=��ȎT6X�̤�p&R3��T��F�B
o0梜2kP6�b��8B{�����8�S�� �q��sl���d��)Ǿ.�	m{��h\�c�R�cwxS��s�^o&c�O>�(U����K ����?�]>	=`�+a���H>j�q��R��Eg�Z,�A�NEkH-4�f�^��r~5����\33�P�����X�79? 9��{C�?�m���w��[E&_ ە�e�:��ㄇ*677��% ��Dnbc�����m��C��n�tԑ2� ���߲�i�(8vC 6�Z3���TcLK�PT�G���䋩b��a�	���h�@6=��m���C�Q���a%�M��w��hQS��A�l��y��t�E��D�֠�m�>˳�h�?�D3VO�O�X�8���L�j �9t�,����Đ�W�����O7i��^�+
 p�@���JJ�<��@u���|V�e�c�Q�@�s�Ѹ�I�4W����3��H�_�^+�M&�Z�_�]� \���+`��d�=�v���,�u��>���_���{)��&���K�Ѝ�j�CU�G��?�1ð޴�P]|[����Gx���>T`���N�G��Y���o�t�PU,�x�*ň��Rn�	\���� u��Yr�(_,2K~��$�U�w��x{F0�7�,唥��s�<)�L��52ۏ�vr�c���.��I�;P�c>)��<�Ć�9M������,]���ؓ�^�cNAd=��j����7l�ܕ�Kz�?hr{�j�D��Wo��}�=PȨ�ϴ��8���-���iw��5*�b+z�|<��-���{��l[��� �I��-k�V�M'ٍH������8����9�������m��6��!��,���98�a��9�ҫ��(X��OX�.�v��ӝ��Xov�J��� d>�����"s;�2�6I r0��������m�@j㙵���#�שd��o��]R�ьM�B���YN�^�ʕD����O����Ӈ��C���cT'�aL8��W2��*kz��q�.<E�y���Q�I��/M���}�{��SV���m�Y��4X��2BZ�z*��fnC�8�sRה��	�<�~�]Ѕxfs/�ٷ�ަ�z%X�H�h�ti�ĭ��`$�T��|������h�X6V��%}o40�n8U������4G���xF����8Y�?�R[����|��P6VQ�׀g�f5a���*[W�Z
#�p�Ξ��Q� (�;�ށ\,�u�i��Z�T:Y�]�2);�������SZ����X��Lѩ��f���e���� V�]�]`�oGݞ3���\��sg[أ�Ɇ��Y!�P���9�)7�r�%I����n�j��P�
��{S���E�6I���� �H~���%i��l�sC���6�;W$��M�I���he�i��H����<��l��y�h�G��C�xa�AH_tpTc��B��Uі*e�W򊊳��U������C�ϐژe˭��9����&Qƿ�|�7�ac�Ӊ�.� ���a�krf�^��,�
#��/��G����G�e<��G7�4<}�Ī�6V�Ԟ���bzFUABgKdur�~�I���3�\�����ڂޝ8fm�����}���|)�`����>��2j����r���Ŀ��n�,#I��:yt;2�����*�p���n(��UG�X>������Wb�㝪K�)�C�D��ۛ�����Zr&?�o_�'�Ay��oe�[�#x�Az�<u](@�8�N��m�l��S��tG߲G��	�k� �g��(9�	��!AdWj4�נ��Â>�Z)��c����(p�MELg�pY\��o ������t�X|\���]A��L��A-��E�Ei�p�J�]�d7���m��@Žk?9(l�eF����l|�:#08���Bn�&Dy�Y������7��\�XhI�-���<<�.N7���z��C`$��{�F���CD��V�X׿ddɂ�ns͛%��|r�iwe8u:Ai��m��{+��I�;��1{����2��*d2��1{4=��.U���1	U��Y5{��3�{v������ݟ��G��S���q\�����[���^R*#�0%?&���
&�
�O(�,e�4���Z%��x��Qw"�;��-�g��a@�u�z����#�|^7-6,����¯w.��0��*�Z�� ����͵�0��>����xA�c�g$�ZY��T/��L65���I��.*�͝��v�*��"�@n�{j[4h	v��
l��.7RsW
�r.P.}��GҠ����� K≤���Oy!��UDaU�A��O�Z�80�#�mO���Җ7'�JQ���M)�͸�IU���Q;X+Ѫc�ֿZ����GYz�^!��GԨ�[7��E�X[d�jcn�b��-t0oFan�u��h]�cP�x���qa�N�YTٸt��iF��[N�s�4�F�hѯ����C݊7	b�9�ʥاr�~	����֝ȗ'贼�T4,k`���E��q09D�I>�T��!���zCWM�q�j3=P"��3.��|r(���C�����4�����wz����X$��2�bףP�]�쾫���s���L��vj���3{�V0u��"`E&\�;����ҭO��&LY;�w<�(��0)�%K�xs�]��uN�2]&j��q:.iH�W�K�Z%�X���Y��V01�=$|A��ݽ���T�`x��4��|���[_ڑ�ö��M���㯁i�"��rgP����.�!�d���]<�<FkbZڐ�d y�֏����G�����y����g���Gg���B;yf�h�)��1�gxN�ޡ&S9K�|o�W_����˭��$�(���Ϗ���01���$qt�R�NY]r�Mv���8��.!kK� ��b����E1���wB/�~���Y�:*�e��f�]�����m��|lX;�����2���Txta��MEw�R�H�}6�/L:�L� ��ݪ�?�"_u�� ��^5h��'(�Jnz̤zalr��!Y��))�d��]h����S'x�
��,��E=��wO����˨@������6�X����R �e.�wU�i����6�����(��VFO?VVlΰG�*��㑁f����y��l .e��s8����|��_?�����^��O�({Y�֭w^;����Χ0c��,������ט AEw�8��Z�*����_�ym�ʄ�Gj�Rn�����х��hz�W{��ā�3�˦ƵF|ZZ�"�� "�*�#�F��<TI%[�S}�sb&(1��Pȡ�4��O�2���X����Z���R3��q33=����m'#V��nHq���{���/N\I$Ti��Kj3��T��$ �L�<S;�Q�i����?��Ǳ��?���5'��f��u�R̈e�GN��SSO�Ksz�����lB�Vb�k�d<�=��N���&ߕ�IH�S��|�V";��k$�+v1Ì���bm��ڏ�c����Zv��aɤ�mC
�J�J��J4H� �J ��r�b������׭7EΓ��^��L�j0]��C�kwo�ߑ�=J��!5f}	��J�0#���p����{'�X�d���4��KS��pg��ڷR8��X"#�X�3lR�SyG<��C��`�KϚ�A��ՑIt���g�&�6�t� �d�v&��~u�",��3BnR�1�3���<z�l��}�G�%ڥݯK6��t��4ڑ oRwx�C8E�N:b�~_�Of�`Mt-2����C����,}��N(
����2$O"�{d���ȬUqwЭ�߅&�_�!��KW��S�~�<�e����aWҶzt
ԃ�N.��C��H�e�u�/xG�5��tr�\���aKn~B2J��\�̑g�2�o� �h�^Y&cD,��&F2���ڻ)�=�{�t�+�<�R�j��r���8l�+�ЃUy�f�T���r��AIEJV~�7H���c��e]0O�r�������������ofLw��B���"�eRq�z#f�?0OॹB���>
+��~,��V8{I��P5̩�g�p�~�1�J}��OT�!���	EH}-/�\{�`�����ߕ-�g�&}�J0Iyt�J�J�c�'�w��v[�2(��N1Ʀk~�lDd����^�?��?e�Q�Y���֔���\�u�|Yb�ot���XIm\�E�����W3t�y�yHh�����9VF��^F�.95�к^?�'�1�e+�-�m(l�u|�x��3�(�ɛ��]Px�c���4S�Q���n�A�q��A�>?�x�7v�������xs�W�wP���g���L"��_°Š� �4�{��q�YQ�.��J/�#���a�d���b��	{M�^ {,'���@~jc4�^9���0�@�\7�[m��"�Тf ��w�pu��"���ȝbd�`V���
���*�L��qx�V6+BF{£�l'`]u�Ix�%F1����J��.(��/:���3���֐ђ�D�3�6^�������#�\�HW<�J�ܪ�/T�"�F2����7r��m�� ��2)��d�IJ4c|����I�(iUQ_H�����|e����_/��v`�Y��N`�4̫i)��ؿ\�k��c�r�hN�0��C����q!`��bL0�<�tl���g	�,P���3���ZJ��4N=��l-��c�\�F���ex���O(�*&i���aݐ��lԑ�U�>��5t6��e^���+��N�9!َ��(�OhHDJF4�zb1D>�x�q�@
���n+�]}�g��gQ��g���v�q�i0�Q��ᩩ����r��(=���㣏z�������hZ�*��hxZA�N�5"�SNDd-ja���=��T��wl��C�Zwu�x��!*ptH�in���4�ᒩ��\�*�o#�?k� ����ӓi��WՌ���_Tj��&���K̭�E3 8�͢~`J�l\7e�Z�ZB�K죭� 1��U:"��L�)��m;���/ ��@ozF�6�G�R!q�R�2��U*�&嗽��R����T��M2&��D���Aٖl;T���Wpy��"~QM�k�t��F\Y�:#;M��4#���@��D�$U;
a�h�*nr�)��^�}�;΋B����9لɒ!k�Q�,0������>kH������
��2Z;�K�ي������֒��;&��3cр�Ŗ|#�#>��� � j���! ,�A��42�X�U��ɔ =)�[Ɣ�����5S#k77æЁ$���"�`CZ��<�E�g}�������n�o
���Y|�:|��x�i=;�P�K�8?���.��8'	�{܏�3xE�v	!���LBvry�����_L`�(w��;�D��`�E�l�f�?	�c��2�^fy�|���}���K�O�/�����tQ�iI��&�C��2�>�<��DMT�E�ο�zOO,4����<��I!��-eH��x�H���r�����ǝ #G��ڊJo�ib\o�̐?����F�a''
|Z�u��r��e�xˋ� Ŷ+��쿦�-e���TU4�q\�8	��{�0zS����[� �Ρ���rUJ��5v��^@㥤~3�`=���q)2�����~y�g"V��z٪��*W���o�K�Ex��n0�g{N�����ih�h��2� ��[}���<U^R<>äT���Yy�=ob�o�|n�(���͕rj�E�+�nW�+Qp#qu�Q�0`����%�������mx��eВ�g�Ƭ7�;g+lߚ�V/��v���@��@I��{q��OV1*��x"l{��{[P���4")j?+{�b`���$���#�WU�>�H�|}���ggj��������㔉BƵu�j��M]k><AW���{��fm�8�?Ve��Fl����ڬ)��d�0��Ϥx��G��ȥ��7��j)94]�gOc3W��*�XC�v��_>�~ag���V�o�0ey����R�~������ R��� ۀ�d���%��A7׀���0�3� ����QZ�0�Ag�vu�4�?�O"k=`��b�nِǎ�&r=w�̠J��l�ؼy�=J(�=��#_'\(J�N�0&Jz<iR�I��UN�U����!���շ�~�2I[[�Mߒ yT�W�;~��A�9'����%���8|�6����ێ��C�-G>i���r�X���q<�Cb����3�??`E�ڽhZݶ��p���Wp#0+�x�lM�o��7��<���/:�xJ�x�����Zz2Ͳ��m�ݣC�+)�ׇ9+�`���Ee{"*��"��D���c�õ����$�gW��7[l��a+�h�S�S	/g,<e�E0�6츟��P#�x>M����
�ޚ�'���)��%�p��qɱ�jB� �Z���PT�g��3�w����d �ŉ�GM:��eH\�h,B�C�V��|�R\�%,_��TM7�8����`�ԕ1�]���o؂R��ҡ+����-�툁�-�����*~�^L<��p��g�|$m/����EF���M^�V(��&o��l�ĵx����e,Ȍ*���U�J��3J�>6w��f�:��Fx�Ǹ07\���1�n���c19��0�D����T'���X�v�B�0�3�R4L�|�7���~*>�*XN��ԣ�\�h� ���|�*b�٤|���|���@�*�Ɛ肵*�wl���߿��ϻwgN�C�}`�\A�!���F�5{-yO
�	gP66
GI4�z���W����$-j;2�����y��JQ!��}���!X���!�ǀ�%D�q�'w
�3�	Ռa����}v&�]��]�\��b Ϻg��7��*ebv��8�01�!vRy�D��یذ��,�D��g#��E� ߑB��mʲ�ӄ'o1�y5ȞřJ��^�i�����b �@��*��1�H�}p���t���|TPL�QR���������ڶo몓__�4���9&?~�2���.�+<��k�7L4}ɵ�d�k�Zi�(��<*HM���͗$+V�}������ά %��������f��X�&�\7t��.ʇ��9��C�b���`n�3��C4�$�9�~ �ג����^{�R �r����ݣ��M���<C9$�g�s��k:y ��|����6)ũ���;+�o╰*3�w"l
�$�E�h�끝ƌ�.��5��7��/��*X����0�V�Q��M�n���4�S��
$� O�|��P�i�b�m��*9-B�9d$�چ�������r���bH(+��`�k�?٤�m:��).>��Ͻ -�@��j-2�g�49����LUl�A�Ёy�U�<z����8m]��]�Q0�2O��G7p�dfd���混0+QFgUc�<���I;�J� ���Ohc��JD��x�	8u�������߅�E�Gd���_��c��ԣ��'�Q�p1�8p!���(`���l��U-r9ӆQ��ʲĲ��B���/(��8�%��7Ǻ��ɱd�"��ҜƱp�>	)������X/d��bNH�h,�Oz�P3a��Ek�Z3���;YUm����4F��~~��y0�B��(3��f�9c�c���T���C���jGl����~;p�ihI��5��1�����b"N�& M'�O���/���O7���I���N���D���ij��S��N}N��s��� �dVH._(}ܫ^Bg�s�3���>���Y�5�YȢ��)ż�a 7&��a�~pr���[qx��[vA�
�s��0���k��g`�
@Ih�S�"e�� 3��|�S�]�ۼ�� ����� � c}�m�YB�@�]�ҍd��G`l��t>Z$5�9�+�W;��������;! �i9��㭙�Ґ������wΛw��{��wJ�u׭:��'	BѩT9f��Ű�Cx;G�.���kĸ�"�Zp��x6��G�Zi���MP٣���ވ�]�rYW��x���(��,���?��MA������µs%ֆ�G@FZ��ô��o���&��˕�L"�N�e��ŭ��]���e	��6~��NFeT�!�a(��O�b��0�P%��LS����<�*�Iۃ�l2��<@%��r,�`��M�7�H���W��V��F|�F��D�-T�԰_|J!Ʋ@ȹ�x��y�7��Y�pk����~��𾯍eÔ�Jܬ<�Լ�G���)i�_�����&d(>�~�3���]�P�|;�y3���⾱��п���m>� ֹ5���h�������G�6\��*Gx�BBRpǶ�6uѦVR�̅���g����:51{�.ˬ��g|�5����H�;����Ά6�����%�Q�k�\�	��g�>$�
&vdTR#]�hmѩ�\ȹ� i3`	_"A��Mr�����o,A�(lPBŊ�s8$R��fL�V��OeH�G:�/ίa,&]���ݡ<�fֶ��[��?E�<`����ɖ>�C��qq%�"9o���K`e&����gTO�V)~਋,�
P���Z��ُ�kc��
�?bO�?,?�2K���/���g$�ޢ�t_�"�1�w�SqR\@`W�L�
�z�e���u��鷿��[ԙ�����2Ņ�A�y��hl��d V��|�T�!�kuJ9��J��A�ܹ6َ�Y]�F�R��]�:{��/�	��2�Y#��-}6���������@*���f�O:�єC�x�fw��La�e�TV���Za��%f������Z����^S-�>�S����DW����z�T�&�ѳGb>��~�_���z)������e��[�F"�Y$J�o�@Z�1�|����b���3û�@�������O�r#ƪ\T���W����}}��C~�f���q�;N❋�Z=r`0`!��_��Vʬ�φ�����i����f�ʗ*׬�PT������i��Y���ѝ��G����m�z��i�v�m��0^v4/gU
� 탵
�� ��lvko������ޮ�7��Sl�%�J��<�q6�sC�r\�A?�܂��,�Hb>c {:��&\���S�؜[4�!VǓ`ɐ�h8�z`�Ι.�,��y	pR�;|��bg���O<>�#��j7����4 ���[���?9|��7���ֺ¨
�)sr�����dŦ-M����~��Fr�����m��
����N3$NQD�85X����
(H	���=�l�,�����~toe�����G$rR ���[�fo�����=�p�(��?��&��K��ɧ����E��7dѻ�o��]�h�N�ևܿeh�B\����I@r��_DQ�#���Ѹ�9��b�sI�/z��*Xeߧm���%e���ă����5�r+h���L�L�8���gb)(��V�k��[�{ E#��CK`��`�&�S��uhr̤��>`]�V� Yi>�x�F�\e�]���%��,�Qʝ�����yD7#��4��[��|)s��tSDI�gX�y���b�;�f!�@v>�oEC��������ӓ�V�좚�t܉�+<<H���bN�F)ӼTi��wZ|��o<��b�d2��>��ТTQ�5!:#�dxT�I@�t��ͬ^���}�qp�nX�ep���=��
ٳ$�`_3&ek�1�j��y���3&R��FV���q3<�P�]���n��M<�a4E��[�VG���k��KX���vj���V��~bJ<Poc`n�g�#
s~LwL��:|�}Q�� �@��l��g (<��)�=�&3z��X~.�Ĝ��+�탌��TBBg���X�Ss�2�Ib��S	�-�5��l�ڙ�X���s5	V~�muv��>C����pEYM��PL�`>۬N�E��A�_ �' 
EY�M�e|�s,��GJH��~��=��� wi 6�S�����|��$���Ctl5�)�>��h'ϗZy$h.��k����@��vF�f��v�',�OMB�%�@qK��s%��l��� ��)�$.m�L�%!�i�@��*�<�!�SJu� �>��&�02r�1(�2���ja�����z	�7x{��]�����9�:����`Q��jx5}�Qv�S@�,���������bŻ�a�F���SX��1A]�s���t;Hm1tX�]�6B4�.2�@z��#�ѐ����	 ,!L�\I�t����R�\R�ք�#Q[A6_����j�,E'ۣ�OI�qD~�u�֚�:=i\��Zt��ld�t5f��y����Kܢ�Ł��'4�Aoj�D���Af�Nӫ���@P#�n�d���	%��f�*V;��,k^=/����kЪ�Wa'�m�����G��2a��'����N]�����+��gz��>���������ݲb�\�t#.p�2��K<�=�LX/$3�F�at"N2�� 
����'t�����rv����!i%U{2?*kQK��$�ȵ�_1Lދ618P�J�������L�Պ�~B�i���f����غ2h�j�ghϬ���0U�p����<ZV�"q�|���#ѡ|�Q����d�3Ff��4�q���M�zQ���?t "�s�C2%xN��#�Ѿ+��k@L4vM�B��}��:�`E��X�MWf�^ą=-k���e�LY����?G%�S��C��Dn䡂4��d�pxb��=ș�vh���'L�/�R�3��o����ȣ���2��B��:TD��To��mРmn�yG�P�X�\���Z���nR�'Y؂y`Xh.����}��c'���ܮԃM��D��\%9n=""2��qo�)��ޜ��zS��p�2�B��cy����C:a��A�σ�bC��3����`K��S�����-5��������9��A��D��q�-^��t|���Q�������
����@�/��:�#��P%2�oӢ�%�S9Aآ�f�!�c'�:rx4�4�����Jgu�e(cڥ=��N֭��Uz���ը���@I��v�����3� �U�9w\�D���e��.�kK&�Ph�"my���v!������J�`C �p�ar�]J*�If(�;y��)��|�䖔�/�Ŧg�h��2��>���Q��s��pg�m��1��P��6���� ~�tL��� �>��˸�KW7��s}��5��N�0�hj�H>�x%�p�����>u� ��h�R�fSD�>[��� Ȁ���������[��8L*�s�08����t(����������<�����$ժ�`Is��6m���S���%�#s�q����DQ��r�l?}Ty�����{�B�d��4��p��ł~�jO}��My�K��*Q8|{ult�
�؀�։gyÊc|Lt��c��V\*�+t���)�apB��
Kç ��Ÿ�܍��dq��_��#Z}V����ɀ��3fe���5t!��,�,7+
��P -��5�yW��� %�XQ"б�07�,(���]1�K-vbc��`�V���{�)���J�'�S���/�:P�-�����:×�	A�U3L��*�,�3�Wg���EC	rZ��c��0�4���U}�<�5�F{��.b%hw_zQbU�u��?F��,n�&�q\��P;�I!a	�Lm\���%�|���� '��yRq���qL���e����5I�}3_�U�ꢢS�� ���H��p ��C��W���ۘ�H��"�{��-�<Fb��ؤG�m��.o�zY����lL�f�Ք3Ft��V2Y��� =���\�J׾�#ƻ�>������ Pz�>�ˣ�^�l�zS�~G�+d�0J���늖婹o��F�L��qT�G�yw�!p$���f�ha���PB��#Ȟ�W@����Ut�\#��2��A�ꣾt� �զ|,bIho��������|�v�Y�(/�����q�		���	7Kg�m
<f�TZif�֘��؎)`Y�E;_�c������Z-��3�Wou�&g�ݑ���Y!�������_I��5l�M[��̭�L���@E?�L~��N�2�_�4�im�R@<>/���l�n�]+�
XN;�qV����[�_Q��n��>�RT^F��`����l������>&{��Z`��N�������hF5Y�?�0�(tT�Tz�Ƈ��d�b3/�ۿ�s�M{-�B:�D(NB�;���;S�C�e���p0��_J��G2�����������Ծ&�_�jі(�Nb�l���G� �,s������P_%�E�ҺZ�Z�n���$�2������+����h��͙l��S�;5[CO��ӌbJ���h�5��i�e�Ns�����E8�3|=��Z��J���99�����?�%�k�����'�)�m���y�E�˫�n�����V�Q�+��x�[kv��;#�pq����3��=L�/��9*JA�MJ����n�^�7�* P�/{����{[��A�|�uZ�U|d���$��� �CH�v�)��ޓ�ꐭ�epi�Ή|	�w�vk?�/A!@�M�]f!-h���$�.vX�ꀚ�0��nD��:�l����gT ����j��:�>���b��}b���WI�L�vl#���?��R&�!�+]�.�H��˲���<P3Q'���9�N'�&�L��#.0�����۝�C�<�<�*����i�"�KBB�X|��{�j���P�t�J|`����ӹ�R2�,��z ���G�H�f�(_�D�$����ad��E~�t.i۪��h1�o����G��*ChO-�3WG!�/Y��v�C��m�]��e%ޤ[�/
�������)�i�VQ`cu�S��_ݮT�\_Gj碌���k�Lҗfk�	B�t��DI�,��HQ^�Ľ��e &k�{Ȋ_G}���ې���=&E�J��1�i@�)u�U_�݀��&I�j��t|�@��щ��YC�:�C��D�L��y�R���,�v
1z�ʁ PdF��:�tX�u�)�����Xg�DFB��QwS,�}4�S�1�I�:y�PNތ���%��ԘRz'�#G&�L�����EA�-�`�0!��Ta(xT�����>.���)}�|�f�V�ĞG�A�i�So�[0�V�cI|�7.4X
�~��E[i+�'�a?9��EִP�Ήyz]��@� �����\BDo�:�q�9� sRӖF��� ��פ��� E`�0V �E��웏��JR������g�~=��[�jz�w��J�T6|��o�iO ��A"�NGﴳ# ����iu��/̲��	ϟ���þDAV:���[N�:\$�U�N0˒׳��/���v�K�f\�<@Ң��6��D�b�c+x�. 80��_ |�C�O����|�̘w��ΥK���<�CN]\�`4~���Ҥ����e�!��K�a��"�$q�$�����n�e���>��ҽ�7��0�*�c6��'��{�M�zh	{J)*t#`��F��_�Ш+��km��������������y-J"2x��*��	v�ʊю��v��L�L�Z��(V���$�RwI����m�٘@��&/>_����}[��a��
�l*�lŶ��*�fB �K,W^Dz�X?{����(�ƁckQ:�[�A�Mҗ���Q��>�wy�<7�:(喐\�m${�G}������nnӦ"�jhG��I-�A��V#��s8�X�Rc@V��D���A������:��{=�,[�*��6���~E���Wʅ��� ����[�QM��"�J=g+Bnn�o=���;ٲ�������s�p�N$����=Tޮ�L����%����u���l�g2>�@2ͨ,g�zIU��Cڶ/�&.�Ό�"o5'���_A.�XD�9�k78�WyI�����^eT4ߢ#3Ҙ	.;��y����-����ұ)D�|H��v;6�K6&�ܞ�7ͤ���c�@d�2?��D�⪫��"~�-c�>+vB.���<ݿS7e0+�q0 3n�ж\�>C�!:����wH�rx�����J:O���8���T_ǻ;�Hh���\��!1��b�1U(o��LC꟩�#�8$?�p��-�q��`��]�������o�n��<�4V0�����B=8(���j�~��~~�^(�<�Vp��z��@w�$����ws���zlv�
�[��uWf��'��L�S���Y�����@�lmdj��O�@F��WN�J�4	�5R��"K�&���-�߷��ܒGK(_�:�-�)��i�Ă�O�#\[�-�mZ[�W4��{A,�-���`��O�YK��&��2.,�L<s2����	2�1�M�����b���8��͖�0�m�N��yn)�9�cw����*&a;bD?�ǎ­�o��zu�gU�?!�:�w#@�**<_�B��/眬�ߝ����P�v�V�+}�P6�0�HĠ���8���s��sřR��R�6�銻8}���:�G��2=����E�y@H�;�W��B*ݼQ�;��D�2���e<����ҭ�� @NJ��U�I��￈�̖���=�?�k�|	 �a���A��>)�}�y�ɘ�g�ԯo�ӱ���^WI��/�p�PF�G�z�俔��JM��,�AH�����eKYt�$R^�P�n'i�.+��Th^(Ug��:>H����ΟM&ŀ¼L��R5��4�x�?|��M]�������w�=�#���G���9�=��|�]!�<MI�H�Rah��3�KV���~�ƾ>*��>J�������-��6�c<s����f�� �W�*j,�t;���"���%�F+�jǩy9���J��	��u��N�U�0,���ڂ����r^���gI)������~UD�����mG(�����ʴ��T����>B�짦	���װُ�h�(�)�s~y8-R�@�d��T �^hK�����H.��bCͳ��@�\�.��\U�!�8{o��j��Jr�Aa�_���C@T	n�i:���k��NI%�9q��ϭ�M�[䖖�^qm�J�>D����SM7��v�0�����u���ϡD]\���6�ե;}A9;zh�,z1AGD$z:)�jp��翩��B�r�!�k��& �+�n�>7m'pfF��X�vR̈��PU���I�� C��ʨ�y�}#��'��_ڡ��Z]��\īY��]��6����e���6:���:�GZ.}r�lW͇�l%�h҅}���ѩ1���d/�����x"�]�RE�F�ݚ��D��^�W��^����3.+��t�E�]�4�$*F&K�E
��c�R�2܀��<��O�e�}���sB�����*�6��_�\f���d����q9��VE�΍.��2������?�K�taF]QlA�p|𦐇�R3�\�B�r������F�!��k�bR�1^���U���O](����8�[(�C��P*�ǵ憩�~E�b�䊤IMZ���fs�m���)	/�:�*�D.��zT"����TJ\�<^�wH� 
�1�4#����Ŝ*+�D�s�^P�;P�7Q��Ale�O�j�ǃ�fY�q��:|�ܔ[���ٜK!<޶a�X5Հ�L IIꘀ��˺c"��i�a#�Jj�E,Z$��s@�N��`e���L�� ���M��G���0_S�V���.��`aG�,�s�Tt�ԫO�c�3N.@��n�КN6>�z��� �hƱb���?��m�%��1�.x��Z�dt�-ᄣ�'����*Z��U[��@o�
<��52BHM�c�d���O��A�[M|D#�!/��Ԋ�1�'2����t�d���xu��U�!�0��bvx�]d%�i��i5�����"䜵?�IgМ%)!��OQ�er�!K���P�*Y�Hc��ƨ֡-4���]��ii��y^t��<��R@~����{_A�"P��E`��"���H���<�⥗2B�P
���y�VU���C���Dp�=u(O6dUBE��7��H��f�T⏂E=��j��	���8�{�^�m����4�lu~���gk�o��}������)����c�JX����qSO0��CXY��9c�Tw�(�m*�Mn���S~�=���B�E��UY.���"�Sג�Gk	qikM�6�L�5^=�wS���r;�Ȅu����z�?jrr�,�Q��觶r��
�6V�� fI7���y�F0��rm_�΃�:�uKtޔ˥Q�"F�7��������٥p��I�q��F�84�ɻW����t�y��M��ܗ)���9�J�0�:�Q85�KJ	Cj�I�c	4����ST�텸"dk����7��K-X$"�5����K'��a$+��<ySZX#�G�b�_����?�H��ݻc�R��~U?���X�`�*}��ծ;�?�Hf�ӄ	{s4?\�?���TT���z� Xc���YW'�qw>�܉�8���Sی,ČN=EM��Y3C��b�!ݶgKP�pB�^4#� �wUƼ@��^�dj˧��aW��w�	�Wn���~��3�~��rب0s��ע���cn�zC=I
�[��&���5z�!���'�ĦL�3���ў��lU��8���:"ɨL���;>y� �v�ł�_M>#�N�U�s�ʕ��q�ZuOh�������R����e���r{G?1g�����`F=�|-1%�>xH*D�>�fʎh�#�c�Y�!ڑ�`ЎPU;#��3�4R��1G����b=�B�~��^
��� �x ��N��E�z�i l�����bn������ͽ
ܽ��2Q���q"fp�G�o�������{8|1�m�Dݷ�f�{�q��&.y�C2d�h`.TKn���z�q�x2�}��D���=Qh ��%W�X�o4���|�|�#ӈq����ߥ=xiLSl`v����5=m\��^֭�]��$���_ρ$%U'�YJ|gL,I}F�f��皶��Y�u��̳���組h�vT����uڮ�pN#�tb����?үy9Qz��Q3b�N�֬e/��b�M��jWĝM���>�N�K�K�s���1%�Kcq�as��<��A�(��9��#q��wɹdƏ��:J�LU��qM��M���T���0l2l6�k&���u����װ����#;>�ySe��ފ��a?��:
�g�K$+g�F���m��m��:�&Q}�ǵ��edcJrI׵:X�D�~02 urݯ�ͫ��1T��,U��&)����bo�+SIi���!�@����׾%9��և�*0 ��/5��e���44�h�� @�(��72�����߻s����W�y�X�Z0Ν����[���������r��vVm!k��H~�'��P�fʴ�	����c'H���)f���(�<C��R[�l��w|ʿ��ۀv(Z��& �>c�B�F��vTe#4��'*�4o>�n�p#2�+�z�ښ��X�V�:��Ck;/�F�ā��#!�Z�g#�ߘz&��"[���b�0��]����n!Q�Uh�lf<����3�>w�^��ȧ����b��7�t�5Q�oz�\�9zJFqխ󺊹n�g=���<��&���}`�ndI�����`����h���L��շ�+��;�C�ݝ���������k ���@�[s��o�	]͉5>!A�Z<]�ǭ(��`�}�U����-^#�_�&ґg��v���9����R��+9���1�
g�u���Vl�n��H��ڐJ��<�%f�b6�,p��!G"�OeD�W&Q��2Cf���*}�O�\l�c1���m�D=���F�<�����*�y�U��S���K�D��d+�F���=X�$�=�F��R���(\#5b��}��J��JD��S-dMWq�;RkU�^5BR_��.�R�����\B�����V�!��G���G�{d�-��1満�nov~��׼�2�~-�Z�I������s�JJٛ�91{2䄥Sd �3A��H�-�|_���,�'�ѕc�<�s�0���`	}�{r�wG{5̀|;�W����i��ٚ���T��#��൰fH�ۂ^§��<!A�vT�G�XU�Cj�+zq���=��He�m��g�{��[%��9�<g���F�A^t��Y���YI��]YČ�����I�HO/���IԷj|,XN�"t��D�ִ�C��!�D�'i�M_Կ_{fƨ���;}z�o��#�h�W�+�c{W��;�v�dY�['tV�
w\����1�9_i8���vP��#wξ����W(}�+(v�x�_������?D5I��NԱ�&y$d1����R�]7���_�Q+Hf�+;N�:��T�x�7��Uؿtĉ�O��zD؈�f�t��4�'r��w�L�W�]q,n��B|�K�ʹ��~��
 �Gr^[��!�:|��Uw���:��[� � u�l-��Hl�zY8�_Q�'t''�-�=X}g�~u��fP�%��?I����#��q��Z{����I�z���{��S���§g�lq�=�j�I��[���N���:����&h��Ɖ/8ϸ/A���z�J�"�М\��(�ǥĹ�K�����vdYݗM�0"��o!�$[Np��"M_����ik�آ;%%�TR��"dJ���2�1O4�%����-���[�mD.�d���5�i��!���܏O�V�f4��R������u�:��wu����G�4���~i��ְ J����כ ܈��l��J���v�����LG�5��j��))�io�������x�9�P="����?d �S��}����_���آ-�g��"駆ȫ3OW�G��>�!�$�%����( �a�D��b����b�O-F�Hc���jV�.a�h�`)������.���{��Κ�����z'gm?4�ya�L`3t׭���z[U��$���b��$
�&�e8VA}i]0�,�G����(��"�؍�Bm�Ϛ{�=�s��e�ȸ��oxw�(�?�(��e��H���$� j0�kG3$��:(�\�%qf���8��^��4\_`�RtE{� ����\��l��:�c {�_#!?f�#qF�&�wq'�	�'R�i������f���+�S~����(��&.��@E ��{������zQV�XԨ֥7��[���������
�[�^�C欕�G�XViPo���0��6E���tp4�ڒ�$\���MT���l��X�,�����^��e��*�p�s1���[�+��(��o��xd�V����cٺ:b�nA�_=%8����k�e�]���X������S�m���j
=G���+�R�"���x��tX���"�-��P��fBW�G�ۖ/�\�wf�gT��r�}���5��k����Fi���xj��2Y4G��Z��(�B����g�D���a@>ק+�u�����Czh��y���5ט������n��|�t�T� `L1�+:%+�I,-S-$ڝ��$�U�W���u�Y����5f�tqW�.d��GB�F�'�q�il��U?���֓l8�T��8������l`�uA����c.�ʝb6����|=����ʡ-QۥH��o�d��
�?s��(��B�[Аd�G������ǝ��|�5�9�}����Wq_�)�u��p�΅m�M�\��S<��!�5����)�'s)χ<���MJB2	L�!֔�i�:Sy8󴹐��ʬ!{�U܌�ۡ�"@Ay�ސ�z�if�~-��N�?I��듉��k�S	��[���I�����ꅞ9��	�c�P�`�K7>���]z���0|đd��']37�*�p8KyQ���uq��{��P'���N��֬?�+���+%��r���W�#�����ZG���2�U� _a��^4Sչ�=V4N�8�~�M��=	~A������)��� a|���rN�M<��vCR��9�0�����7Z��p}�����݁��B=S*g���L��E������:�wTx�8��Vf��-��z�6���'�>c�M[z���'D�DP�(�B�,�bX�ĩ+^ew�mu%IZf�i���qB©5U1�NW�G��:�^[��*���	����,U,��sc��w�M���E���]��P�)	�*�AaK�Z0l����;W��?B8VW#�+�u��ZkFU�m�C�LZ�E�-�>��\�.I�B�%c����8S��4��iq��I::���v�L�����֊)Y�������η�,��>3r
���`5��L2V�_I�gs�I�k�̓�6��'-F�5B��t���\ƴA����!�$ڠ��'لB>�R�s�A7��<���)�x��SɜM������l�z2���>���v�����L�Hr�zp� �a�"%��R=]��ǚ�N��G)
����+����Nd��-{�^�����^5VS�CUJP§�1bAE����O��BOt�)��%z�eά��u~τ�'�vvv`�iM�^�tXbʉ͆�6? �4e]�e��T� �	~��5k�{PV[��69�EUk������&bK��m#�+ ����!z�z8,m�z�Ҏ@V�5�W
O��!Z��ֻ8���⩓K/�����6L_8�A��	0�4�\z����/��W�f���'[V#�Y����Lr�ƨ
�sn�A��0����r�{,^�d-@Spph_��������l��h�tۺ_IP0���OE",�M�\S��`�$�ۺf���&�\����dc��0�ʚ5�*}+�zW�|����AS��$mD����`����e���w���,�X��|	�"�Lʮ�ðF��]�I^�nGUG�I4fh�?Ý��:��d6v�F��U��5I�Y�i�;��J��YY������jf�5����*��E����������:���NnY��~������R��
E��(�T��L:�V�T���ԡ�w�%Z����ɼ�K{�:A���l��\�tm��0}?�<KkK��51A8,����S�hNԶ�+!���YN�P�$�?z�T�xݩo�{�`ʇ*�����. h���!�Ku�H���ށ�a̓mY=S��h/�ݒk/�r�+6#�,1���TEo��:�� �2Cy:�)-���>��2x���B���9OCAJ�L�j!H��S(d�92��vP��n�� �₀W�@�MZ�b� �i���C�R-VνO%�|(�{SB\�d4��#�60���M�
����h��/�Uz�1�y6��b��KV��Pd�M�#:�`�J��L+���2��S��&|�{2����кU����R�=p��O�f���V��h�����x�_����+(���y�^�aa7�Q��|DM���"dz-�˼��Ԟa�E|w;�u��wv���rD�~����c�3'��J��#�[%�-+Lȍ�5&��fL ��� Q�^��o� �1��B��I�U��Y�_5�!��q��g������gb��	�X/�t ����eh�R�S�Y�Q+��B���1�ak:!�i97ٜ�J�ʑ�PW�{h3O��d�[}��Ȋ���*�&�Sr�lpu_��VS�`���\1Tu�[��F���9�	{���:��^"*�=����y�
z!1��^������ęY4M��	c$Li�W�B��"��s	�X����ߋ�#$��e�t@�V��zV͂;���iFnHob�I׊��y��~ir�-,����Z���HZsE��N8Yo�
��޲��!WG,�\�)[��Gd!�\ڪ~�)^�~���GN�n��?;ѷSW��Z{��N����'J�5#oX3���Kc�y�ϬUTc�" w����j�T[����"����g�O��W�=c���w�e6h��Zo������r&T�d�� �R eMD�K�:0B�Į��))B��a�WG��9M������D���W�=9Q�7|�U*Tc5���+?���u���x����
�[��d^�G*D#S��q����]x�=��ݰJ�A�9ܶ�x�:���������N�\U�rͮX�2*a�wY>�����k��h�D�M>���06Bz>TB��\o��!��h�r݋�5t�H#������J؏d�{�C2Ȩ�D�/�MY/fx��>�{����N�����-b���'��V5-�G)ۂw�&诽YdQ�$����?W�s6-�0}��ySw?R��*��%BQ<6�L�3��6*w�� �Y�N�"�����L�����5�ڇ WeDUş�nf�
>��-�� =��Oy��E]i�g�M����3�4�x#�om�)I+�(*xdA����P	�  u"$=�&�3�S� �ER��"��ךX��@+`���$�Z�2h��2P���bpC�t�B�w>/�.�&��Z���ɫ�ͩ����Yx|2���ls.t3!`���{���ؓHAZB��`�)]�y'"bf_8Y�n������:��9dN��h3T����E 1t��`z���]�ڌ�芄5�S��_	�_F[r�i�|�`>K�#��+jn,c U���L�@�|׃���!&�������B�Q:X7a̪ӦӟX��Z5�ī�;?�ʛ��~���<�逾���ÿ`�Uᩍ���kS������xM��_�y�=}9�-�Y�Z�!�_msP��
+�[�1�.�������u��8�x_�����׉�%�l�LV�E�$���.(�>�)u�oN�2�ڣ�N��A{�ܳ�⿫���ήG��y(�#���Jj���zz��@@%M*�*+6+� ���M$o��8��d/[�n�U1��lLi���ת�����xO��2�k;���0�*����[�������}. ����J�o}Ǭ�����kxLV`��0t�֜�i�KR⌙���mI.?�XQ���i!`-s�9�ќSzx�)m2����ˇ��J���"4�V�ǔ�*J��e�a�R�"~�;�g-�}L�4S/!�Ă���e�C=5;:~8�= h��S�0mh���a�Ŗ��N�T�l���~��6����md�4ޑ�)4��]��YCـ�R1���+v̪�%Y8�a[��'\b�(�6��j�)N)#���p���78��ȴ�ޚ$ 3T͈�A>���`�{$�
z�5�+w,��n&怠bF��T��	!/���Fh��-|�W�p���C�Q�a�G�_ ��a���H$i0���rf������0 �c��ayf+~г�:�)�A�ok$�ND�P��&�T�eՅ����-�&h�s��ʧU�I\rD��w){�>���ӣ<:�\u,qW�\���t�	2���sq���x��٘Q7Аw�����m#������0z�f�YI(� Re}k��N��o�a�xMD(���l����yg�	u��L��0�N:��?$]�[-U�H��T�����OS��:S�M���q\ʯ|�٨i��Vy��S�q�N�bjc�7����H�¾�S��ᅅ���Y�"�uY�]���w+u�;d�T���
��;j}�j>@��-'����IEJ��/��D9��_���>,�WE����y�l
���r�Z�R�RO�#�8%p.�|���W��P�l���zu=�;W�\�tz��%Ju�`F� ݿ��	��}����
ɞ���|G���`�Q�(̜�6<S���z��
����^nj�fN�̲�*���
��c�Hj9}2U3�Fd�yR)�v��?�b�HXU��S�F���s�h:�\jS�FZ�B�� �T�.�U.k�!Y���\R������Ŋ�����ޚ�r6�0#�/F�ɇ��?��8bd�\�9�C-UF7�$����\��N�	n�3C�L$m��g�(��ෲN�s �M�
_.��L�ƽ.��\�4�:� ߋ{�����>Ue#��U�5K:� ڇ�?d�ejr�Ex�������ɳJt�J�*yjj��A�uER"� &�M�!��Di��~�,Ż�Ct8����pU�7	|�^�u�@��P(�S[��n`4��5�Nq�+�؀dF����0�����"�hH��ƚ�b�Y��_|�+�,�醾�lhRp�A����:V8����q��Q#�TyNy��!$V�=�+1J&
����	�6s�D͟��߅5=2�E�[�"Jz�qD4/�M� p�yR�8���FcT�(�dÿуv���{��zU��ET-=�<D��,yDp.w1�B
�o��������_)��γ�6��r��G�ǭ��)����x	8f�}:\�y�d����0��BKa�Fu�r2�,\O��� ��\����_@��j�]���/��b1��n��>�[٭�?h�o��丸�����,��/�\��q�a��N����<�mu����b�jf��7����4<��{��3�8�C��ra��y���pU�Ec[�J���g�;���P�b)~=0=��7��E��,'��3���D�@{C�e���eׄ@�*F���.��Y`8h ���VS]��u�5�TV3��>�Q���d�#��"�Q{�jϭʎS���sJ���}A��ɵ�<���j=3�&G��21������ǥT�mLf��E�ƺ�0����PcC�M(��J�%5*��~�	x�9�����ͅ�#ِ�$�,��#�lR,b@�@53ܙ2��N�$�tr�02=�+�,S>��'��.¡�B�3�.A���B^�1ںͶ��%�>���uId�a�b�Cb���p��h�r3���N_�#W�g592q�j��6�԰TPĺ�����͘ۊ��_儔�����	i��s�?߈�ᩤ�4�\�eߎBa�U�/�H:(ö�D<Q�q^����5������`�!���%��g+
�i��J2s��Z���{��p��5�j��=X�����{�	9	�Db����xUD�u�^7|ؽԠ�牜���E�ɉO5��A4}�YyŠ܊�`��ro�tX=-õ´|��)`�N%7W�$�7�5�Ar{u�q�m���R�|����<߀Aں�]�=��4�cxq�sRV/k3y�J���c]�˜=*G`�m�䞑)����D���D^d��!_N2�!�X`�&�NԌ<�8u��Pc���A̣���F�~.�pem=Y�H�U���@���?��BFs1�q��K�������ꨧ�N�+�S�y�1�o�UpWS��K�i�5��*S�k��,ŷ�<�זp\�&o�n�W�ܷ�7$�'�ů��аV�\ ,�(��,V|�R^E:d�]zD4��IÅ������D��U��C�0�ZR��"�CW�'�J�(�ƅ�lS�m�<=�W/���,W���籝#��+��\�gܜ��c/+q��[�W.,�Fاz-��pd�x��(B�����6`���%`R�k>�e�29��+��	�O����.w��4�eJ|��;fֿr,V>�\���"V�:Y��(�
�Y��~�?L�q�3iSx8��v�x,8�ɱJd�L����~��"1�a� �����)e�:f�~�|�`/hB�q[]#��D�*#LBo���������>�uDγ�f[Pq�^���dL������sT�)&�	��CG	��qyኧO�И�K�:硍9Q�D��G#*�_xP�s��\e=+��T}�RJǆ�8��$]�%8�������o��(ʯ����7u��g��	����)��7��4l���ׇ�����[��=YG;��K8(q�r�ZN�����w��Ų�D�>��
�O�o�c�vLi�X�Qz%�n���M�B�S�-V��p�(Si���*��;��*�wV�~�?�!Fk�	yM���,�d|�Zt��a�P�j�KwU'�u��W�h�F��$- ��r��Zt]�w�Ct`��\���A��|?������h�vk�F�V</Rr&��p���{���ϲ���?��,\�[�1&�F�2���]������n��^�L�3g^*JV�;��mM�� Y�>�v�7�M�hw ��`��qh�b%�����9���,1r�9���ms�UUM�dz|��,�]Ƭ��I�!Wv���<81-2\ٻ�ga=�|P��RY3T�;�
�6��\����w��$���j�,O��C��8���g�
c��Sr=ig�:�F[�gQ�Y��
C�	��ojeX�@�8;���@�&DQ\�.t�(�ҜhJ�Wl�N�,�V6򗪑$�k�� :Q����F�q<���[/C���x�-8��k[�Q?I��V�i�V��;���A-���wz�fx��P!Q����BV���<,�+6��S�v�d�i�EA۱��yD��4}7Ќ��:s��xg�>1l�e��Ͷp�Tr�k��?��#�U��Ő�}rb7L�bU� Q ҋ�t���.�6�hr.b���\�l����%����Nӂ*�A��/�Lo�)Yf�\��	-$��0��f��Nd&�@�l������2��ė~s-����b��"kᯇ�c�|�.�=���[+�x;�6��H?��7=%������ԓ&�*�D����>��Uy�p���b'h�ݛϏ��j{v���p�����%@*���9����v��GEt�����L��}�6�~O�G�Ԛ�֗�|���gAE0�9��ecJS��'�%�1��}�&H�n$'9�q����^D����i�R�apo��U�k����P�XOf���cn�0vm9����h{�Mt����2ޱ*u5[�����[h�<�e�`�����We�BTx�y� ĜK��Q�u���������I�vZ$2������R����a��R>LgkF2*�L�LL lx��d���3o��b��e��k|�m���H2%�C�q�>�!J5�	��z�;��Un�]���_�8 �>Q���C�9_�`�P�_����wJE�٫�ED��ũ���{k�
cw���黗#meMk��l�T4u:s!̏,�~���:���R�O=���䒑:ns��B|��J��r��k�@����A9@dr�4�!!�m&L�y����MS�|�D���α�i̐�T��f�H�1i�]�L#�0ٔ!�ZT�<.����C����� F����!��lcGɒl�a�^.R4��ܢ��1fS���E��]:F�+~\%�a�ø.8I��J'�ş�I���z ��K��W�����Z����t��WN�c��U9(F�!h.r.*}c��	�E�"�}.Ԣc�6����w�ͩq}��9��5�*����e2P�-5�hN�Һ	�TO�#�ӥ�`��''ߺP��Xt�J;L���:�njw,.��
�ΆJu����w'���7y7�d�:���NOɓ�̗������~;���(	�+�fs�F$�f�7�b����P�W��?|����uߢe*hҒ���aٴ�ftIk�&�X�1Ţԣ�k�n�8*ت�VH`��0Gb0�M$ e"�~�
�py1��F��u�����H�����۠��@U,b2�i���S�N�4~D�ϺA��u�O�MK(O+�[��.ǐ���|�*��K��V��t��	z��8��K�8ˑWT�D�L���W�Zk] ]>����wӾDLcCt �\PE9��{BxD�^����U�DZ�ִ�F�9�������g9�z*�Iv<#���~N6�!��`�Yj�&�1�/գ�e�ʍ�v�����Q�
nF]E�b1���8�.�N��=7AY�b�������7�=!۟$������7{�՞�׳I����Hg�7 �D�	�x��ij��JzY���B.�c�D�q����`���$�P�<7U�.�D��uͯ0��#J���5o��?rS��؇�͒5(��)��?��fFr]�N�ƕ]�� È��XL�l�"� ��ȩ��ɫ:4�6W����g|�������p����!e�OY����� S�q��k"rƞ��x�������oS
�c�J(5@�z�.�>�Po�_X�{UX�¹�p�a��+3�=j@�.�I]Q��8���O^�Y����z��W��L��	MU��w����f�cS��ۡ�lx�8~�*�9L�O�A]\5��=vv7m�<N����jn�A�Х�1�x,�҈���X�`�G��LԀ2eq׏��r��˃=��=I�s��.S ���qx�`��~�^XM�z��?�-K�;zD �B�3��^�<4�g��3@)�o���K-���0�DE�c.�54m�N����-	HF�0�4	d�F o�ঋ��#n����m:�W�d�,��f�.��Ȫk�={����� .?]7�P�?J�o�5o�(���@�ז�����'H�v8~ߦ�>�AY��i�s�H+�]�H�O�J� ��.J�_�j3��ގ�[�M��}��H��&	�<b�a�?�lX�ج������WU՝�m
\�B,�Jz��&J>�0�,�+ ���S�jv�7)u/��J�RRg.4.粛���л�Z��pwv`�W9�Y8�x!�ԌBc(��4�b���2�X�{��&����T�d��#Օ��E��I�@jd+�2mer�����}�{l�����S���L��kҦ
�y���q6�3�*G8���Vb륗ʶ����5결���I%g���,��_\��v�߯WK��0v��%�(8� ��M����h�8�u��@��1t�R��<s+��.%��Z�h���N��(�;�F~"퉹3�V��\ǝukޕ�`��L��P��_����%���TyA�K ^{l��`�Hb����9�V�;m����~' ��T�rB�z?5,��H������o�n'@��B�K����u����o��?��p��-����1�$�I2�"�j��#v�ϥ��#���F�t� 5��A������-��\�E)z�y1*�V8�3N=9�>3=�lFw��r��{��"C�bI�9J���DI`t
4|��+\���[�k�����:{��"�x-�j�ÃlX!V�i�X�~��[Q�)'�I3��O0F��A��7˘EB<�V�Vq�n�/�G�z��8�ٵ��LO��}�E�P76�'�,�W��vd]�h��<0_,��9�\�X�2Zp sB�Zi�f��6Mx��,G�)�ygÙbq�$���d��	:@��u�U�oλ�X7�i�c#��qR��W���l��iu�Y� -���WN`Ï��Yxb�8�T���� ���&P�\F݊y;�amB�U���)0��^Ŏ36$�.�j��!0�g��<��Z�R�g�����D�k}=���hk���R�4�� ��cʿM�*�l`�@Z��
m��}9�����l,�'n�g��ɨ����#�^�ig�%"��G�!�ԍ����D%�WU�@m<�Z5	C�+H�0O�>f��d�
џb��aqY�3�2F��<N�1@MM�j��g����8&}(M�`-ۑ�3��+툫�����;|�g �E%;��[)~n�/}dl\��$�,�[e�_���8I����u�	��z�
b�q=�5�ïdI-��X�u���x1��\��;!R��H�.��l<���o<������;�:�<��cZM/ڽJ8���ha|ê�x%w������}��p��n���
��[qp4<�I�Q�`���<^0w���%r�MVm(���ez�W����r�_+o�t��#<��A�����u����������^itK[���|���s��Պ-h#;2�����M2`Z��!���ڃ·���@K���k��Q\���ڑ��4�����0B�h���#�>tY�jL.��i �����g�d-r�Q0e T��m��O��z��
�UC�InflCv�m�<�:R;�8ڶ���E7TGgȤ��
��{p�A�)DF��6���v����` �^?���bfa!jJi��Vo9�m��sy��7Bϖl�<z��aC!�$�#���ö�N@�f��pr۰:Y�P��5}$Z��c5#Q�I��DJ�V%�XS����8��t��ı�`���w~m�PI�]Π�Z��$ݿ*WZ1񞨙�ͰY���v��#�<�1dz[��"K����2�"�3K1O��h�s�O_ևFW/'��c�T��6���@��-|b�<0��t��z+�}�@N[d��5}�Hq��ن���B�|F�S�p.i�5 ��E��F,�ݍR�c,�O����hh�8$=�68��T�l��{}���%�Ol8�JCy�����1�c��2IV�px�yu�� -�VnM�0��(�ɕ|���#�|��p}�?�X8�s��wd�vՈ�CZ��Ñ�JC�X��It��;�4���m�r.�-� X����fuz_.��5�Yjv�>)pᡫ{�y7�7���7=���������v�~��������C�d�R�;2n���֘`����V�^i>݌h#5�k��Ģ�А齛U׳u I�*Y����/�F�ǟR�5+̵�/�A���;bit����P<˅�7M��0�PI+�&G����`�*��T�:��q��s��2�b~�3�;�'U��#�oɇ$��J�)�����^+���Pj}k�N`����u���7�Z��^
�q�4��0w���zCӹ;<�Jv�(�� ���q�B>�����g8Wr��	��dىQ��eQ�ԉ�ǌ�`�H�#��4�j�j&��/˽����Y�C���,밌tً;�ĝ:H��Y�!���o]���F�|"Lv� wbE�v�-+��u���,��ԥ��l��ː�L)7o	�2�É��Ck��Ɛ� xL`���r����#o���DPȈ��W��/�7u�G�ci�;?�+D��}+ْo,��bB��8.����xr�z`l��v�X�V�@�q�|g����'���h�jR��V��1�7���}�Y�+V������T�����V�#0L*8G`���=����Ce�eEs�؁8���,h��!�s�>��@�n*ӛ� 8��7h~N��y�H�V�&ك`)�1����^��?F)$�C����|�fa�S5���z�G�Ė���q�����!#ӟ����Ev���� j�����wz){�Լ�A��`���$�(U*��I�q��WHq�ɭȐ;D�=����Z?N�.4)�O��{w�a@%�u�?	��<h�`�2��>m^�ܜT�ZQ�=��M��D� �����TâB�p�����.6�<�I�P8����-Hrs�������q�3�Dy/�$�KC|F��zњI��o�Ֆ�?a�
����5����`ҟR��Q�ln.���+&⑸�l �v�?!�O���[_��Cp�4$ʌ��SJ5��!�i�ڏ<^�Ԇ�V��t���.�u߾� ��W[�鐆����yD_�� �֧�Tj��L��e�@$�@t�܅./�r'�	D�<ʲ�k�b�o�c8���7U���F�9%�D�<Q�/�N��GL��Ɛ�j�{��;�N��3v������cO.$k~�'r9�����{X8❢�� r� cdS�$D̦�t�NJ��`wʟ��{�K��G��u�(ͩ"D[_;�4�;�#���jy��,͏��[��&�e�G�xN�N���#���e��J~��xR��t��9#�Ĭ�����}�Oe t�wJh�����>􋉣5�o��w(ܹ+������8�A��<�@:����Yo��]s��/{�Ќl,����1!RD�;�� �t���0�=���|aB�0C˟��KX��V6|�0T�Q~���*���wIۦ��T&��>~�F��j�Ob{=�]��oA�˃���*��r��������a:a��X��\`K�)W�qCQ�+QJ���d��+f��M)��u%�����W�f�'���4t�ӣ�WZ[-�6/��#d���ʹE1�o��l:$Ux��g��vy�{H������_�#\rt�۰07Vc����0R��T�����M��I��;�aA�{o�,�|�7N�,^�'�\���x�OU��<:x��R�P	�m���"\�*;�~Y�3 e��r��iN2�Ş��W�$�(���>e ������O�lya�r�����]��{V����8P��c1C�XSr�mj��y�=�_��7�=4$���j0��2��}�i ��Av"����.K�\�W��|7z�k��i4��Q���Kp6W���ZR�C 	Ԏ��g
��@B �#��pɔI�Ȍ^���
��o!*ߥA�8��&�)vU������7��{��0�
u�V���hy$\�P�v6��y�#����>*§��mq��)mK���$��D�f�X�I�%�x_�[_�{���F̗��HS$S��	6Q'`��|h3���a7ʍ���W1	�(�����@����h�(�"��Y��W3c_��&�:�D3g;=��1�~\5��o�4��
�u��XFh&+)*���"Ϗ�x��h]4!Ɗ�| �p"{ʜt��x���'%���ƙ<|b��C*(O�/zpj-s��n.@�D�̣u�n��[�?��0=hiv4��K��<���5	��"�C�B��V����怹�� �`�(f�F y3��1�N���
�z##:Sh�!xuZ
,Ew�ȽĒ���a��8}]�Q�����U��r�ş�24E�3dXI	C=�˂��4I�M�XQ
s�&֊��v��\D/����?� ��^�=�*p�^�P��Ƀ\]z0Ο��[^����Q��PP;U<)��d�p����=�l�C7�VU�Q��jDZF?�B�T%�i���f֗�{F�<�;��c}����UA�UP�lˑoB���)?����C푢�{KY���K�Z^��@o�jmQWEX�����Mj6�N3rc�»E.oM1�z���MT��T�B��t�&��Ȑ����=�qX�38�h�*<�Ȉ9$h_��%�������~�>��<D�R��/vSe]�\+@B�z$@!S���w��~8�΢�1�r�q�iذs��H�7ȧt��xp�)����(A`))E�Y���T�Rr�m�c���ǳ���@7G���ׅ�?J��QK��sz`���W���eZ*�Z����	��fR��v:�<��ty��poi�AQ �VN�U�*=K��=�kSdf:��[AF�D�G����|x;�Z(��#�5�½f&����������X��0���=� ���k��7�.e��1�pzj7�c����.!������O��ڙ��SH��5�P�x ��W��Y�Z�����9��\����I�ii}WK�;�u$�Et���\��/�5.��H� ��x�1���4�	��x>@��P��J��n����c��Us�A�A�lְ5'QP�#�9|}��T�y��V��*���!�L-��,�i,wO��Ĉ�Z�һƅ�%��v��!GQ!*����a��}wՇy����I;2�Y�m�8� �L�^������ ���e��x.2�I���D1 �^*��^���8]������Ȧ
������������
��X��[�v����Ζ�T�F���Ͳ<̖���kQ��&��([���uͣ�&�a��E��h}��N��31��{4�6��S�t�
��~;��}z�U�g�����qq��f�9C�9��|��7c��\��<��/L��u�V�P��4�:�E���e���'���m��6z��.�@���E��s9K��y	���Q�ig`H�d3�@ǜ9	��Z Q>
��1Qt�)�QL��(�
���,��;
�v�9��5���8a���\�p�J�F1�<z�����_���z�M�r����}Ԓ�ْĈB�9K접�v��b4�����101!������㾱��^WOt!�.`z☞�1  ��YHuؿ����)�p��s��C����>�K�9Ð~���j��2���x��⇀����,�w&�?v�ƞ3�Ȣ����0._�@\�s�$~!��Цz���>���
f��^F��vT�Oc�����iY{�y �������Pt�JK�2���3(ӫ!	8�g�0�[r㍜��n8I�x���k�E�vz�X��k�P�'ui�O���j����h��c��O�/����;�bf��ۦ��m��3�%DڧWn�L�p���� e���N�a�\�ր;�.������Ȼs x�Ŕc�t��C���Ki�񯯧�����2�Um0������#�����z�{!��fYC%_�W���3�� Z���H,FU_da���_@�98"P�n�"[�ǵO��.�Y� qL�^�=�/���,�T��f��*��ZŮ3�2���oU�=bc���̇�Ƚ��K=QaUfO���<GO:H�KH�&0���K�hn`|?�ɣ�oՔ�c���DH�l�����rV�/X-b���+��R�{~�
FGj�����^����jP;���Ź��[��%*vb��p�3��^��
D�*]�?W�G"*,�@�`�������W�����/�f^v{�g��=LS�ϊ�'��w}�� ���o�+G(��.`|����|Yi�
yPḋ�GZB�xT�L6B;� ņe�v7i '>W&v�l�H�Ln]!�NM��Z�lP��SSE�����x���iש�
4��7q���#���(��恳�?J�xg�uW۹ T�n���H5Q���^|>w�M�D1�j�x�m�e`J��k�T]b��riȨ�΄0h�]-}�؟��}�d9��ݱr�iǸL�Y|s�,s˯�|5���'+U;��O�%�SRR����FL��uЭ/�BdT��_���z�,�C�ΨA�C֗C���h���@������y��O�sgR�5����?�����Z�C�y�Q!3���R�� n���N����vRrԖ�A�g-7�?u"?�E�i�H�?.x���m���Ӣ���c�f�M���"Tʳߑ
�M�T!������Kx��;��+k��TZ.���5-t�`\�~�ͻ�<<Ǧ2-+�_� ��"H�1���d���p��gC��}0.A˻�w*���3�M�)����£���f��'ڞ6�j_��v9�_���x0���o�5S铨ĶeGS+0�,<���U�_�ֱ��u��� � ��+
�$j�F�K���}�N��~�/�b�����{�Xm�!p��+ۣ���c�ad��ϣ��u�A%DL^�4r����m��mC��5&`kjH˛,�0�[ݯ�u%Y ��
fh�N�M"	e�F���dꛈ�p>�YNE�9��/9��h�ph�S���t�<��;P?� ���qoo����7��H4�}��U���+��!�2���q匴��䕥R��w8�(��:�����(� ^y'_r��ΊT
]���;2�`�*/��q�0=�*�p�j���j�G�5�I� �70��-���Ue�Z�Xc���=+/�����d;��k{ ��9PƦu׻9��:U�N'�a$��T]/)����<b���j�k�0e�q]|Z}������������J�{�L�Ӡ�����{�f��˵d�%>��j�Eh3#��|��S�n�4�>��9o_�DI&�j�� x'6�%�]N�4C��f�et}?�2}�=� ����e� /PU��B�:N9>��	|�뮾���pdD�ow疡��$8���a6�T�^�
V
�"����&̧Mwg�H���!�����k'+�אJ^��? wRݩ|���j]��aD��خ���d��M:��Mzk&y���U�>mq�Z�~�%(�r���Z��#iq�
̨G��G�D朁��w)z�U����0PF��P���B c4�p0�oi�m�@ޠ�W2�2��-��B�,�l��.S����A����S<�~�"��8"�{�.8rI��q��;�n��m���m��C�c۬��dM?]����b���;���E���s����wf��E��л ����۳�����"^��vt���3m;��͹�ND`�J�L$��`�̵���?24|��,A������6m���D���`2j�z�8�a�3�	|P�dJ���4xr�eU��s,��-׻�v���b*��q]��q�^�=MJ��66(��w��j�PK�RU���c�/<��<�/pL��y�(f4��B��E <@%-`o��5@hCz%�ti?%8u��
��e��[�3y9�U�
B�\���Eo� P�_C�����/,5T��ѣ����u�,t>�����gDs�8�&�"w�*}w�����NZ�&���f�R��)��u~���}Ō٭�倅=XH2C����pJ��v�6o
�c�cy
���s8]=��Zb�3����o!�\�g�;6���jq��
}��F��?��q����
��E�3��j�:�7FG�_5�����U�$��� I�B#m\\2���0����1h��7|���{��f�ޒL�v�+�3|�詯z���#�p�p����oAY%�>�kh�'R���tѦ�)�jo_�OπΈ�$����`���'���[i���}�����vm�w ����	J�#~�� �L0_[��'�(w�Z�_��`�`�����
��ɗ�p���M`u��4uk��zس����g֦W��������xNY}z:ó;9�0�d����׹����wx���1)�L����-)~58�9jx6Y�I7(�Ơ🸅^Ll���]d�5.��?X�#������[20<{�e%��m�E'�:��:.$��~��{$,;"QQfW�����x��Kv����9�9�DΧ��e�%������&e��|ƈW��x㗴b#=��Q'@��2�4���c��_���`ӊ,����6J���j�[]��5�/{�V��{ղ~�����MN�U��۵���b�ޱ`�=ޖ�@}�qmt�79S �U�O 6��1'癴<>� ��꽈��&��|35V���N*�@Dfg,�L��~[;�x�&0@5%]�[�!��@m;?5ì�΁.$�|<yf���?����?4��,"�c��'u�i��.|n'��.6���q[�+����op�R��iƄ�P�)��q_�Ӄi��8���cqG��%zаq6MI\r�{=�׾�o6ɵ��ha[T.�,&����C�x�e�nы�A�.��E빳����̓�g�����7$	M�A1�E����'q<�|.�O�,�&C5/���w�ן��$RZC���B�'N���Cpzd�=&�֬��c=��J��odoX9"¿�P	��J�Y �f����uq4���_��-�!(�����n���1D�a��6��T��;N5d|6N�	5l�����e�^���O��,�:)��N7�Υ� ���i9ao�;<�+����O&��7ݾh��g�?���>��i?Wke`�mM����t%�����K6��?�W$�g��K�r� j6��TX?��h�^�~�!�c�\�6���`��t@&ޟɒ;/O.P�,� �dԯ�����Da�q�
�c$�c�ij<"�9|��Nښo@2\=,~��|�0�=,?����74�'�#�m�~[⭞��u*��k��#�6%b'$$狱�ҷ��6�үT�j !<������s���D�����n�J�&��d��9��'�3Ul�e@��U@�o׺A��8�7v�)?�D��(�;�������L��9(*�+u���M�B`���x��󥪈^����Ɉq�j�r�
�B�SŢ�b>��4g1��se٦��(�d�����~~9���B�>��_�g򏔈�b�Z�4��Ij]g��r�>2�<F�zZ���LL�����=���g%q��gr�`�
D��%�#���������b���}+9��@��H<�����d�:
�~{��l�N��7���*����3��q��p �����7�w��Hi�BRt�q���M/���_�M��v�%DgS_��"�j&>��L!������o��L?���>���Ҟ �ܘސzv��U_xZ�sc��N��6:M��89h���ȋ"4=��������ϱ#��jsz	T>�Q`�2�b9��Y����$W�ʘ\=L��r��4��x���n3��>��B���ǳ�ͺU��0��7��MH̶dd��͉k��:D�(T"����L0D����k�-Z�ly��Z~�|����
;���ø�e�$�ʉ�Xu᪇J((�f��ι}�֞Ӯ��cb�Q�s��
If�9��S�h5�uw�8\X=�����H�g�ݴ��	[�Ր�����V:RBilc>��>0���D�^'=��Z|��dB9_�����$Ŭ��˽J����t��������g=�ʡM� |{����]<�X�%;'G��^mE���f�̠P���/���NN��	U���3��D�������ܛ'Zn�93'F�$A��2݂���E����&䯻��K4"�}8�8�(RTx�b������~%wc[���&O�1P��������+�-4o�Ď�z��yt�̢�HA�+�a���Q���8��io^LX�����o3r�أ��&���	I=.�?��n��z׎�$W����c@i�D�a�G�����;m�X�~���
�/&Mi�(�A�}h�����w�1^r] `lʀ�������>��k��(v&ҢZ�Q
����hS�����O9n�����a��g��ZP�+*t��I��r<���P3��ҳ�����G���^!ͬ��j�mғ�~�|���aL�nL>�b�g����Z��/��:�]�|�J-�a��g��i-�[WJ{���ü���F�=t��rL<q5"��.��ŌG����Mq�X�$�>�YС��P�Hc��O�� Z~o`�������Q�a��(�(*c�N��H�s �Y�z*�0���F{�݄��VB�d$�9_�T�ɟY%Z�.�ܸ�-�HG��,iIɸ�����>H1-b�n2)���c��x�e~m�&�+	ĜͶS�wy��2��K0H`B��T=zPP�1���e����	�Y	uC�Q>��x�w�"����}��Z��W^��B�z��Mz8��%��C���1О!��hy�n5y�!�wj&�<R�Liq��t!����5�����G������>��t�7��9��"\��W����n_.������:d��o�F[gS�b\'�C߇N~mߍ.%m#��0�:�1
pm�h�5p��/C���W`~�f��F�Ad՜�O��S�sW�D)g}�/p:���]�=`�yަ߅�i��J���sx�?�{�]]��w��a��H����@�k�(~�&��6#�]���Pvy�����4�[Kp8_��t�E�v�x/���l]?���[�Hp��,q��6[Wo��Wd'�ۅ[R��>bS�K�s�{v(����{�e��.Nxr�d���=SW8≊%����S��v���C�RL4zJj8D��8��v,W%�OC<�v��I��Jp��V�K����#� _耊��CZ�]���ῴ���F_�fW��ʝɆz-�K$���dP9��j+ 	ћ�@�����N�׏Ѩ�E׉��l��r�i������`��u�b%*�L��cH�,ˉ��uaT���ߞ��.����mYu��I��
g�T�w4��L�_��aN�g�������A���2{�s5W�g �/�T@�=���q����W�3�.C�r�}��-ڂ��8��e��R�>{���e���^c9��	�*�0d��]I��1�K�}��ȎI�t}qX��[�y�����=J�� ��X��}�F�Xq]���y��1��x;��br�4�o�p����1i?d����)�_ve���5��V��'���@cZ��w�d���-\-ǒ C#/.�:�g~�ؗ���:D%���cb����>�� NP���榓N���շT'o���B�������ovn����OV���\oD���6W&8��nRs�J~����)����]n9��p���@ˣ��	4.<Լ�HcY w�����N��l��k�vtk<�;r�c>c6f�sx�E�:o�PWnFg@Ew,Ol���6�OKq�R<k9�+z�Th������ �u��ݙ����\�o�T�A}����f©{��4-�2w�����uo��=U����rx���Z������