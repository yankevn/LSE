��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~���n��$%�\V��d��NS���p��@�B���!�B�K��a��O/Y4��u,c� �����'�2#�2v��u��D<g�H'�,��=��IݹjA/>�+���+� �/I���9)F���ИW��R�����}zi�CǿG�`�@���s	� ��$���a��sv����\����0ψ-$�����a+Z{�o��<%`�m�_go�ŒD�Xavߣ���������"=��Zy�-	>M��{�Kĺ�zԭ��1̦�<w�?䅍I�f�L�r�N��1��I�;�NC%I�wM쬕)�������x� �떏�i3�����*�[�|h��[QQb~���������[��rqޛ
4�/g����1X�D��=g�����=���遐G����X��@����\f�Z��l4rXE&��������y��B�{�r�Ї�dVM;ބJ	�M�Z]y	�[�FN�U���ե<u=oj���$�iؙː���j-������׀�s��~ �"'��i{�cf�ɣ֋y��%_B֨c����ēh(x)P��#�F&�nx�� ʈ@�	�߰y�>8��Ԫs��G�g		jx|Ys�.8`��u��R�m�T���ӀPꯊ�^[�*���j�NPN����T��+!��ozO����Ļ�Z��6�8s��G�j���S��A��КY���j�S�`�� k/6d��������R��>eR%�<��3چr!���+j@�Tb���#"T95N��F+_oU�ϹlJ�Q���F�K�w�l�M��\i+^m�	)�W���~{�Q��P���n��7=���xQ"� /�ubV%�w���Hlw���4I��z�xǻ7���r��3 �s0C��u�ٮL��ź�������J��ܲ��-��y� ҒR�mYft��`aY?�o�a͔#�LfQVKd��A��y����	)�%��h	;�I��1Ҹ�QPn��H5\O��\��Z���.��Unb��"��\��P*v5ĥ��'%o$t8�Y����[v�*�>U#��)tɰ��R%�Μ��Am��]���dCd��ؕ���ޘ�a-�՝���������L��/)]��(�I���E��	�;���G$�����P5׍�7v^|^�q��i�^�\��rp�0�a*3p�a�`�o����f{������X3��c䫯)����ȼ�ٮ���@�����G��U�ˠ:���!�q0�%�%�m-g)l�8�	oI�V���4�]=��M(�VOA����;�5���>�`�	
_F:o��j27JBb��DxQ�!��6x����_u>.����Ȍ���;7D���@���-\oϒa�.��|¬9�ޥ��.��(֯,B�+��H��$�92ꓫ�=^���8�����!l�u�6�G0���A>~����J���6��^09-��9��)<o���@i�~�3�c)�7)vs��3�?�䃣����?>g2=����/���t�X��}�i��p�@snj���a�d�h|�	�N�N�$A��\K^�f[,K�ՃlA@k�I��M�+��Ue�f�I �l0m�����MĐ��-%���(6;����$xCn��Uq�E2�K�_VÀ	�:�'9��dܣ���gJ�A��!r>���x��$��m�i���B�t2���kKKj34����7�ԡ�t֝P���!F�p{d�����H�Y��]��4�pj�../f.���v��&y_�rq1$v��X��DX,Z���%CW$�Fܙw��:�*);[�r���u$��/�/��8��g	�G�L�R���`J��H{3�leC{��������5җ!J��[��Z0��i�����k�?&���c�K������,Th�b�嬱se����f�s:Ux�TW�D�*h�Z�#�Y�@�a���3�f?F>�</ow�v�ǥ|�&��s,+�ޮ�"��`�`9|'��Ǝ"*utgH��%��j6I��&2b`�aľ{
��(��Ba 5-��������2�Դ�EhjK��,��UE;7��6��9�L�Ǌ�=z$�%�� ����3Q��tL�K�sv�>�ys=b��3�e�,*U��_#�2���ɕ*���޳|ԝ���sb|V��yO�(��� �t���x�k�|{T6b��5�C���!���2à�aİ����	������v������
o�<�2�&|Ia}g�?ۊ�r��O��U)J�,=�3� ����lP�L��>gf;���&^���q* L/�5��L�A���G� �jB= ���%����{p�7�\�
<a,���a�P������"V1��01�{nѾ��&���?W?��|�J׳<���U��3����2�=ױe���,���o���-	W��� ���^J��gZ��9�EF�:�]���������'��Fu����i�tP3T�(��<3Rs߶t��~����S�Nq3M��=�������ކ����[xXn�|��|��M<�j����mT��5���Z�i��$�0��
d����c��Zr�;2�cL�_�a�~~�/ ɏ�P���N'N��㿴�ǀ_#�diTz�02D=c?H���(L���{��X�9W-a;�m�����զ(�ǣ��l��N���ݴ��Gwx��UC!^�Y�Fi����ƢY���췋sp����gH�͎��mr���I�j�x�����&&;�h�!�%YUS�:������G�Ŝ&+>%��C��<ֻ��u`�Htq1Y~Z��;��nX0CgZk9-X�'zW�e�Z&x�^#����(�K"�su|;V[�Ֆ;-�-&��5A�ɦ ɠ�l�֫eh���^�Ώq�\�
�Rn��د�P�b�]����&�N�B���C���\φ�ig�Z� .Y�Ɓz��Z��
����HgTP& �@1���lP��G��4K�3f80́9I(䡜 �ހ�S%Z*�h�w����{���m�:�fO-�2�1�l�V���뤱��չ��iO��!�&�s�3�3 ή�%!��}C}���,��p�NV�9��A|G��fv�_��l�&���٩���k�v�9��Q�2���H&zbg�Jx��Ӎ嘡E���j�MM���:[��q6����#�طY+�ư7��<'�����R[�Sq�k��	��6�?�d�[�ō��`�:Y�HSO�pR���M��u/����1����/����Y��9k��,�8J�Ux�(z���W�L��@�;I�DK�,q�~p�o�H� �?�F��"v{�kF�g����-������*6�|iU�?C���XK�	H����P48�$���\�`SØ�3��ퟟ;r��P=�q��^�X���)���_[�d!>���R~�RZG6����[Ѝ���]����J1U�����z75n�vx~���-=�0�����O�Zo'Nd�֧���i>Ja��(��@�"���I������)\4l���#��l�	���B;��	�0�����X�����p�iݪ���ި2��Bc7�_§�z�i�|�f���n�U3H������� Sl9[_�8�D�!���%�a�z�L��e�R7���ZơJx�3y�$V�[�v���F[P�ɧzL�l�����N�#���Vm�]S[�/�愈"Es� �{���e��i+F��ꖀUƨ��N��偦C2�a��?F�C(^���D�c�/mf�8Cx�*���+B�\ zm����u��ط]+�;�K/I�L��]ov��}������9�4NCM�d�rS���ԏb��)��M�)o`�Cl�l�rv�݉ݏ��D��
�P�&��~��rځ��(��+�ۦCqi�L�vF����ԺE�Q��]'�\ ���w+���,7�j'^Ϲ(���K�0�����\D���j��3;���Tg��������xm�RQF�w�$Q�I�z�2zaa��>�\i�U��q%]�^q�d����%.u�<$��5��IC���z(��l��c�5����r�OW�OxW��#�1Qы�`��E���RU��"�~/���?���ܩ�FM�p�LI���;��nU��%MĄH�/��\�P��t!��qA@���R��pA��ch����ޱ��	*@R�^�����I~�>PiY��a�`)�U�Vjz���̬3'�Ч8��<ض��p7�tϧ�$��Y�ַk���ێ-n_�*��*�Vs���Ҝ�G��!�\���!�1׳|Y��I������i�*�ݔ�R,Z|�QA��2q���^z�0�FZ&fe���k����o|+>m,��'IX�ϑ�_>wc[]�8]e��ZE�!澀�V̋_k�P�E ��u� �4��cV���#�U�&SiҊѯ&v"��^g��)>�M
��y-�<c.�ˉ��r���R���-��g��������~��}Kj7�Bj׼��9���(3p�������x��$k�g���{2�OK��8U�T~��-@!�����v_��S#���Cm�N/��*��������|�h�w�h�3p��H�62�R�nO%��n/LS���^��0:£z�`������`��Zx@���r�@vT���!2�6aO�9��fE- �_�:��%�A���-�":���'���8�}�7H��7�y��Q�ϣ��M��0�?��ό�s���X�yvuЋ�a�)n�̱�:��N�+�l�ʭ7�ُ|��ʟ�C�x�]��B-C�f�+q�^�Y�8�s�.�N����g��#�,���tlru�A�X��U ��>���c<�xo�j����!��J��d|j���̊b��=;Ql�G8g8"� e�0^oo�H�4�gU�įk�Kj�f�ކ �^�6s�W/�ri��#�����=����3��~�Bm���djx��O�'�U��*�5��P�6waq�헅�ف�J��{��>C�P�n1^w��C~~��#�)5�WQ����ꨔm����W���@����C0�]��N�ĺ����j㞕5�+(s�*��UǊZ ,�X�w���,(��m��}~3�~�.]��R�7�z����f�Z6�K�:>2��MO��/Mg�{pI0F��ߐt@i��q�m��JˮI]5��kw�Qw��-`z�%�h�)�>u��K����W$��=�5��j+xH�qR淜0p$�J
��%���_�Z�&-F�(�������v��z�<z�����	|�=-�M��I5���G���f���z"R�G������K��✬}\��%p��C3�l��~H��m�Os�����5��ƨ0(}R�K�?ú%�s�J:z�&�ȤJ./\�k�a{�Ue	��]��UO,����1����G֮B�!V�R�)��Ϝ��\��O�J��/���h.�<�9C���J�é���ֿ��R�3��gDw��4,"����^�x�NiSG�F䊲o�݉t��A9����>��G�"��\*@@>[�,�L�?D��=������@r*�U�a^t� ��A��B.έ�ѐ���n�^-�c1c�������}�=���T�Ԕ�ڨ1ձ�`������7��Ca=�`:e��N	��~l�3V	F�*�#�eF����8,�r�����:�K;�,i+��nn���D�!^��.r��S���PhVm`��x����b���z�i6W�&3W�5�;:�#��Ҵ�%e<��X�n��q���3��*sU��R�Nqg�G����R.D�ua������z�������Q�ǅ�`�;��z֜i�-��*b��K�����H�.ks��:�c�b9#梔��9 ��K9�����&��L��{�J�n7-�����/AD�dTh'F�Pi�Б��?�Y���t/��Z�=��g���q�Mx��h�h�·"cʱ�	��P�;�<��+*O�F	-�̗xx�z���<Dg	��;�c�ζf98�\g<D�>��7\�a�$K�*��3�̐�9�Rk�:)�J>��L��!=o)��_���
�S��s8�)���O:����ir�l�k&��><L��� ]��a=Y��n�RV#������
ag��Z�X��7;���Jo�$���h��U�M�^�?��-FN2a���J�W�b�v`޲��#��ı�V��A�b]��
J��3Ti�!D�n�TV�W̢o�)�z�AN��a�e?r�0�Կ�Ȃ�Y���מn:s�B�9����\r'
�hh�S}�uDk.:�p� ��@R[A�	ܛ���|J�y\��Zx�iu��?3��������E��+^J�LO�M۟\��;�C��f\W��5Ҹx��D�Uc�Jթb��}h���(�T�F�
_��-��Ar68 h4e��?�?8���)<���a�}�����d6�j�X��r{^���(��j8�B�d�L�{�(���06G��Vǋ*\ǘE+7�:t�pm!��+:Q6<�/4����	g��"�c���6M|��z3a�~���%H����*P�:� h�V�_��A��PnD\u�M.U���)��pBÛ����b�w	�����h��Ďn>�Jo�����'V9�H�J.�Ԟ`�����⛒͝�i�?�h�T��4⼇z~�£9p�����(#����.���F�m�߂�ƃ[ٔ(va��\O�P�7���	~��N�wH��1y�#��Z׋�>�m%�c"��6�`�{�W ����5�B�7Ec�f��#`s'{�b�b�<�- B����W�OC����HmOg%qA3i�2(�	�3�H%G�Ҫ�q�W^c��u[H��Kͫs�+,�aD�z-�����q���ȏ������	��2G=J(b��o�&�]\4#�Gy�\��ypt�L�@�+����D��#��*� K��h�5<
�ϡ��ݒ����"�&�)$�e��d�em�J(k�A�4M!h~`���~�MJ3��/���+�wl@�*�q���]^R�اN��M�������vc����� >n붛�f���o?��.���������5��i������L�ߺ��`����]��@�v�x�rm�W�2�H!Vrx��Ӭ�ӡ�)$W�c���"�_H�n�Wx����k�h��9��<`�g���a>�^<.,�����5�5��<��aV}���$*�����T3`��DS�)4���m +�g�Q�R5�Ȋ�ݯ�ިiƈ�<e�����#5!�I�ݢ���b�\�����3�����ZS(1�o\�t�/�k�I�? ��J���U�B��B�Vrb��8tP<3��8��V�_ڸb.����䇣Ѳ������/���}dS,�zL.�\��\���X֨O�͇�0�/xq����L�r2H�Q� �o:�6�`a���L�(���mLb,�C��m�Ye�Lą(|�-����y�-����' ��☧y���.W)Zy�m�������1���W�d���o4��� �vX5�$�nEӪ���1	X���¬�L;�m���D���p�%h䆑'K�[{��>sm+���7���z��j R��_�!�
Bf0N��qC<\��C�K��?�+3�ԡr�$*p�eȇ�YP���:��Z�<Z�xb*.����.�y��;>��q(�	��e���u�����М?�{VS����w��8�8)�8S�p��i��v�Ck��[r��B��X�a�A�RbD�=t��ʧ["e�����~\�Fw$02�<a�Q&<TE�[�|d����uþ����g�SLy�x��C�M�-Q_Rԣ��T��]	i	�Xo�Ð)D�593��bH�A&�Z�#̏r�B��Vsԁ:SǛ�Å����_ڃ��K-�'��?����։sMFE����xZ:zKƌ�[�ޤ�By?�����e6�1�Pzbʌ���T�\Z┕e�L���#_�����ڛ�õ�/B������ʜPB�L��z�чa��]9��tv1�̅�Ck ���3Y��^<��z��L�.(UJ������{�an-n���[ip���8�������D���(�B[��|�5^�F�z{�l��A�/g �����KL��
�D �A�ͤO�;�K�O����$$Կ�.b��v�aǻՅ��>�������|���R[,	�p|P\>�)dz1{����KJ#��x�TOa<��a�0�����p��!�ē�t�����:����|f]�lMJ��u�k#V�TjS���&,��xL��^��U2�k�O��o�d��~���0�6W������e�"�r��
�� /��*z���z��z�k�\	��(R�����J	ܾz���c�Y����U�J�p�G��Z5��d�&w�����>�"��Ϳ��Q�|��ըހ���`˓g�c��]d��Y�ﻝŋ��Ix��ʼ��M�"ڧm,��s&\��~I���h�Y���7��" sЬ���S���$���M��$NN�<�F��kqa��j8$����\9�[��EL��k�"R�D��Rg��ߎ灇E����V��% j�Ls-��o��O�������� �����y^�H+0LK��i�1b݇_�8��D�~AD�,�V� y��/ć��d<��"�]�D�򤇲�%V+? ���[� T���H'uIF&���-H��a���YH��\�ld8u�Ag_�^�t�YI(�I��_-cgç�fXK�]V�M`-$�����K*/���֔Ag-�Yᲄ�d=����4����P�J��պ5���}�քPaW6�r̓��X���m>%_:ǊmÈ^"2�e��?A��a&�#��35 ��w�H齵f����p/�=zu�h\�`q�&Z|(k�^e��C�?%WJ�����9�Ԋկ���X��$d�̤�H��ѯ&t��h�����v-��@έ���:�ծM�7l�wK����;-ɰ	�k��V04��CJ@���_LV�`z*�bt��qۏe���dr[Ț�x�����~dEh��&of��Vecx���4�S<�HaD��`u�&���%����v*�jD�"�SCs�Q�J�砵{��_|k�{{�"eC�8f��Ȕ�D�� t�[]�Z�&�4�׬:�D�{X«x���$ه)��Iʹ�(~��:_�2j��v�N&q$�qCo�ӣ4�*09.�ـ->�	9�,	_��pƟEu�����!�=ڿ��/w�$���a�^��}���N�[]�A��nrج�J��{避Jmgk�f:}m�gO�~��zS[���
i?���-ֿ*AJ=���Q2!�XE9��Φ�;�a���
Ս&�n4����:��a�pN� T%��AQV>`hJRi�l�e�r��`nX�^��/��:~wn�@�]���w*8ҡ����7�x�?�{�T�Y�1��")���x���W� :<a�����Ϟm�t.U�
�2�=�,f���%M`Od�u�"c��1I�L���[7���]d���T����՛Ţ/�[�<|�*~��Ǉ���� RÏKc�a���m�Ԗjs�I�Ǻ�A��i��ƀ8s��Zw?_O�����ǖ��[&_��ǠM�(钌��R�^�]Y8D�޶I{_�Q�D���Ԟ������k����T�6h���L.Ql���(�U��<IJ`��� b�J<����$os����J)��ݾCt�PQ��J���Gj��rz�4���~��}����+$o�O�� ���]�9�����+���Ͽܨ��)w���Q��C��%���皻�N,�?r����<�Zw����Lڳ�n�̴i���</�lo+[ C���D�r��Y:?c�!�G;w������h	���N˺���L~�;��-�5�籱X2�	CJ��Ɵ�~TE�0��Vֱ*p0t�4�<~�C	�@u��#[rk�����S+��ܪn�����h$n��zx�eF��3�ԹX���Fe5 V��w�¸�tU�� �]����&~��`&IM�b�&��Jm�%PR��*��7�!C@?�/DƓ�6�'����ꞣ����?��>���푾�|x�yw���.C-k�l]���D���8z�	�a�:����d1@���@�|̷�͐�L�V
�g��٤��?���A)̯L�yܓ�
�ݞR7�#G3��S�m�8��^[U���[����� ��}�N�n�`���8��^g�m�Ě�6)�6m���DT�R�~��-�b��(q�v�#7��֏DuB�A�d��˺���4n �r-�tn���¾rĴ��?B�zEH6+���;��'a�8]�<dC��H�a2���#(6��084e~ʩ�U�kP�w/zI/�1��b�~c]0�qI%M��o�gaH��曄0)e�\�œ�]��g�#�������v�'���,(��;��v������>ľ��.���WOeK�I��W�#�U�9�8R��t�[�9xU�v��d�d*�1̔�ɴ�|]�}�L�i��t\�h[��Fa.slCrȇ�8V=T D�V���(>ȹȅ��6V��ܦ �0����c�[uVOyFx�#����wz�xJ%����u�I�}�W��h�z7�h�_p�-��4l�2�fC��Wƽs��2��MF�P�����,���4_�Qz��`$����ą�s��d��操_��I�4��8`�+;"⽖ݟM1�y�㳩��8��a�ҥ[0zm�:D�l�0�QAT���C�
NJQW��l�*���L�`V�A㝊yAͧ����Z��0���4������9���;L�A_^(�S��-����Ԧ]m\՘+�N��G�G�B+���4I���gP���>��G���3}��t�拼���C��
o#i%��;b�.0r�V*L����@L-6.�$+�9f^�.�Ζ3�P�ێ����}�磙$<�
��?A�fZb U�Aa���(,M!�d!	�t28t�{��q�4�|����A�e!�]J�]��c9I5�LY�<�,��n@֑�m$S��U&�?�;_e�n�]�gB
T������|����{��[#�#�ֵm>���A�y� |Iw�I�n�W"(�I���� d�P�k�T���H0=Q�����Q��4WX��;�g�l-�5�m�L���A�h#���(q����6�/.�D��#�5� �Ր��"~~<�jQ�z�9��ª��T�Ƅ'������3&w����w���e�'���v�l���l>��,|��g.�X��DͶ�nΞ��� J��u����}xP��z� +�㎗	/f+��20η� CǺH*�
��o����qQ��gi�.��3o[tq�O�7�;����� ��	�q)1>H��`���T�c�$U.�+��t��g�x��D.��.�U[�t�0�����@ �� DU�M&�SD�lT~b
8��K�V	���\��da?��ױ�}��!���>��EkK|l2�шy�RɁ)l�n0b֩��{�s���=Y���	~�ir�D:1'�T`�z��̒G'm�Rp�`�?aI��f]j;��O܉7s�]�S���=���eI%�ʒ�/qS]�8�A���r�c)SV��i�rjG�iu�'xxF?�Y�r�'0���%�v ���LOV��rԊ�^Cl���=�6r�U��b��'�~�r�4<"�ֲ����9��R@S  ��(/�����0��tL9�AI2�"���r�?$kn(� IK��ZJ�ꀟ�(��0ع:�2���"�\%���
trW��N�ّ���k�z���r7اu�S����֙C`9�c|�$�.^kVpIb����2a�W7�+_����]�y��\�i�ۨ�=J��]��*�7�ą�Kag��m�(�(�w��9�g:�{�h�]���Z.#.�D�`��x�R僯1` ����~�����D�t9:ENI��}�c���8dK誝��Pz�;|�S� +�k������,�@yU���mw%�XDí�Ob���D�(yN��E�:0��C��=�����R�SU�ɥ��y��U�b0(-�����-��п��+���Vk".IP$iUű4����:���V\O��c�'�sOs�&t���Kc�&ի��p��A+x6��N��[�k��ʂyƓ;�/����~����6R�-�=7�lp7�h��Q~rϾR-V2�c�A�a��M��tJ-%�hYou*�9�s0����p���\���hj�Dv�s�a�?�voMfĖJ4�����3I5!i$,I;�rT'L��L�m��C�3���4�\o)�	w~���5�v���g�w���{�Hv7���lGt<�R 6�7�£7Z,�!LG	#�iR-�t"�|����!��4�>Xt��(�u�q�p��BЏB�w۸k2�8��V�G�A�2U�pE��;�UÂxd��:tV��7�Ă���0�ȫ�ʨ������>�a��WDX܏���o�l��lt�y��.�Q��}ɖ��D�7��~�Vp}��~S�d~G�;�Rofd^���`�o�� �֒�h��Ly`>�81�ki��x/�m�u�8B��q=��g� /�B�4As[ 
ٽ^�L,����8�u����$���D�Y��Ҧˤx"R3��k��Ƙ�@��.�>�@���4�R�CsS�)��H�w>G��f����z��N\9���/���P(DQ�j����D,��2�:��@y�t�P�Wd�����ɴFr�9��"U:� ��U���ԇq�C�����p���b�����]K�ck�瑃��G��͎(������0#���AR��v̗*�h'v�Y��p>>���q4�QǇ�z�0��ٍp�J>�Y�21�����9ʔ�|[�οt-~AiC@����D�{����K�n�ǖ��m_i�����C�@�����G^O�7�2��U��9lF���������$�g���|�����6�|�nA}��@?ɨ�1֍GL̀T�+G&G5�|co��|�{ny�wq�=m��4�xN�v,����Srޗ&�%�HJs���U���'$�*�F"�y]���>��}w�!Xݽh3T6���p۵vh�`v�
�x�t��S1�3���n2ca�@��%�)-�IC�n��e��b��m��K;J�:gj��qqq�U��"���وR�͎� �y����4���Cj�!�v��&̺�AC�Y�㛗/-��'�:M���K��-�eNxl�w$�����Q�*!�f�ą����=G��'~�«޴;��T :�R~r�\ܡ�
�˄��� ��i��'��%�2�k�ӟ1[4[bi���䠎�/�C{n{E��v>7�U����"-����i�PDe���(|�c���lg������U��[Ǧ�v��<4Z���c��g��J$*qS�9�X���?Z���D�\s�\pf,m���M�7��k[����)v�"��>$w���Z�0�̧w^�n8Y�S�º����U;�����^B�<Y㪌_�T0`���V��u״�+�z[�O����E*�$حd\��-d�W�Pj.�U�7ǡ�}	�<�j�GO�������t�+Q+H5��./��D�!C����
�8�l�m}u��h�[Q�rE���H:�2S_5)����ͨ[�F�!.I�vbi�Ȅ��|��͓X1'`��bx����٫�N^��t7��c��{Z�ܜO�N>H��e��U�{gj8Pԩ��z�����������'NI��{�`43�㼣J��}�z�|z���?�.��Ӂw7ei���l�K����tC-�jySp� �6qq����3Şk�dŢėp�p� Ö��<�y���U����s��"IMۄB�d���m1�8�*�]�'�nD9����i�\�XV��Bx���:���k��?��r���ݳ�9No�mp q���X[Bץe5�5�U����ae��۲]cZ�\^0�8
�T��_�Sa}��7����D>:��0"��_���,�k�{���5�z)�	�8�R�I��!FR��V�	[�[�E<�ݙ&���{H�\'k�m���p��.���zw�ME&[���oVm�+ͫ_c�"_����>�cv�����{x��h��8��E1E6�h��{�f��o�b:�^W���7͑���M�{�-S
�����H'���"��ژeUI�_��IBS�zΒ�y�>�[���e�\�xmS;m��1��%��5�
���eʓ�1�_�H�:I1��~S#?����K�u]I7�2�����&I�	�~���∉e1u#w�К��c:�mY��C����Ҧ��.���N����.��<�������U��]̻�!�)<�bLH!"��ؐJg��#a�O��R��qK���_�f��d7ۤ��c�X���C�+�$�_V+�>=("���k��sشJ*��äߪ�ǌ��4x��sOl9���AG!���3�	\���ޝG��~΀Z}C�T���d'�3i*^��6~s��d���T)��I4��}���B�%�	e"����Bţ�S4��1r��#�%������n�hCC=^e�������1<��~��s�0L�L0��CRi���c�FM�����ăg�\��4m�l�.�$Rp�c��,�rĂ���^�Y�a�E��<A��Ks�q��aV9�I�>*n#;.�l�`�P-l�rWx�#�r��'�97��H��^"�ɥ!�\B����(P�Gf���w�(�����Fo�#ܠY�3���uk'�K	�sANL�O�͑�|�����DH�j�3�Y7EW�ϫ4%(&����X���)�¶��V�v.$�\S������œM�ws\P��v4:@Dݓ��X98�SUM��0EzTe��T��<���J���x[߂�d���)�9-
��m�k}f�r��Qr	Dz�pUAİ���y��T����
��ʠ����h '��?<����d�_UŹ'h~���I��U��Bx�.\{��#��S�r~P30��~�C<]�'>�X��(d[��#0��	�*1{��H��*o��}���4f�@�:~~qOU�� +�~^��{@�٘�k��Sc�9f:�S�����|�H��`"���*���&MN�n��oM:�=p:��*�A���/2�˾	Ef�7��AGجߪY�2���}�5�7��O",J��ə��V��c�8^���b�`��8xM=ѻ Y�W����f㝜��a�6$V�o�ȃHOe��?M�;>���2���<��O��O�eH፞�"" s%�QvY�"�+q.�.
���aY��z�fv�qj"�A��mƑ�/=���%��H�}c�������{%*G��6�K'�qUk#���"�[��9֞���[R��ӏ�3�v�&|ʧ��������牃M�Б/3��0x[J=�z�z���M���"����89�������S�A"#�k��!G�6��D7��S�{�0珇Fť�x�����d۸��zv�Sx�`8��x���!X�?<���Ns`�I�htI�|���'ADu�5S� �4R��D� ��
p��H�.�ϊO"�o����޺�hU��\�(N��&:"���!4R5͑P�/��?�o���8����=�����4�L�Ө��d��fr\��=��<$�<N4-��rՀ_��%�HO��;���:���u~P����q,�tS�[�%,�s﷣�!���\�S���;�?V�W9�p��V���,r�7��i~�?�rRr�l[Hj-��� ʑ�y,�C�|�=��	���㱎��*3ֻR�8Cg쏀j��n�T��ّ i��I^gR�j����td��3N�u�{R8���:�u�F��bp��so RZ8�4l{�np4`�S�I,S�\D�3�g���b4;8���x�}?�X�	��	յ�ӹ��)�g����|�z��n�'�����Wps���6(���Zg�4~>�:3uh;�j�ط�Oz,䥏d"O�E5�ۊ<*�g�:�xW�'��(�+���DG��+2��q���i�J$a����L�?��pGy�R�}^o�R���[^�47�����`� _:q��g5��S�ڬ�-�:"\zy�d		
��o���$W�����O�\�:�R���*�xqB�SD��5H�W�n�j`��z�e���}�P��'���Fc.�]�vA�V(���}�V<�����n8������J�rz���D
V�n���_���=����R�7]����ٵ����s�%P�u�$G�/\Rq�a�W۳G|�	��}���y1�h��]���t��t2�G|w�GQ����d�=�'�խ$�r��j�X2�O�?v,�݃�%�/H_���啘�ȇ�X���n;��P��An��9$���q��2�3�H�z"�w�K���q�Ț��>'�?�� ��KJ���h䖬��M|랈�X�czbz�����߽��u������σ��c0�������b�1�1��:�~�m�����(RI��n��瓔S7��ɐ�'�Ca!���[��\p��M�)�	C���̑p˧J���j"����Qۥ�֮$	J��tbO����y�C8�je��<��;��
Cn�LS�� @�Dq��y�k���j��@��cu���2��ly�1���˷�/5�lI*>J=�oЦ�g��N���VJ^ؑ�<P�>�%��Sm����1�j28	V5L�e>>�s�C�˃��ARF4ĩ:��I5��L[\ܙ�	����j�3.r�7�[��F�}&2�k�wp����H0�gLq;?!!�B8=�.�I�+"p;��`;����j�������I҉2�~3�^ �g��R#g����ng`��F%�\��洔q�k^
���s�h�D@����XP��gs!=Q?~�jqUЇˎ�l�s�^�����6D(�C�v5���s��ﻒ���� ���{לm
#7� �������h���|���O�KP�D!2�Ll ã)t>��U!��}:S�.gl�8�ju���*�zG��b��0���x��I�x�k~���<U�'m�2
�/����0�^A��@��p��]|�n���0�u\x��STR��u�qca��{'s3>.������^�a @�k��2�W՜'\s�ĵ��-�:~IvX2���Y1j0R����s6o)I�H�<V��5�`(��a1�}ߪ����Y���5���W���kK�P��l�7?����?�q��E*�=�;�������|]��4�YxUF?�3��kRk~���8�ӻ@E;�,"5;�ܴ�	P� jj���/�aA6�%�O-����0nh" �ί8U�VhR�k�t�ܼR����ɢ^ȿ���u��7@f��Dk"[���Q����(��ȷ"��U��T��B
��/�uZ̤U���7&���ӵ��_����A��ng)}�n'��P�i�L�1H�����C��ߙ�C����D�G��P0��F�w��D.�w����Őz��'Z�^ �ס"��ݣd7�9-,P@��Y��Gx�U=�T��'*�U�]�Mm(/,�&� �]29Q|��<�o��O�C���V�>�,��EhR�C�~B�H춭��p����C��7�����`��0�/Z�� �����*���a1O��TRE�{���������\|R�`_�u�$��dXX�r�����wx&$m/�����T�=����Q8����S��/�y�C�R����uk��fp�e�e�f!�ߦpm+Q[�7Z6���7�<���e�,|u�ۍh��MxD���g9n��!)����t��d(��r��]�����H>ΫWU^Uq;R ��U�E{@�R������&Y1	�?Q�i?o�g��P�i2���O�{�fФf�=V�K=5ao���I��%��1�L��[hJ#	���4�@�����G�
  �ȱpb�� �� ��E�'�엢��fǸ���?YިL˯b�2i/��t���w��.��1��;�e�Ɨ`�P;�+�]~76J�Z���~�
�?�u���QKY�S��A;�f�<��܌P��O�A=��=:��)i��=��� ������$I����E��D{����/Gҝb����&b�4CJ�ʍ�h���e��g&�y��5%?K��zb��ͺ �Ď�qǐYM��w�M��5"	��0���8��_��e z�ʻ�Q�KӶ�~qX�j�O�'\h-e0�0N\�!���A�|��j��� �;�;y6����/?�K��=�SF���z������3�L0ey*UԒn�s�:z �q��5� ��B�-�"����)_���w6��җ��c�?�KE�}{V.�z��e� ��K�c?q#���u�G�K��3"�ZmO�a��WGL���5 t�&O����&rP*1�|�+��U��g�Q�g�,�#�~{�'�&א�w*F�J@K�b#Qo�܋����u�6z�B�x��6�OG��_��f��n f���_���Y�p�Z"~$!�	��9k5K��T�А����&��.Ox�c�� �FX)�;AhJ����Vb�w���
-r�������P�ҷ�)h���ܫ���u&0�ZɌ�"�H��$Nύ"ŊZLƯ���a���R�D�1����n����ʀi��n~yN�_�'Q��ZawU���4F��:C&�)�E��R<��u�j��9�k��m=oi���ݐ�Ǝ�����S�h�]�	�P�=����\�F��R0�/�l�oF�`}�*io KJʰy�_n�=��av��cۥ�Ov�����ʒ���������25d,�id�S��PU~��CZ�Ɍ�1�&E��%W�GUL��W�/�����NS\T�*�hĀ|��7��WN�!�����Ǆa���������S~�әX���nx��@j�!E����#!�*�����-e�`>P/��4mշ���s0K�^ͳ��2��rBS�����b?��Yk�
�W]���#�񫩋 ���A�u���@\~.Rklj�(�qh�u�±U��w i�CL�v?ܵk)�� zv9�*M)����ME��^sF��t��f�,�|��H��T�ٱ�A�d`\���.����sU3mKXB�<�҈E�ZV��GK��A�\"Z��FqA��u�����/d��s����:��f�r���H?��Y$�ͱS��F|!�l���FM�9�@�=��5nCC���·2!eMbT�����ɛuf{��<�_��)\+�42� ^;J��>��OmN��"z͑N�@zY��-l�����_][j��Afq��a����g���*;:�d�6�0A�ۨqR�|�k����s������zY���̃���7w��
	G��4L�*�����U���F�A� ]��9b�I��cޅ=��!���8�� �Ev�좷Q��%]Oq�O�%�t�O�<2�LM�p����̒�a��
9���z�!f%�����WX�w=A{���:gS%O�`}Q8ף^����C�{r�M����\K�ЍQ2�!E�}�}9j���%i�)OJ��M[�4��" ���Y���ds�ߍ��l$>��Ű&���f�d<�Qo
�2
��n� �)>�9��9!�Ë6��ؗ�ᅺw��yH�Ay k��F)k�n�6̢�3�^�<�r����R{�!�	����Oh�r� ���Vx��Q�E�
(�+�MN��3P ��i�H��m,R|��w���Ii�ej��!�Jy7����y��Ed�Q����B��%�<�)Z3��`��4��|dVR�o94]���4p^a��>��`���gU��2�e�/���|���$pb��f(^�a�]c�d��	ڈ��Xw(�JMx�H�E����F�J�|o�M�,��︨>m*�n=m=_ ��<����������Z��N�����n�ʳ�͉��)>��-՟�������x�K�T���0]�E���=��,�����8`��>1��� ^�{����-�;l^(�-��1��������M-;b1�.���m�}�˗�%�"�k:��V'�=�; +aĚ1	zA=6d����Kc�z�ԑ�]c��/L=�f��~�>���O���9�"�1Ҵ�kU�$-E��'��詳9�j-i��b=݆�ئ�_�3��Q=����w��~�����L��󤥈����Rn�:�zh?R��K���ݒ���d������A���DOe=T{�BqK�	�oJ�kA��= �H�M�PNї�� h ��\���|`�6�G�$�f���&��v��N$�E�����ד�u�ڒ�-��bdf�m��Ѥ0�������w�% +���
D; tw�=��9~s'�b[>�q��
�N
`��TWڱ#��k�"3)kϥ���D�� r�^V{�UA���M���_D��[�3 A��Eng�p�G���n4�x��×��yp������Lil���ެ
 ���6�5�->��Ar�1�H�����:������p3��v#���4k��H�+�M�Y�$�3v�s��>+e4h����%�;�Շ�d/hYJ�$ʮ������xY`����k�g�V�kc�w��m�̻�XGj�f��tBr'��V��&����'��/�~�ȕ�G#Z�.
Qe� :�{�?���1A�#�]���)93l�.���$eF���鈡��P�iI!!W��|���ry:��� �Fr�����Q�ht�&��'�?�6T�s_�{��r��r�{p(as���x�)�C�[�"���P��;��	~D���0Z�td_�2�o��t�Y�w�T��ujV<�ƀy�J������#��>%7�49��a����W����ې�wG��0_N�vyH�����%�@ص��8��u�2B Yf�3����Nst�j�6	�	�FkB�<��SWR��$�7��Z�n1�z��tQO�2,�X�k?[�SCF�U�e}�.M��I��� ��I�� ǽ�ɌH�W�ַmm�~���.�z�m^k��]h��>*���X�>|B,�ܥy4;��/j�M��C�Z����=c�?e�hH�Đ �o��z#�TS3Sg�\�+��b��3�]X�?�<��P%�U�������y]�x�^8R�n�h��H�?�QVh�i|�=+�QN�y�b��}tg�V8��-9�E`o�� ML���MHE<�U䞮�v̛��E�Yb]o
�qS���=Io��񦚥.�Qtt����oK���h3���?�?�#�=2��S͠C�� ߽���������4�c:� �qG�z?�g�3�<��s'j�!��`��v �'l<�DG�(هѿ��Y�?k�Y��e�L�Ĳ�:Di����k�e͸�)*-b�W-~0��9.�F�����}kݵf�ؕ��)�����Gw���pJI����%<����ߏ�.'�B!�
�#ϙ�4�.0���(Ϳ�wWJ�<��}Ql�R3��0���Zl��w�a�������0�hf����VO\;b0�˧�RT~M	�����k�.����`����a�auWR�BW�xB�!~��N��!c�F����aN;`���m�X��S��.D�_��K�����O��J��@����e�4���U�p����,%r!���p��<�5�F�~���ب�L^���Q���~� n&HgRs~�� ?�9�2�ć���_g���˯]����s{76���Gu�����j���;P��a��G�Y����·�g����O�F'[�sN���EQ`���:��#Q���|�Cb>��-Њ��W���e��2����U�C�,�g��6Q���$��x���d�Y`�4�����q�b�/�}�4E�^{AΨ�O����j�c���=�8
P��A������&?LEx�cH5nчz1-6}�!�
�&7O�Y�r�N���"ɯ���-u�2���%�z����'�Zz��)�Fȳ<��P.m�p��R1����+@���ix��G֜�f��3�l�q�s}{�n{�L�e�R�+D�d}&4Ӛ�"�(�1Ktú�o܇l�P�i"S�f//��mwK�5�ٟ��>�Z����m���腭�y�nv�mj	=���:��X�."v�0����/����ҳG����5f����|��f��� gލ���캗�TR�^_f<��q���Iz��Z�2l.n)䟇�a�k���g�� �qj㺍��� �?-�c9$��5�@��2A��r���ߒ��T)�Ϣ�����c�	�lc�U	N|T�K[m	�%�\1�a��������:;�`�~\��/���Z�������H]tMw��P��kY�M5��8Vu�T�Dm`|&hsZ"�}���)���yu9n>1x/u�GӅ�6M�(2���r
CΦ�_�p��& 숒:����&����/�&�H!`U:�XJ�p���5�|�&�j$؟���1�AyiSr�!�k~�Io��^Ѵ�Wkb�Ã�1+<���>�j��FM����`r��ѷΚ +��5sZU�vjf��r��>�5`���d����6w�_���!j�Ը�1��yKϳ��Q��gZ�d�G�Q9�4-�T�D�!���*
�< �[�5H�uM7y�O	Զ��1��3�PS�Wm�"��N��ye+5��3�"�L�Af#��/~�S��r�V�/�÷J�Q}܋��}���{<�B�켹S��kA7.�W����7;vq�x��.��@�!�	���ɢk�ڳ���J�;�е!0�/u&1 E�O���[���z��f�.�!���卐�&WϦ���t��#� ��=��j;�cy1�$(tNb��~��T��v gp:S&_>�T@��}><o�V﬽Ve]��ُ�: �ܥ1��[�D
�`=�nb���!�w��UH�J�x����Kc��k�Λ��j�oO+��4���x-��I�a`6�.6�u�c�4ۗ=s��Mi�2\`��YHU#�"B��V[Ei��ǋdV4�|��%팙��#Aw6���s��αqa����V��Ɩ6���铜�.���3��t�Q+JC>`�A�<��e�1m���ć3Ǌ>��d�*eɵb�����$�)O�G���Bi��RFi:�	��Y�c]D�׎ȿ뭧��l.]UfRE��@����s����O`L�![�Οr�h�O���C,�z������@�k�{Ϡ`���:��]9����U!f�&N�w��P�+i�dcM	�s2�P�Vj���k�o��[t��OdX���%��4�*�1�at��O�x8T�����K�v=�f����$O@{�;#����-P��+5�Hy����ݰ��y���C���a�Ym�4�"�/Y�����8����Rc �ڿ��u�k8�Sp�%`�)>����rʲ�J��c��Sxt��\�rwy�nn���"+���OL�M.@��`���l�!�2|�[�&���4Q.����񶍵�j��Y�%����$��{:0��ٻ1��Ƒd��a��̇+y�a1�����&�W�y��R'��m�P�������gcU���-���#��2(��w�������<�8�d�N�S6�{N�P��P%�u���H#1���5*��W����t��w+�@]���R/A�����oH� ��y��\����D|�IVUT&�uJ�M�Qlwi	�&̲9-�J3-}�]^� z�X�-4����Vn�T´��4�7��=y��z+�]�'�vr�
Ll@�d�g�Q�k!*ڞ�f�޺R�%�EiZ�������P�M���<s�7�A��?4=-2�����6N��H�R��A�ZF}���5��Q�:GD�
+Q�O��wu�d�D��RN
��	�M�>m|�zx�h�����	�������:��@�����LQr�7��^���;(�XO��+5����oY(N-zٹ��S��7���x��m�!��q���ʳǕ7VX�l��ﯓ����`�z��+���՜"����gE�L᝟
�>=�$�3�n�	P����%�^�c�ZN�����O$���M~ N������g�M�p1��P�L�#U����h:y�s�߲�~C��UNL��|_Z���X�{.�o6�����x�>4o��+���m�B4����� j��s)C�'�����L �ff�f>�v�P�:�v�����+(��H���#fM��Tj��"J�C[T�߇��Um���1�d�|���͠iG��_�����G5ڊ�'5���
�4"#��ԭV�Pb|�������25��+=��)��m&��A��X��.\E�ZK��"]2�ǵ�Fj�!uE����bY��D/�{��<|���P$��c�y��%�=TwC����iۂ���;�0I�C�����������������q9'q�!\_HY�U9�B9��D��'�;�*��6�#�N��h�>��|2s$��
d���e$MȦ������W!��'}��;h+t#�V�2�K����|;*u�娘|=7��`Y�Ed�/QѬZFz�U��ԓ,�\P�Pаƫ��뺧6�����LEO/�.�.R���0�:�U�Gu�h_�?��*�o���-�9��I#��BfNi��\[7�󬥨��=f*9��jeiE��G\���XX�Ն�=�Ŝ��A��
.#N�ۍxW�(�V�G�F��� Y�{��n���0_�ℵ}�aW��1V��b�<��lμ�e���\��<��BUK�O�pFZ��~�G����b�" �f~��}������b=bbGQ��h��3
f��!��>!�gtR�!�����NzQ
K-�������ڋm��CS-{u����G9�įg��f��%��)�=%���ݾ��l� ?��R�O9����	>���Ã�Ufb-��V��Izf.��O��(`���I���Dץ�I�H���/*U?J�Ǉ�N���on���n��td���Dʪ̷�4)��]I��O]���#�F��AM���]�/�3]��,+Ӛ�uASD��P7���*�hәXf�I�������A/R����|[��Ha&�� �J��sq�n\�ڈ��"�]3 �2��� ��*�������d9��nO��
2���p����>[78w��sv!`��w����[�-�Qm�2�T��0�6b�E[2q�i��p(oso�kﾗ8�uy���'b*$�	$	�\�O��A��\ރ�f��*���
��M�Bq��/�r�O�,��]u���
�]3q���Uʷ�N=1��}��5��rǍ��_$1k	��|�u��
^c���_�\���Bj��w���ZX���+#�KJ��x�<k*m�uē�!�O�	�~j���r�ga��O!ǖxҋ��Z��"��SJ�vJ���ǧ�=p(3��|I/(*u�Ƣ�I����J^�k_Kz@�����R32���GF����Y�3=�Q5�k��[�r��NT�yq��h����P�+�KK��cl�Z~eٱ|��y�L6ݸ�
�A�Z�]�!�z��z��@r�d۔�Nlf��z
n�"�AD�iE�JԦ��ZH>༚��O������[����(�vԒ�I�Z�����MѠ��_L����@�K����|�=��S5>��ؗ`!t�`����[���[�A�m�ov�ag\�=u�s��R*�X#�hx�2�ɮԔ��ȅSa���Rt���Px�/C��7t��fy�Vw fȉ��.�M=hnƇ����'��fU4�Sȏ�>�o�K�N�K��XYĔJ�s�R�s%��m9f���<�,b�L��U>x�E� WGR��|�E��T���4��@<a�l���q�������aّ#��fwI�=��w�^� �y��l�)B�������V˲O�j��9=�C�Be��j����.q����%�G�1�m�@�b����R��i��I����������Aq������'�l��y�Q<9���ؿ#��-����8c�,P_$��*G�+�fR������y���ݱs<�|nJ7ee�t҂ n����+�����v�&�m���v�/���3�9A�jy�������5}"�x﵁����l\/��=>�H��s�w+}������L3I�/|\�����e0[����yz�0��d�?���[��H8dJiD"��Ք �Or��o�<ޏ�f��F�a:�n�6?��@xq4�y��w�f,BA��ۤ(r0��*u�V�$�wJ���k��o���R��kT��-���b>ǎ1����r?����BaY�Ŗ��m�ѯ�?��s}<�^��B]�|��X�����k:�r'�M���W-�*�:�:�˸�&倠�4���_�K�S�@V����5|�ING~�2%�H� Rڔ��|��
~��?�hdTt�4MFeA�9u�$�t�UmW���i���Eq��>�ʎ��{.�Ӥ�]�{�D�9T{�IװH��-�,3Ç��ђ��������j����G�iQt=�*Ii�i�&i�;z���"|�<�>��F���O�j��\���*��wu�ҥ&�X�Ȉ�k���(���*���;l�[lT�g�J�3���m��A�e��^�n�����	�~^:Vp������l�����>+�?����h�4c�U���I ]��[#eLI�HI�2+&q��M��p�
����>��+C+��߈u�҂�uR���|EV=�L�����A��ճA��~
�|iJ�p ��K威�O��=1{2��C���So���Йm���`�X�]f7d"-��o��t}�*S9?pVWU�>�T��Z5��uHP�nj]ęЖ�����͜�i?������c�¢疹��MSV|u�l�����S��cj��ۓ4��\�䢗{L��V�Oɚ

��e��P�i*c��/u�e���a�Q�0�ϓ��Q�t�[�q."�"���V㝕QSM������l�V�����Բ 8n�rt�oȾE��K*z
��B�9�qݽ����^�1`�rm>ܥC�e�]�9hKg�`'���c�XG��g��v��sv�CY�����x
Z�F"�1a�u�K��#-�b�mT 7���iJm���|a5C8��3��^��z�^��V
@cb�Q�����Wd�SҼ�ãd�N�B�/�|h�bh�r�[ߔ��㒛��N�	�2�n*	��B�`�ڠ��F^��r�#������	���;�����C���/M��ޙ� 7,Q��Ug�ET�g�S��I����1��!:��EƘ�������;��Fk�;f�a���nlp�NY���7\�#���v�B���0 �����iI�Q?hXv�����R������铘�A^��� �d�w[�&V�����a �:	������RI+����:��O��Ҕ�������袠��M��8V��Lf�pP�][+�G���fkZS�|�_4�	2�����i\c
��I�;;7��;_w�6�V�r�}ux�/ĒQ���Ł���j�k�,�[E7^����EBY��Y
�gK���[�|Yds�P��)�fx�� �!4��a��!�Ⴢ��-�	$ٽ!��Y���_����DZ�i�rk����o}���c�=y�la��qθ��3Bp'���c�!>���}�H��L��,�~vw���b��D23�~Bz:����8��� �^���<���G,(G�3C)ƽ�%Pe&���\�>��\?�R&�Z�8��q�65��]L�,nenS��h.��oD�YC"��p�+Ѧ����^P1�NY���]���R
�\������hB��M˩N���#{�������q+1�XUc�J� ��?�S�����(�e����$�wQy�4L_Q��C� �`#߂�i�T'-	YC��m��i�j�ދa٩�2e���okp��R����k�F�E)�愻Y�Aߠy4��E�c]>ϵj���^R�:Τ~c\�L0�5�5����I7��a B�h�O2LTV�C1,̹"���]�� �]X|�m~�#4�,�*K���4sM=v�;�/��nt�@� �cќ���?�ɘ3S��1�M����Z;ɂZ���q�2 "���V(�Lj���huc�IRtt���`��c�s�S�Y����0r@G��R�����b��:������^\��:U���kvz���Q�w37���+��m��a���:®��u�1	�(r�m'�2`75����@��)�����Ǧ{�����C�)b�r�)�+�ɺ�0SЬ���3�/Z��,�)�q��i�6OH|â����J�u�U���}����������)���>�%���@82���Yc3ʿ��Q$@�V#Y��Muq��38��ͅ��)�Sy��V[�w���J ��2�Q+�8�����)��.����set��L��Ѫ���3N�D�e�=�@_|c �V� g�	�6.@5o=\\Ĩ$d�l(�-FI;N?e���P.��*jM|�Q�����M�Mˣ5�3��9+�y0ϻ
�.��C��i fq���cA*�W�n�0�պ`�:tw8u�r��+�^�l�cs)��vA��9B=cqz�ʵ���rcDo6U>��=H��'�����.T��\a�m9� ��M��І�������Q�0�!��a�S��M�����x V�?�H\9�m�������4描��X.�-w_S&-�*�ݍ�`�-��=#]�5�Y��C;J*?��n��,3	4 ��;.�Vc׷���#��Gh�!��/t��um���\����7ru%:Jص[c��������Or�N�B���ڙ�K�F+�a<��ѱ ��⮎��N����]b��Q�׬�ȤQM��S��e��؇�@ܡEտ����NʲC�QIZtK�x��շ&�n�c~�/�6̡��|�@�1���3�k�E
���K�e�1,�N\l"���f���a��c���f�P�7|�s��*bpE��3�������!�.�d4*xAu�Ubx��)�6�8w1�x������NsF	�?l`kд���_�f�*_Lp
��)��`��8��EAWQ�6+xrg��v�}�nu�,7b�E�L^�I�'�wC��|��RCWa��sQմq�s"��9��H��lKOf)_M��Z$�MkS�0��^t׆α���Y��>kh������Ќ�1YU6e?��07bU�=�R/�6Q�մ1y�3� ?4��1��2�y?I�!פ�%�@��ig�~w�<^[ �N��U���P]I����[[�>Ah#�A��4	(��8�����H>����P�J����Q�j��J(=(����*e��D��r��n�1��^�b孙��y��~�P�è0�h&
��a�!�)��)�F8�e�ݭ�qr���e�'M$L�' ��(xqK���2ަ�n�f@�8z��ʓiB�ĕ����x��ч��3I:��tZ��$�}�T�}Y�dж���gitOa�������H�ݬ�((��P���s�&Gq���(?�Ȓ^�3���O[.?@��'H�7`�9[� ��dq�n����a��+ڼ�?�E0��z�Ri�`g�Pc�����P	)j�SA���E�A��:'�]��1�Π�4��U�Z9$�5ʐݙm���s�V'���gUR.(�S���5g��.��V!J;bxɌU+�,.܎� y�g�t�LW;�f#¶r�5!,�Y�<A�O+�\v=ޤ�\r	�.�d���ǫ#��3��پ�@�u�#.:�D!L[�����s~_]a��|w�<���FG�u�#5�5�d�\kQ�e|t蕇�b�^�f%lsO�.�v=x���tuEB!~�o>(�q
��>y�^��D8�*���hQ��π`�-%�����'za���3a9�8�V}� �vxd��8�WRKJ3u����|l���8<�_����46�±nI�g��#�6K���T�Ʀ�����j'��	 �p8?�v@(ҭ��$r���'����-��~��g��`�Ǚ�gx%2��9%̟�$UA�MS��D�Hׂ��-%��ě%I�Ө��QA�tL6��c'X�����x��=A���"a%�T|/��Yg��v�7.B$���I�������S5�Z�*�.�_�ڈ�yB���p[E�l��x�fqSE��عF)�̛4��;��3�� �6�.uTsaN�[�[�=�� ���'t62�{]W)l�u^;����7pǕ&�7���RP�c�KJb�SM��g$t�z�Pǚ7
f>�"N�^{�C���U0�(���i�d�v�����N��g܃}�� W�u�ŗ�
{x2�׺uO����2�0���ش>e���1���]jL�f==�]�b�Q�_j��O��O�O�d���R�Ta��Uѝv���p4q:i �sQ�B~�C��YVm�t�:�r�K�na�z��]����z�z��YG?�������!��y��9G1 �3!�܈R��ͶKur�.�� ^�����T��޸_\nq��������=Gv�6�+VlR��y���APy^:5 kr�T�Y��٘j��.N3��2���8�8Fq�mY����f��������"ͫx?Ͷ���E$L�{/ŃƏ���g�g��R�V�"h�I�X/>~>NK±D˥������%o��ޠ�(�ę��������UkG���󤓌�,�d^�q��G��6��;�8���UJ��>,?�O^�
��4�$sB���9yr
%�����|��(�PA���33��\�
�T�hP/~�\�l�q�!U>����K��ig;,�S�������Z��|�[��P�3�ܴF�g5�߼�7�
�#�ca����1~�"���h�[ԅ�I�$��6R��)!�!K��x�7/�u��"�6P�	r�ة��pRu
���Ǌ��]���=\cF�+����+��P���`8��ux.����5{44����ZH:�����3��}ǈ�a��-ǲq�mKb�'�XeC�!�qg����}�L<�v�(�D~%Q����}��K��g���M�49h���;�h�B|ĝ� �Ȏ����y�y�~�������D��ױ��K��+�oi_�vF�*H?��yB�t"�VG��u�5�&��v	�M�M��=��9w^l�JRh@g�,e�"j+}N��� s�������|(xA%�o�dZo�r���D=&x�M�V�}�8���I�S��"�;�	�{�d�E
�l�A�9�n�*���)P�.����������)%Y�"̓�������c��<YO#_�8�{IQ4���ù[��Q=*��hN�3ΟY������>�- ��J���®�g��\'�
��ց��o�K)���G� ���*���w�����|�ѿ=�n�V����F��?p�Ba��*��~j��q��n���.����^*�O�rך�v��_cA6�%�X@}���v�$�f�W����u�:������e���:����`��<�\��Y�:�.9Y��a�,i$�a1�\�	 D8Vh�h}L^Y��S-t�|0@'s�_����x�.`­Hy�� ���i�P!���m�&�dSV�ޚ� �k�;�ka���u��	���T�~�Ҿս�L*�0��H;�%]��"*2̺oL�uA9��v�m��&��r�/c��iS 6t��u4_�B�k��nsd/��X4X��w	�Q���d`���j�mc��4Pÿ�cL��U��\�� �;�,���=�sB[�j��6�?:k!���{S*L��|����F�u ~���e�Q6�6�½�}υcG�qeCc���﬜�O@����&:�U7�tZyKGl婈�#h�}vJ9��E�h�x��=�JT0>\v�Ip�M6-�+�1$PY�6�r�p�����AJ ��]T��sh��@��'�#8!����Av��*����Yi`��	�@}*��:�]o��i$�ev")<��y��ҙ�pa�=?���!7M`�m�/G�غBߦW!ik֪�j���՟��m�� ��x��h�4E~�5��Tʏ��-a오�7,W��q"�?4[9D�r4�-�͢�wB���#c�I@\������0�6� m��k2�n��TrJ��$eB�xc[/W@��!T;T����y0%7ˡ"�_8�Qg�ё�DG˩^T��˗�L�4�]���c�:O���� �������!Z�@.���'���4��lq�%����8�YE�=�W#8�V���^K M��Y���7H{Ю�+�L�Nbo�U8����xk;*鉹v4��IPۙ�D���w��(wؿxE5�ր7��.�"���wa{) 0�>�^@�f�^��U���HVB�O��⟔h�T��[�e$���S�xo�v�9�o����r�NX�ۺ���nX}j�G��q��u�ѨϠ�\�G�c\��+9�Bc�&��i^S[�[��g?`o��u��x
����2ȃKq۟��;����^�,.�D/��ڂ*:h���N��{���0�o�Jq���e�R�/�\ާ�����$i�h�����EL�k���"�L�gNr_|��C,�W5�X���մ~�����n�]F6�4{�Q#������B>JQw��W�w �����H+ u�Ӝ&;��H�������I;�h��D�w^�;�K�!s�]
����y귣)2o��`��c���N���!�M9OD��ձ;I�ּ�.9������_��%��0���am���"Gs������׹Rz��O?�Xi���:�h"����S|z�,Z��j4A}_�ou.�4~F�Q^T�Ϙ{#��g��m�����������u�=(��{O{I��lm�O��d}i�e0�������%$���o�#)����J��ͽ���>�j��"�̆���D��0��Agˊ#ɛ�4��	bl[��C<���֒엃�!y',�97)=����Q��/�܂=�7�ɜ�D��K��9�2���{�@��F�qR�ح�0E ��v��׾����aά���	�I�� � �.�DCu���+�����`�JVa�z� 5`��� d��L��A+�o11:W��>��L��O���R����ǈ���P�3[��מ��v��\�&�p��-.eӬ6�Z �|4l�y�9�hb߷���ؔ	��sBgO%�l�P�A��C�m
��Yi��#�4^�cO\Gjf����=FtQ�7�zzг!d9��
���� �}��_�Mџ�;�V<u�Z6^����&�1���k�l��t��ֱRD�Y͎�S��;�����3��Zb��G9�V�����1nL/������i�71-	����&�E ���L��������N�3\����Y�$�G�IsG%��&MZ�t�8)T��������08oM���Z�%�?,¨k�*��A҈��"�� %?I��EZ�
�{�z��q�$Uf`���V<v:ڞp�8�P�t�ôT�0E�/�%gW���$9�{�&\� ��Sh��V����7��J������K�EL��̞�(�r3�::XO�V@�n&ו�&aƿ�)#dyp�ݷ��^��;��8Z(D���`U5=�ZOVE&�jl6Rfh�.�EO褿ň�E3��;� =z��i���U�q����1�����U �8�ꔠH.Rŷ��`7#0�q�;~NB�˭Kwf��P?9��D�IO� �b�(�c	�T�<�u��9���ٻ���x,S�ij��	~�I�S�0|T���i�Z����L�OT-K��m��1�l9��$�'��{ !�+��I��t�_G9&c^����..!���̿:�*>�q���ETS�闀��V����E���zDNF�����?2�"ߎ���l�ݚ��(��_�����6�B�ޘ��G�е����!���&P�p�r��ϑ�=$E�
�b�x)�;�@�wU�`nyn�&����,�I�Sn��w�ZV�TM\|[�CհKH�(5f$E���G��KPUb*HN�s�)����t,��F�Xcyb�q����^�HX�uUn�=ul.< ��I���v�@s��Qz��ך��M'1�@���g��
5H�V@��Qb�x*����)����E��<x	M%�C7+�A%�Ӄ�����c0��Z�GL�~���(��2�9?^��<�K�ȍAԹ���*�j�o�H������w��s!x�������.�~ ��`�Z��ĉ�b�s3�ĭ��.����\�0(�������'8��HB䞎Gs�L��0O�4����b��09�{Q=)�[~�����y�c��:ng~x��C���k�B(�j��*I��|�`p�����z��u��b�T��wW dD���3P���A'����g�k փ��X����zk�+u%k��.������rl1������ɟ�����}Bd�����j�j9H��>�	;%y���U��:+x�7��1�c��n�"���G�ur0�f�tj��b�Z�.�O�k�v5e��%�2��]u�U�B��)��VM�-�I�Dݗ�i�
O�`8�:%�,޿F��p���?n2s\ �o4�ċ�����X���3��H}G�`@�;�g��b��]�d�[(G	g�`�Se�~\�����u�*s+�ҧ�QaId��v�HvT�(g�bP�(`"	us����&��^��ۮ��X��Cx ߊ3�hSidj�<�؀���E3&��B%]�ж+u<�*���^X�I �����8x8��^��K�3��(�#�Vٽ����Jr�W@G���@0�b�F	;���g4_�J�'���\2B%�k`���j��4d�{	�d��$�8q da����||��s���������0V�,��e���k�e4v��9:�Er��}#|A۲2�u��	�9:�T}�P�&�?�U��G�._��� �߷�t�1���[��]a�t�kt�v
ij�G$��V�B΄�*[��ߪ�f �H��b��@��Ԧ1rܹ���S��uX�u:Q�.@'~�'�	@qG������� [�}"��?2ҕ���!Ǥ��'�xߓ}�#5�ejD��v��ښ-�f���ԾS���Hxq���{+m�sO�AzdB�D3 ��և���Z~1k�bwq��TJT��H�a� ����do�8�TSux��A^�c�]jT����^�X|���� ��%�M�Zlى�%:\��L��&6�<#oB�֝��LT+$;���2Al�ˇ���M%����d2f�N�NsacJ�2v�y��4�4ђ��أ�%�A�9=k���k@y+���gf8�����:�.�����[^�}Ɇ��v�y��H�*�B�z(%�Cм�`��x��Ln�h�< 5�%
����S�#t��P�o��|T�-4:@T-@�$M�A{���L�t�Ŏcڽ�m��7t`q��/wT���T���(*zي��J7
ة�0�#�*6O.���3�y�6�ڣHB q
w���2a�)���d��!�y���uH�� ̙�E��hC}�Kn�w<�_�U���mL�|��K3�pIN񡗙�;�����j�LP� ��'����֕��[�G��/���)F �C?	k1��J	ˈI��ԛ���θޒ׈+�	f��d�;�O��H�H!����$e���wm��nuI�]��9�H	3L�$b>�O�@��b6��2Qc��-n�r���R���`'B³|�'Og�3��?�+����~�W���ˌ��#8^#]nF5��7��������i�c�Y�D~��sv�L`�YL��J�����^9!v�2��8E��mA��~�:M�mx]��[WյxR�'���w$�����۰���@��i�6�ǰ��w�ȰB����R��D���(�yn��Ӭ�O��\nX1������������4�E����J�:�%o��'ۤ�+�t��4�Dީn?����c�u��Ub'@��^�7oB�V��7����\�+���=<�gy�2�k`��]��Is%��bxU c�k�ܻ�ab
6�!�_�`KM-%��Io��%����zv�X�����$���dF�q��Uţ�e����C��m9f��$[`���xk]W��*��j���F����T;�k%\NiB��D��P%vS�dW��j�q�l����Q�5��Յ�)zk:m(Hs���w��,ʌ�&p@̱�U�B��x��-'1�����)�A�o�;}��o[A��2➳�#5PU�"����3Ǥ�3'F1+����v��F1��~���O#����O ����ڵ��2Gu�M&�`!�$'{ϒw��q�S���5�$�]����t{�O�	�\�7�G
7��)K\���x� ̎:��߸���?؇R$��^CEGeM�;�ju��֫�8::�>%B��0+u�hCx�_;B�V��i���b-�t���D��F�#D��=V�%�s�ױ�U���<�R��	*�0GiG�홂�ә�n�� ����]���	�&0�+�K����0�n�v�;�竺�%�}��[�#���o��ͫl�����!N{h���I�;Q�0��|;'�γ��~7�Mk�S���~0<��B� GmJ���b�m|(���x����)���mq	M0������ggn��77_�=40 �!�X�~oh�Y�����Y��lC}8衷� ��e��Jv�>�K/���:\-F�#�th���+07v��d������3��R�Hlz7¼��bA�z,'K���%J�Nl(�^� �P~.DBL<z�I5.>S[>󒄨{����`�����q]4W]Y&�����
�"�ߞ���0�4��ɕ��2}ݷ���B�LcLV�:��ǁ���d���)E�]T�:���u&e�Qv��Mg�cyK�IB�n��Lh��,�ƛ��;��r|R�̏c�C�ǹ��\Kctmr����޿�ɱ}�z�BMՑAȐu��Yk�*R����gN�l�SQ�pHPqc��3*���R�E�K�~`�60w�����Kx�n{���6�V��FJ&ٷ���k�n��
J�u�Nl��R���bq}�|J���y.�\�r�57����7��߶��x�}�FK�P-7̋fˮI��H	En��=��V[�˭^���@��e�ut�~O��+��]��ӏ��(N�������>�����EL�g��C��;gb:?��k�����V�
�e?��N4��Ezo4�v�\�
$/@�Z�2,���3��O��U:q��Q@��ߐ I��SIA{z�����ݪ�"s�h�m�=]��$�-Z��Z�f���'[iXZ%3�
�m�Yx&a�]ol�7Ǉ���� 6��{�(:��M�}|�@��o?)��a�8E��C
yى��OlM���
���	�BiO�7z;�О�g%�0��%�P���k�!��gە��K����nStDq�:��o`@�C[��6��t��p��_���k���P��#�k����T-����jx���A&�ΤU���
;�92�5���{�������n�K���r;�:T�!Le�@*���
/T�"2 �Y�+rp$A�#�z��UE�LBn�7���c'D7���EW�֚���K
��U�*7��'������fNf���q�_Ј�`�H`��F~͞�B.�h�ۈvH k�9�;/���k����oX��+�b���a���5�w>�U�ީ�SM��O(n�x4U���V)O�^��'�Y>�n�@,�  ���������n�`:��Ȋrj�{���-�.}�y�%��O�������0F�ES<���>��Z�}�u�SS�	+�ɧ�
�C���3q�@6�V-�L�������8��ħ�l�/�C����D,���Y��ܲd�PG���g�&㦭H�7�#&]n�Ǩ�'��5>���Հ�1zx1f�w���Ѐ�Ż(=J�y�rf�L��u��^tvC��Q�/�0`�A]z�+p�5*�ಟN�Cn@�-&�[�F��ݠo��t����$eQ����r��z؝|^�y 6�kn��x^���z��2Jx�8!ph�4�$��Q��(|^�*���(B���5�V9���_G�6zJ�mn������.O4a?�v���ƾ���YyUm�M�����\�v���C
;�t�j�Ck9����Wl1~Qu�ɪnqyy�^d[[w��QNF�D��zbopaJ|�����w+6��OJg�_g�ļ3�!��!���l��ܕ�ژC{q/{bA�D��U;-B�]��j�&� �[�����Bc��m��5�n<z0iN>����p��{WH�V-dR[l0�$ۋ�4`��������߫�í�]�R g���\���q�i%=0�T��'6T���t�M��=-��/���]�k�Ҧ��ª>i��բ��މ�"37*����ehD@z�7�UE������L{��[Fi�<�F{�o��{�n����V'��Z���'�Pؕ��w���!%�������~{?4f� ��?h�Zi��O�����&��OF֋4��i�E�s�q�%	�f����zj� 8}Q{�.�	o[�nP�*�y������|\��1)>�^g_gm�$�P�*@���2�
̟��|��e{�-�2�}�O�v��(6׀�]�ߡ��E)�H�˓�R�;Ro�h��.�sv�>�
�ߧy��`�o�Ҝ&�m
��0t��aPOv~��AS!�fr�xzVߨF ���Y�L��r����cL_�*�^jD�\^��j�*�7�ÿ����!�c��G{�`���夊q_u��h\��?�r�i��$�F�r:�f
>��M�)qy^b��A��Ik����z,��%	��x�^ge/t%~�O���dIo���P�����a,�⑟n[��Dp+��>p���7��x-��z1�'�gd�Ԫx~$=۶���@j�U����I$�d�f�<LF���;{���.ͦ����@YDK�9,!7���,��K�`l��ԗY��uRT���ߊ`�q�%�����
tv{$�+ ><�TKL�7*��N�H����a�x$п#�&@ōH����"�$��O!B�(����o!Rj����F�|QR����m�\�I���]V��<�)�vN��z�#>/X6��� W�52�[Z�W���Jwp��'k}�ʒ�`�̜!��MP�NB*�[U^��3��$�7xuDU��se+�z��VB�GC�E�4o���E0�v�R�0�i��^G���h�.��=`Ϛ����r�vP��"�,�+���@��62je����U�Y���UWnb�b9n���,i^@ �����N*f�0�������@ev&U��%��z�G�1���M���!y���Lg���{�UP~��p��FĚ��t�m����Yt`iڙV}��Q��	���D݋)(�M`*�����y+BZ���H��t>|%���IJ�:�t�!-�e�?x��G�fi���mN���_����� cv:}�!&ԭ���	��h��W>m��EE���J�p��^��S��C(�7��s��ţ<�-�n��o��dp�FB�{X�bB����+b��%��r�'�r�W��V�vl�0sMԾ�����f�H�tyY�,g9��\î��g_�U|�>��Œ���kt��(��'�T��9T�̐�z���ugF����
�?�ǺYAC��ˑ(�0;�`.IdjgV�s�G:��cQ�� ���T�v���#8�G�m$�R��eEy��%У�N�v�{�TϮ}&�`�93�A[Gw�$)�S���7�8�䌻>rC��D���^"�'#hƊ�zm\��8��P6*<� ��aZY��r'=M��]����5��󞍮qxA������)��>o�e����9�!P�$6�iN)�l���`�#��Ķ������f"���i���~�r����59�H�3Ij ϒK/�ԥ3��	1�m�-���iKP\��ծx���P���FnS�D~����D̬U	 ���(l�H*��XU�00��F�Z�0�hj��zE�o���pE��Nb���N:8}	X7:�KB������u��Y��@@V�b,,V;��f1��#�:B �2U���WbϮ���ڒa5��14豺�U�mtAc{�9@�5����L�PK�_������T�J�`|%2v?��
VH�t���$~	B��tzغ��Qŧ̴�?gƼh}�W�Y*`�������>)��Ʒ�	�vUܶ�z�4��hd���Jm.˷�d���2�tM������[IƸ�r�FDƮ���e�Q�$0�MP9�j��γ���T���VC9�����<�΅���ug�֣՟����+XSy��
j���<��F�Y�#��/r>�lV��:0Q7��������I�jO�	,3�NUg!̞Q	D:}��S�N���#d�rD��w��ˊ�3?R���!��~�)�ZZB~j�P��
������އP,U�Z�*�5�<t%�nؾ9,k7��Q	�-a�k�c������7q%H�/���򎨔ɚ�%
�kBa��������`i���Ua��V-�!p~;�}1pf�tG1�j%G	���v�3�?�C�es��ۄ�+,m[�oY5Q�9Ù����SJ΂`����}����/�����L�K&�ZaO%`��� �X�"�;�Y��!��_����{�4 ,"��[@EA㹳Qc���������~5��쓚mUS�,:�����8��s��O�X��&�X}����f�vFٞ���	f���_J]�&�5��-�G 8lհ�<nHg$��c
J��(Y�i!ĳ7�D����E��a �{;#Ԫ<7�w��j�g��Re�S�R� ��An�s�z����AH[�{3<��ψ��g�e=�#ߊ3/>7�z���Z�%Gv��;u�!F�c�������<-��|1�(��Yဪ-�����Xr�i�$p�A��$�����v8����u�mm&�;� 0��)&1:�ȁ"F�&P>H�+�f�ʖ�>�Ԏ����aʙμ����g����%(qŔ%X��?�ܙv�?�'�Q��\��J�`�c�I�MX\w0�y{P�2�|���E'���7RZ@��_�p0��c��AS�G����w�̝3����6�/�3JT�y��"NVN�Ld(�z{*>X�pì�_?�����3n���@�\�'lR�t%.����[h_������s�j��*sƮZ��,.5��u��:�g�'���������{�)g��Y��UPpUB���]�o>f��V��Q)��'�D�\����KqF����ڶ����㎒� 4���E�T3
7���K�zv�Z��,i]�+p_����9"�H��P����l6�N���89d����,��bz�ˉ�b��ڡ�:��-�_��nt}���A~+rY$�L�D��,�|�51fT�5��[~�rO��/��62p���G���Q�����,I�����K��SE�n>���_����;7��q1��I�6��vO��?ޚ4�܄� jՆ,縣�	Q�@�>��N��!s�����KK�
�s�(�����P�kƔ� ��ڵ/�~L^�Z
ƣV4��ӥÞ�5NJ ���e���x7�(�����u�o�j�V� y�f7��S~�-T�-��{�{0�I��z�ʃ��i(�_���aԼs�H#N��V��If�iU��T�������W��!�W�;i-�ںp�J]�T%�����D�Pb�q~|5����-6UCP�E�8Ҏ�:�����u{��;����XY��]1ï�@��"d��YK�n��t�,��Ƈc{U�=sNZ�W��f ���J^>��a����?����UI��/���hF{� �܀R�i}���AL�\����<F�Z��tL�a��?a�}b	�s�&ae<$]-[������.z�F�a7:����I�jXkbnDR^���]���
���Ͼl��5��}��'����XGf�/�����Qx�\���)�@�yBj��܀B�7o�ʘ������t�[������r���ao�.����Eՙ*�tз�;��9b�k6%rK�)`������^3t��	�S�xꦤ�_j�Rw��o\��?IPCx7R�ZG�c2	�%EUa/sm
�$��4b������K��(>/i������JD��^���,�Lݸ��5���m�|56k���`�SE�S���5���k"R���H]z���iy�q���#�������Ƅ9#U1�GP|��'n!�n��(ףSh0�uFe���y�K	�=+��B�~���$/֙I�K"�B�c�q��q���D\p���42�?������=�	���X]y��P�􌖉�$߃����ڸH�8��j��5�o6���D��	ޥ{����~W�4� �p�e����`0b8��WŖ���aO{N�=�,igڭ76�Ժ$��qgs�3Ͱ���ښYhϣ�$)�ltS�\cS"'r9Sw���dnd5h��t�&�� \����%�$>�1�Χ�$A� Y$|C������]�VB�J'+�[rx�M��]�_ ���J�tJpQX��̦<7^�'�K;�U�-��pX��)���hM��W��t��%B����"�{)�]��XG�|3�{Ƭ�E�F�����kP�ц��t�������m�Գ��?�x�(kθ��|�EMq�@�ڂCsVw����]%���l�C�,�	m&&㓪zUg��a��O�`l�����b���2QOqŃ�仐j�1\�wZ�βS��f�����RA7<O�[7-�s��1f��|k;(/񺄒��*�
@�(��jzA�s~�8i�R1m̡�F��K��LX�bI�ƥ-s�����
��4�ۄY嵔^������G��jvo�N|�w�vg��e��`�2��.�1DM��N�8]G�f"�8��l6�:	؟��$��GwUv�T�a�{�㚳l|��D�"c�S���؎����4쩶���3up���1x/�&����:[ ���lun����4��A����֢��r�X�2r͍����!�����Iv��+ol\9e�z:@��aJG(�<�}Y�W��#�Ғ�1:�<.�L|d-*m����`Iq���;J�Z�qp(�7���PB���Ă��ťz��ɶyR���z��B���!�1<|Ta�]�~9�|��wr��<�>���i�#�;�E�?�+�Ss�S��6���<MF�$��莬�w��kf�:�����,� q�x�`� �C��#��I�"���'�g3:ڡ�B�(:'����J���a�CS%m���i���\��������h����t%j�Sl���&��4�se��  ���P�Dߋ��23�:��/�i@�%� aQT���>@f�]�@OGY~h֝y:R}��KjM|��1���Q��S��P������8� �#`G:��)U�Ģ7�������Z��%]�bx�~��2;ӚԎ�F ��%;V'2�VI�;[l��Ig���}���f4ݱ� �_��I}ͽ|�Q�B���R1c�Xy�J�4;�5�h���>�<CA��Ma�k��D�� �,<�$�
7B�aWE��'P{�h���[F�X����`8�Ro�$���e���=mt3��ڿ�A�'�ݢ��S{��Z$M�6�prQ��\Q1��ų� η�f�@�Պ��5
9����`���)�B�ډ�����Z���n��R�˨��/����uDHP�s�{�Ws�t�Y=ҕ]�5�?[H��"(M-�'�?NR�D-'�{e�����W_�l��s��&j��b�rJ{�C���6DX-T���]�2G�����8�ݥCv�Ƶf�
/�7 0E����e��l��p���(N��d�$�������212�w�$�$��V��U�D����YҚ��� ��D@��#U�q����w��;q~?N�l��������)���^x+��]a=V��Q�f& *�H[(�Q�
'�%����^t��J���
�`��J ���ZQ�ث0�y��ڮ�q��7�ݔ�QC'��/47z��AQZ����������H+q_�Aza�� ��2=b=�N����1h����H}�d,��H2M 4n8!��e�8���|�8!�u�\���Q�!����	�����	�4^-��2<-�Am*?�u)��#�4�6h����'���)S\�&<�����:y�IN.~9y)�4D��8&@v'���fNt>�}t�;qx���q[ߟ�d�`����G\#*�e,��z��Oۨ���1�g*��OH&�����\���7���$��0�$W>?K����L�@ڧR�}�(+�� ^ks)��8(!�ٰg�?9��t��6��YS
6z�����[�&)F��6T��RFS�p�?!8� ���MF=D*f��a����u���X�o{�4�@�.e�X�}c�;&�aZH�J�l��W��J�q����I���>���SC�缶�C���/�=�2
����II��s��A��k1�P_�.��klڹ�e����E����	C�ӈD������5��nw$�Of��9~��t��3=%��/w�ӎ��r�K9p�<ЯU�_�SA��OML��):'Ӽ��hY輥7�W�����E��T�i�_?a��9���K�����AT�*d����Mi��n9��>yR'M�'�ݦ3�|��=E� B�{�D�4��DV�Z�Tɔ��L�'i'ώ|��DQ�=&� �X�D�9���n'?ۈ����g:�c���L�%��Ia���$���n�
� �'~\�\ZՒ]�T�h�[@�2��ėj$bُ���=��%�FtLqX���׭�'Y��WP~�����>��;4M}{k��O����*2Jo��j�9����83��Mr�l��I��R���m7f����XVy�L<+���-�R�M�P���X��&9�%����#2ףj�S�jڤ�-N��J�����8}d,\��~�щ�M�`�"�8��=�9�x�́���� *��B��:x~��c�����?�
Yo�:���=nOs^�\d-��w�Lr���G�c]6��c���Ir���U'�Y����z��P��E��p���+�,�]ϻ+!�h�Ƌ@��7�TV��;5w?��{��&��B+��aԷD�ZI��o������8�1�i
X�A"���{Y��M^5:��d����~���.X�z��z�7�#b v�C�5׊q��-�݉%?�lF��[��Ǵ�-Aase.�+Yl� R�i���N�?��0�qƴ[��8z�r�E��i�_7�C~C�܀8u�D�?�n��a�,��n�$�D�ȅp���t4t����V�X7��>��NT�0$#�'s]��E�%P�bY:|��T=��c�#��E�u���_Cu��0c��6�0xҟ�Tcr�a��#V`���rw���Q��`͔��W\z�s%���@�[���C�O�	���Q֦bi��RH���e&��0����1ל�EM	ܜ7
.�@��D��LR�vÌ6��e�80�+ܕ�(��ڻ��c
Z���u��Q���a�FAa=��q~��Y x��T��<H�<R9��g@�#�q���>������6�T[�.ʋ�
��a$��P�BI]�o)D K���q����kH�f���2������O�tU��О�ۛ[61u���w�T� �`m�W%�����3�������9'�s'�$!��>J�x[�ˣ*�� �U���
��.�Q�I?�r��M�-w�Ǖ��q����i���u^��2 ��*~���E�"�F7�O����E\gȚ1��'��B�\l�)�wГ�U"10�Gݳ����� ��,P�ª���\����Ҹ��7M	e𰵹�
�ը��|a�|�N]΍g��v��-+u)�80'_�ޤ�]�{�R��&�Ol����{�Q�����C�2شV�@�,���dV��Z\���"!YJ#8�ӑcö��g���%�#e�C����<�Kk�/�c8m��9�Ւe�;��"^�_�`n��]~!��{��aKɇ�OfY�Z�J^��	��氞��h��=�v'3Cn�9�Ќ7�g�b(r.�#���A���G)�ʗ.�%���G�78��Θ��F���F�y��/����vJvϕ���g8���<ʿ�ڧ/d� ��d���)Ǎt-m �J���6E Yǹ-����&O鑑��qT?��ݝ@[�^5���Ŏ4���Z�jz��
e&=vXU/� ���ϽG��I�RA���a�{��5}�mHٮ�5#�'� �q ��wں>�;�OfY<s�3�ҁ2��:̘�h;��;���ߤ�S{/�S�5�S!�i�~�iV��a��@͉���V��B�M�(Q�m����$r���;�I��	[=?�'��\ËeN�w3k�$�Д�N�2���d|��_+]� �p���)Q�xN��\삧I��J%Y�sb�����:��8�zb�Z��R�zZHn�s=�K �l3�'�D4�%��M?�d�1AYn�Y��A��^��K��-$
C���q�/��H��ߚ��+PҺ�'�m�����L�zQG<��% ��P;�u�(`CA'�U�ǻ�ޛ�'(���i[�e�T���)�N��_�3Y��L�"��O�G��c���H�FgO�B��� �[BHmv�U�<C�w��d��-�l_�z)*J�̍�KT���:�y�?!��cJ��I��5�T4�,��8nd&�������kMO�ջ�S.��eİ��W�(Fş�[�,��C���K��oR�G_I`��F�����8�R.��_�/�UF���'�r�6x9�"��0]~b�o��>�9$�R�,?Z�6�n:�m���n�ai21miXPZ�oqq��YJ��MXa��vF,�^Y�ݢ,�� 7��4�:ǆD�曟�� 6�7�@㧕�*Qy\�t��(�Lq5��%�T��!��w?G[́)�쨀~��9�!E�~�	�/�c4�A��		�(�ɺc�����Y����}I�C���dlj����4�nFu���;s��a�%!-Ipv \D�����9�iC<�q0;-7���c�7�v�0�����qx�_�JdX�8�t �����~���(���d���FC���&�.R��l\3�E"����=�
��,V!�'��/���>6��ݝ�$�Z��sxO�#^ s����A���23MC�L�e7�k� �k�
U����,���1x��?������Y/*�
ͩ_�6�C��u��N���GV�vw�7�&i����{1ҥ�O�8�6�Y���[	�?���H�c)���WBT�{�q���z<-��t�2ꧾ�z���V��Ҳ�N�m���N6�C��Mx+���ĤU�i׎��{%�c��$���sp8���V��F;�o����	��?>���v��u���tм�IS������ǿZ:դ��m�6F%4�]H�t��w$w���+��5��'�y.�����3�F���A_���i�s,�+:l����7TRI�1�\n��tcP�?�d4�!:�z�C�m&�]�W7���!XMb���PX��x�g���I����5B�;Ga�؝�"�,�x���q��W�x��8)<@��� vę�Ȁ��=Y�>�t �cω�<�1�XLZzԔ7S�K���p��?i�z��g�1Ԋ�K<ĹM�ڧ[�1��2Qo$�"p��XH�n����Ӎ�X�%�nb�x�����?�����$����UN���K�4;D�'X�-�U�zV�2<�7�$��B�)���ꦤ�)�ob�	1�D���!2G�{�\E�MR��yR��΃�Dzܮ�l��[��c�)P�u
�s
��+���JJ��}��=# ��`�wm�cV�ン��e��Qo�{�^��&�esT�b6(�	�Uǽ�}W綗��> }�e�\��	Q�^����"�vp�(A%�M�Z����C����hh�8f���G�@mα6��F�� ?x�wwJ��'��'�^CoQW�!0/i��$���A3gl�-C�s�~��i"��B ��]ǷӨ���\���?*�5���:��XDƲ&����97�h`�+�
�1D�p��JŤ��Zf��/�iE���){�������pj�@t��퇩�s�-h�d�K�ʶϛ�C����y=b��s�`h����G���<Q�;��0�.��d��wj��E�hM;L�r ����f؁�%uK��S9�� �����	��뽈%X�'��f*�X|��䆟��;#�>�H����xoNV,|�����'���2��� �N"H�Y�4y�BO�`#z��EU.9�[!PZX��(��3a[[k��w���gኅ����� � �J����	WXsےz�i��T���������H �����F���QF�����]0�z,�a5�mmU��_���A�>rg��/���o��*�!D�{��s�ŭ����M�]h_/�G3V��Xr
{~y��L:��m��iAgZ��M��--�w&�s�@T�������װ�LA����K�ê O�
�m���Iz�}7ӻ$�r酀������ɷ߅�C�wR?ҳ�q삆\G��ep�e�1^�m�]չ�_�����庩?��ΪY��jX��А��f��k'&O��HO=s,��r���o�5��2�d{n�o� w�``���go��w��NA��z_��,�Q��a=,7K�k�ky�cDgAw�Ǧ���	0�%�����/�xs3��BJ��-0�����ˈf����.2/ �_\�*�9d�G	[��U1�����r��w��d����y�5KTQ@��0�2Q"st����<���h�_�p��Zб��[/ʔ
���RV��nӵyR9�bZ1��e�%�>ʝD���lMύ���6��|��������!�� � ���ɐaR@���Y����ꬩ�1|�����ൺ��fVHj*��W)��Y��g�D�[�1�R�P�Ɉ/>��\�71�7����\d�:�@�0�J�6�ڟ �^k�f0D{]M�gO��C�$��2��E��P�.�G� �(-f�J���3`MG�E�
�ߜ=,���3Yt�!�tB7� �V��B �}�7�n�d���M���paWQ&^�> �:p��A��;�?-�R��8uB��2�a|^@�r���1g��sH;���YW�)�O�=��o(��ϳ�3�V���jm�mw��fݸ�6MG^響r�"�u�F	GK���>�BZCJ$�@�Ѳnn���n_J���C�?�M~=E�,��j�!�4�?O7��]覯���O�.9x�g_D�A����h�W�S��%,��O���V�>ռ�V���z�S�|��H� ���:���0��%�,W�-a
�'�m�|nO��%�T��`#Ơ^Y��R}��4 1+��l��@}Sx�Mx�"�-����zTR}�h)rd�K�yDx�j0�V���1֞Cd����wA(���T8���~ľx^���`�����K�y.+o�B���aw��+/XF�k�É1͔�)%ӟ�;ņ���V_��XT$"0ޭ0�Ws枋��^�����x\,�L �1QN�.�h�,����Su���Le��ᷢ�pr���$������A�#��1������}��F����7D���N`����`fZ�e����~���-�հ�cV����008~<�bx�iZEʀ���V3Qp�A�^�,�������#w����`DTk~r2v�{�.r����i$�=\�8��
/WQ�W�4�X] �\^%�Dᣯw��ۅҜ��h�c���XCJ�/
�6-T��SB�<�C�M�9�,~2| M�M�~���`��Θxx	���;�s��_��#��
օ�R�띪B�z"t6�c����h>���W0�=��"b�r��<�M�'pΣ�N߁"7��������UN^� ���TAe��2�i�N�sj�蒼��s4�Ȯl�#��� ���͍@��q����z6�f�*�]���m^'�e �<;�ɬާ��v7?����[�u}�A���7u�Pppjx�����dܾ���KtW��ޔ;� ��O��l�b����&+'�iV�@z��%($�.W[Z��\�U���	�҉�nd����ib�6��1?r�44uY�~�:q2�5 卸��P�:��#w`zGi�U��0��Zd�b����k5�b|����"�ꚁ��<C����ڡ���i��6	tR��y���o:O%?�w�k�܋ߕ:�<w� "�׻�o��GRyCL��/�@��n�)��]�Bg�r$����# >�d��L􋠴��'�m�h�C�����8wQd�d�z� X���Y�"`x`-�;���-��#�GT�!Ăʋ��p�p�['��T�V�����<sx<l��$J91�T���h%�i�0@x��:r|� A�{�6���W�m��ȵdЦ(�N,�.���h��z He}�x�v��R���$��<����k}�^�K	�^�q�Z��YP:�}�uV�O���0��8iVcS�Tqs���*���*O��w֧��Rx �t�Gߪ�7��dG�G+��8B�"�ܪ��]�/fc�b���p/�5]�2��RD�v2j��e��A���(*��S�'&	���|�ʅ#ӿ2�&uu~e!�s���e���n�[k�Z�� ѭ��@a�Ɨ�6�����ծt�=.c;�WHU����4����>��\k�?�gL�^2��9{2w����^�qf�أH��M�@�;+)��(��l�������,eEmӓ�xo^�mQ9���IZ�$Tz΅��f�?:�v(.���6���Щ��c���ȳ�?۬�l�codOw�}ep������3�U�#�|-�@���V�kݦԺ�4��z�_�Mo��:�p����;�\�PS
����'������.ـ�>�~��S�����N�����<�;z�a�U�|��(��c�(@�p���l9�z��MS��ᣛʈ�.�n����=�C����'49�~������>r� ���ݤ���=%d�f�c�2>�OB��Z0Sw�e�?�mſ7��B_P�"���2��ݞ* |��0�r��Er�zIEDY4xof���}a*L܃������Ռ�&�Ⱦҡ%$��g>7�%�_>���_1�k��gcz=����d��{~���;�3*��e �G�\-��lgG����c`�g� /�v&G��o8n�|7U��6`�M.�{�I�����$l��g
������By �o�6(,&!�Z�oj�y�����Cn@O��׭w�rI�(rbr�2M</b�FE�J@ڔ{�l6⥀$d����}yر4�~�T.a���l.���j?å@T�^@K#"oH0��d��A�=Y�� 9-r8�HzT%���
l�S�q�|��韀Ej�w�U"��#ȡ�ʾ"��M@g*�[週<T�b�PZ4��7|>�v�[~@�d ��vwVGb>�O����/r#Ww!�AX��ۥ�#����j�S:ئ#���׏���s<bm�͘���/�]��]'�p$6������[2���*�+�-w���a�ç��K/eH\X�{��gCr�@L�3a�3�I�m�=����k�����d�-R���n�������X��ǹό��-��*�/ϰ|Z��<E&v�����a!��%���%n���d�둤l��YLͿ1x���#7�\0�	�68���{�(�����m�c��% y��jӜ�~.R|@`�"y��'�7��7fu�,��r�u�JYE_���kG}�{������.1t��(�������`�bu��9���bs��zC�`�D�i�*Vy+�`}j�pF ��)��w��iw!L�Pu+�����o�b[�Cj����W�~��N�W�"��da�R�ap����������iy�mn�-RD������̞�2qy�ɱ`���4q}8lA��� faf}w��<n�8���m޾�_�m�VcA� ���Dr���!#O�EsF�6n�����fH�n�(�X�B�@���)r���'8bfA�Ӻ�(Ew6�I�S�y��x�r1͍�<ʖ�\uʺ�&��;�+-n6�EDQ"�y�z�g_���J$���ad����<g���շ_O����Jx^G�g��'լ�� �[� ˌ j����c����4[�������#ߙ���R&��A�(s�
�{T
XSZ�o�v�p�����z�����`Hn^quc(ߔnK3+�G�~�˾'9b~�r�Y�k�"���g��2*`�`ڬ[ppW���l��[vb�/Y����0Ƽ�j��1ˉ*<���d+��A���dnR��n%s��~}߹���N�=��6�1c�'v3��H@�<*��X��2';�`mwyk2���-�3�g$��44IWc�oB�v��1M���O���=&��q�Q8=���_��H���<D�F�R.-G�Q;0)
������`��P��Q�3iD��w4�x��C#ml0��Ԥ����mb_��9�X�d{:+�G�����:}�xO���:�������N���<$���$,S�2���?/|�VsC���O�����v7_�i���n���0�mſ^ǥ�b���!�@ǔ4��*n����}�Ш��a=����L�*��Nt<Q�TH��Kŵ�
��h�yQ�nM��n&c:9r�`Sv���+�1���?b�@��ʊ"��(@��0�	�����n�˽n�@�#���:��XS�U7�6@�����������7c��yĖa-ݽL�֤*�L &�"ؾ���H�hx�q��eXqS�510�B��	x�n�#}t����d�� "�����8�>V*��@�^	���0^ɡ�o�Z}Jgjs� ���tЀϙެ2 C�(����;�}�w���v-=xh�����-�|�G� ��W�[sc~�{�D��!��=�i�Ɗ�?X����T�	��j��#XQH�TД9 ���8c1�7QP^�FS��Ss0)�ph���6kX���7��[,��4�#RQ��,Z�Y��E}���d�I��5)����0T�^~~{r�ܿt�F/��
�$��"D�s�xإ�n�����������x�ϋ���P}#_{�N�q|�tР��&�f�:�2F�����~o f�0�"W�~��,�&pV8�c��
V̻� C�P#�l�t<�c�Sp9wC��>
��. �^��z_4\jxy��a��b-�S�p���0���kF����4=)���k�tt�H��������,��+Z��a�H�&[lR�k��*���'���菒�ݣZYT�UYgj!%�y�6�[���tb��f�������I��t��puI4-yd{��65�'5W����4!������/�@LOİ��Լ,:y'���1/ٷ�@m�=�'����*I4�PH y(������w�p2���`�M*#�o-�p5Йc�~y�D�Z��!�N��R	������_u�ݡk_ ���'he{Ѕ9+­m�b��d�Z!�	��nW��#�M��Y��3�խ�����]��%ԝF���5H LJ��@�8�ip���T���2�r����4���8@k�֙���Y�ʨQq�h�g)�Jl �`-�
���Q�R����(0z���M���y�rI�1]V�
�V�f3KRIߡ=�lbw�"L����Y�tip�I6� P�&��8���*�vGp2p<J!�mqUl��8H5f�g|�����6��8D1kĔ�Z!��[U)�F�N�|ɭ|�g�Xw7�&}����BW�|_�� �U��)n޽.?�"�<�p�f�g���D&�e�ZXB)A1�����^L$�k���a�f�Hr+E�P �;���O��5L�L�8+W�>� ���%���L'5y�9���/pf���FA�+�ε�+42XLl�u4`�K�}'��~;L-��ХXF��^�&aœ#�Q*��N����w��k�슡ypii�ҿyC�}�i�+Ul��i����s�Ð_6���X�%0��� ��l@ ��~�w�ֶ�P�٫� ��H檮ES{	�'�W�fLe�N��������2S��Md��kV!�H/��"	!x�@J(ªq�2^Ku4��(���+Z�U�❉\�de��r�,�4%���5Y�R����E/��	�����/ڭZAQv��H�3N8 d%�#�?/���б�H����=�Yx<Om�l�՘=S�;Ss{(�\Ҙ�"Ί��$3m?������$b��_L�5a��	�j�(�r��92�J$]���C
`�y�I�!زQn�H�n�9hzU�Y��0d���,��Ma��Ֆ��9�F��p���b��.���95l��o��?�;��@u��XΝ�����>G�����U��#Y����☉
^��6Y���*ʠ��cD+�ڌqyN��x���i;��T�_����?��76�5M[��UT:����V/��������Э!x*���q����h����ʩ�
�ߊ :�N��g*�,��7�����X�ۈz�a��
r��>�Q��ɖŇ���E������Eؐ�&A�����I����1�1�5>:G
�5Я�J�Y���/��7{"�TS�)N)�FU�[�M�l�)Q��%�/!�no�$��.<B�d�0d�&%�G���o p���Y2U1���B�L�/fK��
$�<��R߇�6���W)2S~��;*�й��l;�^�G~g��[ۨ��\�/��֮�n=��������?�9����̇�B�hGW�䲼�0#oD�U��͓Yj�v���v)�)ۋ��3�\�{>{��Y�٣��h����?`[�x���I!�o�� ���Q�y���]H�N*�w�L1���m0����Ih�<�j�<��d2E�͓��#�^|�Ц�����:߷�M?�?e������oB��_F��0�f�Y�jjEᤙ�-g�h�hi��gvj���J2y�[��Ϲ�����QnM����ժ�Ä��.$�9^�{��TR��%#⹬�ʉ+L}|���W!��/il�Z��a��x5*�1���������wzc�tQ�k7���/U���
7E��%�����;�2�H�x��3�q��wX����ӧ5�ڞ��q���eQk����`9֢tѓ^T���G��I�a�%���aR��)���W��c�Gqǋ�kl`�Y�_:�k>C�2��/� b�H�3̽d*k�Ia)Ԥ�Tc�`�,�|K-��׈��8��2�^�h	]�m@t%ԯ�8�*%�Y�Ƙ$��Be'��f�N�|\
�rg�K3BRw��X�$~c�$�zC���������@V�<���r]o��P�W���$����O?�H�v֭��jd��e~U<h��|1Y��:��a���9L(_xk1x>���~���������◥28I��#��)����by�ɹ5��b~*�7w��2pn�S.�H�\�9����sA�y���AcWGN��X�"��l��Vƿ>Y䌻���m����&��ϳ~CE�}Ȓ��f���rc�j|lG�I?ߦ��g��2{���x�X�(
�Z����
b?Gc�}�ǝ�|���#�u�^`%Vkg`�Z�s��}��C�um���wQvt�<݊P��`m:}�dM��R��h�ַ��vz��kG�_0H�߈Z�X�'-����N�u�4�`n�9��n&�V,.ɋ}N�8w�x�·����-�O�*���JW1%����p�E�B����DD>|4"x�k	����V�D6�R�r�c�vW	�z�p�q�j�������!��B�E�ŁBin˙r�.�=~��'Ɲ�Z�x��x9���_��l�y͵ܳ�g�W�����3q�b:34�vK��x�g�Ҿ�cL^�QXq����'�O���O��E@e���?ꛚ���&Ya�Iy����`��x��!����)��0��'���H ��!�3}c4x��y	K���mV�����s�����}��}�8������±�ǡX�pg{���;x�Y��?�:�����|N��~��5���`�(���\���<�ϥ�-`�t&"�����)¹�$5��ww����6Z���3a���`��a7��84@�Bjb2�ڏ��x}��)��e\��V�e)@�����ߟ��{���L��#.�:~0���y�xo�w���ӷ�BK�+?��0)5ބ�B�dK�[���y��,��t�]��BD���c{�H��"GK����0�O%�P	��\XR^�+1WR)��\|\���i�nhZ��c��{pk�Q'ZM$��c��@�1��;�DJ�Z�)[����&Gy��Q�isfs��?	h�9&����t[����T� ?��ʯ�Iȥ�UZ(bf%?��~���r"|Rs��ԓY��{�!FE<�Q�����Ћ]Cz���0������q%׀a*i�'r���Q�7�mɎ�b�坩�[����ħL&4k��\t~ܿ�K^����~�_"��wwc'1�婿��A|a�F8ą�C*��6rn��n��Aw�<���NG�a	��w���)��yӣq��\�� 
w�%��n�/(�V��1M����x������A���F2�Jz���i�	bi�۽�����N�D��A�l�ps�J�Ƭ�H��9�Ɲ�W,�墡.���(dZ�jX�Cze��\�d����H��f��"	N���#^Ȧ����9^�jjm9�p�U�mC��GbgYr�y����[D����۸��nŦ��bЍ�}V[n[�^e��t�m*�ǽ^Ӷf���㵳q��4����'.H�=Lg�z8��(d���@�.���LMYS4�[�i��
�y�-���PE�ex8"�<��+�U��)�_�\@�}9�-����5K�Z !<���I�� ��4I����b����xW�.�B��ʏ7CD|�oI����X�\����	'�1�P�%�7�.[z���i�8/8֢_f�d]z��g���B��,����p�������C��qul�n�yO����C2VLѳ�L�Rn+�h����,
��X��ٲ��kT�bP��)�!�j�n���<N�\j��_�'�f�~�1�Wj8o�rd׻�{��
񈎉Kص �ۚL��-ek5����$�Py�OX1]bq*�N�K����e�A�W��������n��5�~����/HS�}�����[��ߞL�4�>"�K���>�kgp�P��r��ɪ�5�{�tc�"�j�	P���.��7�ї�l����n�15s(�#�
_xa��3����UtpC��}F�Mc��S(��& �x��#/|8¯���`����~�e�S N	/d�D9tQ���X�Vf�M�|�NV*���~��SD�MN��Yz<�����\���C�2(�|�A?���=ٰO-�6ɬ�z;X�U����-�G$����^ސ���0�o)��Z�T��B@@�3�'�\c�"��5��gf���Ê4#zsL.�P�*�U����XP�z�D2����a��]��\BF*�㮒��7�[/��`�"^Y[}��;�㾠�KÄ�^�Y���)`@�r�՜<�H���N�'�Ƽ�,�"_��*8R��WDX_vI�����]aǟ�Щ ���k�{�6̌��U�&	n�[���"n�]�}g?;o	����c:�W.�~�Hn�bL�W� �4}�Nu�n��9�ψ@G�&��k_y���J;ҵ�H�i��Cg�З{ʔ�����B� hڝ�<�O�q�?kŰr�ڭ ����9�B�lZ\ �Z�ZYϞ��IAV��c��Y��	C>��׎*�,��ƙ޻[��5�UiL�"��>�$�IT~�?o���}����6;�H=�$�gG�@�"�=�ju���9e�T4{]q���$UE������<}�`	����´�T�|0�]�|�Q�/����B��R��AA��]:5D�k!uA�0s�Z�'?"����ã����a**����w�ڂ3M��*7�Pa��>w�<ޣ�UƳeV��� &��Ծs�k
�ܑ�����r:�����a^�F���w%����<��V.؍���.�&a5�O���יA������s�Hi��5D	��L�D�]�]�t\z xl]�����;������R��bf�o�9b������F�1��6}�VV*��۟ہ�i�e�a����2_��� 8]�_>Rlv���sj����߰^�5�^�s$�K���:�O�m�f��53�ך^"�q7�bk\'FcZ$��]��shkm}�u�O.�l�Clw�?����Iq;K;�K�艍�d��M�$�����ȃs�R.N�,��g�G��XH�K"�i�\K��+-��`9�j���>��l�9_�nK���k�6�+��� s� ��N�T��.yI�>!p���|�-����	��n1�
��1�F�k��z^��+۱�ȣAt�g�S��֡vA� ��K]�.��b�!�2����� �	��cҍ%�4&�j����Z�P��~cKX+p��Z �-)F��B_y[����<]�G���2�R$�fÛ�)K����Yj�C�M��l����W���C���⵼W\I�^t�c뙟����4d��@����
��˞3�I�r����h!��1 ez��ZgaY�v�Bñ1����#���]�l{HZ�B��y��[<���Qx�@/��)�^t��d�G����.���cD��5֓�#e�I����4�W~��y�h�O<� �H�z�
'o�f��T�V?((>ː�"3�JΘF�J����,�&�9;�����Ƈ-X����o���<�+o�;��_�"~7K���x�3!8U�a_�&ʑ��i5>D:D�S��Dd�T��D�r>B�_q�C��O��aN}��H]e�;�=�1:��!_
X�p���
��D�h�$����>��^��s;��;��c�\xa�q���m ߩx���/Y�B@�:�T����������%����>jG�_��ŭ�Lz�{k��)B_�����sN�]� ��jo��/__PQЄl�E+ꢵ^����E���t����ou��5J?���'(+��INJM 2��Vm�t��n�&�ᾚ��&Z�@*Q�2� \�,l:�F��6q���v-[�R�ֿ3�!R"��r-����T�%���&f�8?��U����}���D<��ɱ��(m��m�m�1.��kTUA&l��vђ︀z�z�v���o���Ơ��'���>�'u=?}�����E���u�t��D�W<���q��(%�Gtn��s�A��c�+�D�֞�����Hп���K�� Xۇ�F_���۾�	]��zu耐Y��q-���n|������\
҆0����L�������C�3�IL-�G��:q�}.j�]�2-�l$�@��3VЀ��ރ�4�#0�Q3���U
 ��������B��Y@�8�N�i�o���#;09�k�K�A-���->�A�AG���	�%�ˊT���n�p��b�O
kf�(������GUB�/��h���&B��0�����!]S��cy��U�+Q�+���Ǖ�jE̖���kƣAy� 2H����J%�QN<w�e:���e����沕5pL���4	��	�O)!I_o�\"��бm��7CeK��������<�K�˝ �T�3��� V�����0�7�8�6[|>	j~t�{c��Eb;N�{��uˊ�/�Y��m�څ̂g|�Z�k��
�
M'�w��Y�%��&��M�C��lݘ4��}]C��6�C4��jo	�`8��YP������]�Ա����Ye_�ǣ���U�'�+��M�
�QP����[Y�K"��^��)���a�����	����&���h��Ti�6./�Dk�02�k_@�*&Pړd�	��*�[J6-y�����ݶ��O�wI��>r�Z�I���)="�(\�=�$3�j����a��}�~P�O$Vo�k
q��mL�d����'tpr���ԷI�Y�g�&����XN���?���-2��49�/�<U�����u0r>ۢJ�C����
-��K����h=����~-MZv:㟔�)�R�fZ�C���K�Z�v�T��B~�����T@���#˴n�������oz�4��\g¯Ҩ}� ��)��Tk���3�Ȓ�sث�_T�d��0{�F%�V?�$d��� �a[�O��ڕ�TiQ�:x�!:rN�P��z_�7
���3qDe?�'b����"��� ���M��6��g��h5��8�t]+�m���M�ϣ�0�C��U��z�54/�W8"_=lt��)�����(F:�'�m��^%�S��_%Oz�o6c�R���2߬�&�K�4sȦWN����ªM���f\E�c�����(l3��M�l\�ՊQ�4�Na\�P��i=c�o���ɜC?p��2�; tC?;t�;��&@(@���d'���{�����60�����3�8����k8�P2�A���=�� �ݥ���$J��#����)Dϒ(޵F��ko���� �k �B�SKZ�C%��~U��E"�nl?�ү	;�H�Hԫs�� }�.7>�pt��$�2�%��JH� �P$�/��ޅkn�bHӽEZ��1�&�G�i��A�;2���/�+s(I�S�*�h���_"��a�&ì���ɡp|D��flf��2�[�%g����e������N��&�a6Q�jO~Լa�,��
��qi�Fv�
GEѶ&�__9�bn��a�X��pr HX��ă6�(j��Xdﾙ�ع1���O)��������{v5ఙ_�C�=�����>���.���w��Ū2�8�L��R��?�1����n����3۾�A/V��_*L����ތc�v����Q�fc� ���dB.;�xF��N�.Be;n=������/1Q�+�x��1�"��Y=���'�E���(&!͕O\����$C�����>�d�.�(�#Mg�Ȣ�+g+�\�"Q��vĥr׮��G���=���8u1J5fi�
dNA��_pS�jξ�r-_��j9id�C��[���f�p��C#��$$�I;�,�'�#5�F��G��f��yM��(�Z)t	�)����s�Oi���������[A�"��Z?|U�\̚�q�΢i��փ�z�o�m;{9���J1e��V���TU��ߪ��6m�t����d�V�[�� ��be�社�(w=�Z��A`��"�9�ץ�Z�
�r����ңU^�>�|��9�~�3N�`T�*U��(<w!���L)ݘa͞A��6�s��%���;_k�{��nF���2���Q���^QXj5�cc�N��/����]X#��\v�~�mp�>Y���;T�XK�����h���}<J]i��-$y<�a=i2{U�u����#��y����eXf�?6� �%q�O�?��hx�f'� �V�GKC{t�EH�?nQݐ|ʠ�n8 =ӽ;�eqg@qe�Q�3;��I��< |+���4O]2�����͘�pg ��m�ق7��az����=�|1�Z��Z��E�"�@Ni��g%��m�N�|�d-#�-2F��E�Z�h�ǣT�&z��ݴ��tsWc0R?��P(�k��ZQrR�d�u$�M�3k�\2��YjgϓW�"�ٷaA�,5����;���v�,�粹��JŽa�sw�ѱw���̈�/�jE��	'DHp�#8�����,Kw��#��)J�PG P���x:�p|�c��q";8ϕN���z�	n�@6��89cv�)�F��j1w$!���F��+�(�����u�wd�f1��*a�b\�tE�"a���}?�D�z���=�	�ϳ��H�C$����2��Bo�}�D�l��S��@��`�>�JEH����\P5���"���.F��������!� n��&RT�2�[qT�L�@\�*��2�.���9��<Z���3싨*#�30��S��Wq�<��\�$A��Y䠤Wt�番�u�6�97����uB\Л��)x��	u��]��=/��<�{S6|᷍������� ���Y�t�%��w�v�u`R

Sz`Yf�	���9����x6m���V�&Sʨ#$���C?cN��R�-�Wm�|����1�Z�yY	��������ߴ���ŭ@������8Ƽ|jD�8%�qP�D�.���� ���("��^@��0�E0{Mh��HS3��ɡ�o�o���x��������w�Ib��YU=2����c��''-j:XP�����=˼��ꔢ�8׎�>.g���h¸��� x)g���T֌����B� 3���VB�㺥goz�����0
�ɖ$e�Kt��J_A!���[�} E.��L�t�6�xx�Ge�����+�cƸ@l�4�[wy�$\SM�Ԋ*y0�=����<�8t�,%܇�U�֘}�;��b��f\�*� v���M�t�D��;��u�����.�F��#*�&��E �$�s���] �6~�C5;")j������%V��u��`#��s@�n) �����Y�X� ?�E?�3@�M��EFH[��ꅼ�a;��Hu�@?�0�����]�� I'�\F��"W�O(����(�;���b׿�k�h�����N��N[�0��C�����IP!k4s�Y�&@)�pg�ȭ���-�S��[+@�o?"6�Ԑ&,��0��Z^Bs�H7v�d��)'�����l�H���Ko?�_`\4�-��%L�:��V �a	��-b�>���t������Ӷ[��4���Phr�����_!=�y|�R�,�Ħ�[,`_v��h�&=e+F^�M���V!�����{Z�K`����.��Tv���)s�%�T��B0�q��t-<�����F��zG<���@#<f��>�E ��:�N�B�U�OZ���v��#n�O�r�ǖ��
Z!a�?�3֍8���=c^yL��7�8�������ѣ0e`����c}A�&r�3���[��𐵪�{VX�Ji��{Wĳ��m@D�m���"���@�A�&����PO	��pg|��'I"��Tu�j�"���J�B��Z��&Wz��MjF�8�p�l�|c�V�f0�-�t��l`��k,���VEݝr\<C���@w#ڷ9�<�O��2l�Cd|��� �7�*��Z��܊�:Pi,=$��l�b�Zzi@���1�:��A�[�~ 'y����Y��t4��U/_���A�8�;kKe-�pw7&'�!H!���El#t�`�G{B"����[�g�}Iņ���*��H����	�-8�l����r�܆�B̛����ER��C�	�5.�j<�,Z.���N�9a�"k����9x����K��?��{�$�S^(�Ȅ1V���]�����6�v��k���q�C��_�Yr[Z��n��8�͐��*���@�D�N��%�{�
�!¬�.I�4E�m����}��A~���eO~A�wd��mf�3�z�Z��("�}a�Z?�۞�oa[T�xu��p�ӗ|�A޾���I���qo<��t�-��Q�K'^̨�n�fJ��!��q^1�&����9I�=���"
�C�1eL��b�X٫��]��JU���X$9q$�(+���Q�,�o��X'+��z����+w=����=�䈾VL�ߕ�r&���ӵJm~�>g�c*�at��r�i�*���Cn�[���^�^r���c�_���U�Q�}G&J_��Q5F�����
:��ܐ��
:���F�?��;�Q5`���ڣd:i�;���k`0/a�~0��?v�5��F[�"eer �m�䭄N���6�(���FUY�:+QL,� ݅�c>�qN����Jd��+��K�?�߹It�+�>J|`���;�3�>��z`WH=�e��T�;M�����,i�C�j�<�X�I޳�K�*����;`8�g��TX�@��eʕ+������K���Kdt�&���e�:�4ڤ�86>���A�s���R��OG�Hh�=�ԇ���Ɵ<]�M;�z?��k��!$��D����+$J��)�>:8��&�U��,14A��K�@���<�B c!��|��(���egS��!��)*O[����ߖ�����I#rB`\�Е�.WJv��r�<`��SB�6Zԩ��n���c��M��R���zP4���,q����bˆ���
�� �qQD�r<���`��1 Ɲ?��,'P���fY�&� ��o���5<��-�2�#��=��V#��hA���3I�ghi���@T)�wD�����Wq��[[�}Y���ly�e@O�GBvM�B"u�S;�]�F�h�a�=٨��Mb��%|8}�FV�%�֙�5���@��ؼ0vz�7J���{7�3�]���أ�	Ni*���s��^����o'I�ם"|v���ޱ0	(��d&�Dy�!.�:����*s t��6j3�"�Qj[��v�>/߳.��ӑv8�.�B��F��<wg���L�[���A�;Mf���0Y0�D����H�zT�p�s8��)*j,a�l�,&dx�!������]a{_��P]\���7B��}~���Е���ey%~3݋o��09jQ����<c��V4M��Қ o<�*t�������%q���������F����x���j5}���oZ~Q�>9��)��a;��u�۸ ��b󈂻;�0��_!����|��2�_��T Q��W�����g���i#.�V�W����@�D���c�z����k��ͨ1���#���f�&@pI����2�%B	:,e{��~-�e�QB����xJ�<U�6�H<>��[u��;�.4�n�8��M�De��.�[b����Ķ��^����D��q+�8�G���wV�j(k�����&�;+�U�
�+򯈚��@[�+ �`��ZF$���$�h>����MG!�����W��s�r�b���E�&��h��ll)���@�̂������.A��~r
����	��xS3؁���{^:�RxE��F\�����W���nF��Ef�|�f���r�HI�bIJ^�,��=&��%����\�~;6"������F�R���ȕd��� ̇��d�*'R6�v.�0�����^#�6�H�*��8�|x,P[/c�Y��M�KX�!@<��ɠ�m���������ؼ�:nP�ǋ��!Qy �����B��PWԍG:�ԣ�B7���;�� J<r5�3b�� �ہkϨS�Y"����g��i`:��r�Gx^�e�!�&�Nc���0y�����6�b7�"6�_�v�B��n���˯��[�:BT��6�۪�O��?e��qW-�	�ǭ�p.a�zL�7�0W��TB��j3�8M^��k�thsdg2Z���K����1�����ב0d�
Y��ʥ�@���aI/�	h�Tl5��.}�~s��5,����#0�m�����3���éa=c��u������c��f*��tM�Ml;}b�j�+-~8wC��P͎�< c�&��k7y��ێ�OjF4)e-��l��ʨx��sB�_�?o��E.���S�o�~��J-Y�k��yq������q��-���Pi��,>j2�f��7��
�����X!�Uv������@ZO��Kk���߁uK1�aP��kj�����Bz=蔐�|�
½6PB�l�]7�uV�e�+9혷1�S|i�O����ȥE��������w�3���3����Z���l\`�j�Y9s��Ko ~B1��$>I��<���q��5�\���U�i��*ّ&n�,�r ����V�ƂD>��!��F���-�V��`�~�lT���2���M�#�̢���1.�y6�/v�:��,�����b��b��2���0��6� b!����>,�����?1������5�p��%4v1r���2��-�������]�����c�7�^�Ls��:U֧,�{E^��z���� Q�(.�&h�,Ռ�����+�?*������Q�w�����'�Y�ΉQ�Ka�X��<J�������)�gހ�y�A���r"mtH��]6�����ͽ�/g����c!�cG���&�h�8��S!*	0�B�.���9��.�+�� <hʐB1W������yߎ.��|�

���(˟B�n�<��S���@Jai��~r�L1��e�YqN+׍��{!X9�`�1��Fb���T.�!�6�������9km-�T>9_d~�U(k~���-�%{������C�Rw��yRx����W����LA
�%z�a�"e
AN7��D/�k����!���25���JK�+F��s=CM�1��曨��-2.FIO֡6o�\p��PE�P2�^�"�������E��������S�A\:S���[u_bv*a<v�q	�
��SK]���"!d�W��?�0V��Y@0��ԫ�қ��Q��͹oI�&��)�S�)B��(����O	x��nG����`���rw%R��	�zm�}�0�$�Ek>�x|�]oB��a��zJݬjDp5��Ll�Q�i&sj1r�<jT�a���S\��8�l��&�7�w0
��V'�Ť ��i���N�-��8h�
Aj�ԋRo��n5���{��q��j��Ui �}��U�&Xx:��-4w;�#�[�����pYK9���Z�W�}!ߔ4���HP�����H��m���W�4�Ȅ�+X<�I�Ł?^����� ���s���f�Ԗ��[��B�Q���vB^�J�[���T��l5��@�QʴW��Zj*x�C���Rw�HacfՃ\_�ymUٕۥ����3F[����G�v
#mc��K�z��
����m�#���B|�}E��q����5lZ���_w�ݒ�a͋{��d�/h�ΖE�P����Kꋐ;�D�﹓���B�Df(�s �C��m���`Ƽ�3�>R����r��� a����54�[�zx��E�fSLn���)��HK2��wQƩRYv��ҡ| �O�o���ccS厺q@�^֮�qPs��Ww;������7i���{��nT5���l�:m�L=�Z�%�w���)��bP�U��*O��W�n�e���K3k
�ퟁ�\BfK.qTNr�P^�q��q%�-�7��������[jG��*4�����q�A�P�$(�#[M�ǚ�Pu�����^t�i��yA�7�z��E�+{L���~�h��^�����LǴG�B7��y�:��Mg=,���<����,#����p;OW1ֲn���
�F�HI��Z����K������w����].���T�TEc�����G)�Q
��Hf��iK"���z�J.������C5"�����/i�|��s�;<1�|h,���aJ�Bѧ�֘���β�~@��<���b
����?HC;%�������?ƢT�{Z�0+��H���{&�m�#ZI�.&z��)W�!�nʠ������������I"=�;�f��&����Hޟ��D���.j��7I�GY�բ7Z��#^�;�&k��������8Pmd{`Ev�����"���h\�ɺ4=�SX��f#R��7���Y#�vӫ�G{�d�1`#?3�m�܋��? =y�cR�u A���Ҷ�V��I�p�A"�i��j�0����¾��E#\ܓ���uoVP�&�F������ـ�5�67@�a7I��'(���΀�ѤU�b���P�`p"�5��9TR&8k8�vx�������%S�$�-tC�ReIV�i�O��^E�P�U&P���g�kL��D��d�~G��f��ˣs�i
�`�G�*����`��G�Mߊ�j����k�dP�����G
��E��b��}c� T=Be�1�Ƙ�h5�[V{�%~B�3~\�H��iۨ�"��b�|�J�4�o~��=�'���������eMp�B�x�&+582�������;72�E�f�^���|cA_�Y���lGuӌV� n���9@,�gV��Y.-�J�Z[�.	~�A����JS�+��E!y )�@�]�z� ��`�Ъ\i�8��G�W�&] ��jM��0nD-�w��I*c��"�n�R=TҥShV_ʱv�.�Z��S�[8
0}A��2vK�
M*�uD�UuĦiZGy�e��/�0���jȝ��?̖"G$&%ɬ�&�٭�ͭwb��i��fk���i#i9�j;����إ�-e��Rf�2����(���	X�Iy�J_�o�N�S���c����j��ZC����/TC�̸vĪ��y|60Q���)�W��T5����j��$�Z�1�A�ѷ��H��1E�y��DML������;��e���0��
*eEM��2З����ކޕ���Qy\�����Q�*��G���J�� @a��Ά�X؀�uxQ<�u��: �N��v�#].���d��-%��$Ɛh�P�H�`��x�����S���ANɖ�L[�I��Z���u*�Z�n�Sj��m�穹����ɱ��e�p����o곆�h]$3yC�V�ʨ&k�+���ڡ����ݕ>�PS�f���G��72�(����ʒW�K�1Tv��j�'R\J�oٔ�����+�����0��ٜ��d�#��?���P]k5��gܜB�_�<|Ʋ��co+m�l
�Ǚ�d�e%��n#5w�C�Vxt��TD�����r�Q���c^��KG�0�3�!V+㞍�?zM�J���=��&����Ҧ�Wء�v��L,�*ŲP�g�B��n@^j��Rf�J�&v����Im���"E�Pd�}R?ʫ�m(	��O�vy��Q^3�
��#S��MZ�|c���c;|gt@��&��+�pĥ�/T�2(� �X��B�6�,A��$�FX/(���l� \��'�-U� ��`<+�l{��?�f�;AR*�O\�v� G&�Vߣ9�C��>��u�ë�(ſAF�_�rwc4@�i��Hݷ0!�6l��գj�`t�N���9��%:��bo>d���w�Z�p�Fku-��'M�*���t ϟ�5�����GC"�Ĥ���
�N�e�Y���e�0��n�:L��y�2
W%��*1C����b[��7e!S�4B�fG�Sܷ�zkHf�s�3��/"����O\�a�����Ɲ�(�^m�[�a1�Ox� �Ζu�u��$��ހ�_0��N�V�(QG���e�������ct�_N�ȓ�z	:�~P����V��z?$�G��m�r#�����0��2s�]�-y�y� 1˚�� �V�a�&�n,e����*���w��� �G>z���ƻ�qST���!����_S`��î&\��c����<�t�:�����U��HO��cn��췵��_k�/��#�pig�������U^����`%o�{ʣ;0?):6{>���2q�$�x�Z̴��g��ϒG�"�{���z�G�3�wM�0ܞ�w;�z���pa�F+��o�V��A���>ֶ����7�*i��2?�|O:��\��h���������{H^p�wX�-��� {LR�L8@�����vo>Cdzy���#���	L-}y�($SN=���}�=E�k`m
3�KQ�<���uo�qAq;]���*_����t�6�{̓�C���9���4�LX[���^s��nd�v2G���P;5?�wh�7�| �֒q�i*�H�{M����Q��̱�_܊�F��U�=�(�4�FX��=ǉ2⣦?����V�������!jυ�t���f��BͩX�9S��R���b�������I�Z[�Qq��5}|D����������	%��d*�_��'��*�ȯE҈_��<>��8�Ǫ+�u� ����YX�?���cg��=�f�̏
���vu�o����&x,���!������gs� ;�~u�)�	�C��M��B���G�Ѵ��ƠY�L�v�0|l�Qޚ�Vs�ؑ���3�W#���I�<)_�f�������S	g0���TG">B�;��+�z�첼��50�Y�����כ��'Eq/���4{�U������uAA��
�ћ,�~3H� ��j��c��&��ٷ���1͜����o����M/7"*�<���ؼ
S��{���k�Q$l?�K�]�O��xɓ����+��i�$H�<�$M�6mJRB�;����wF#Qڇ�#A�����@�ݯ/�ǈ��;�-~��@u�����K\���|��M��L�v�eqOx��y��q�];n�]�H���:�z�
$*�^?��EO�Jn��_σ�B"�\Q�k�&�6���L�p�\�)x-핫�~�Z �v^hd	�gLl��8��{�x�c]�"��2v-�<�Z博������A�tl=��Lz*Kr�l�����"#<���t~1�b�����:�T�tlŹy�9��-����
����I.1}����s����H=L����׾�a���0/\� ���$x�R飩��v3>I�^,@�8���!-5����(�EU�2��O�΅D��� _V?Uo �/�`3��Y!��<HE(	I)iky�z:�nm�":��C͡Z���v�)�XD�ꮒ��+�����	^�^���|Dud��P�M�o�$�Zw֏�����n}�E�T?Q��+~Yc�bR�eVčh�=cN�c�#�ǘ��r��p�ӯ�m�'<#������eN����:��{lvWn;>��it��t��?7���3=�@{S��v:B��~�/a��o]��W�%8�DвS����i��-=��>&+���¦�<'���?Y��Ϣ)竴Xܐ��:ܐ c��7�H\T��<��{���i�(R��؁׏������	��n�?�CZ��F�Y����uv���X��Y�<��L��8�@�~V�^Ͱ�t'�w��e7�Ӈz�@EL|�^øH�$�J��Ʈ�.(\���ς��_d"�^�~��tʉX��(97�2T��r]ѝ�9���8�ƨƇ(��|�`�ZqZ2]e�Jkn.h��(���39�f*ߜg&h+�#�B�o*�ٻ��Z$7�k9�M�*o�?Z��YAL��[H5���G�n1^�d�X��
��D�k�8=�]�zC���b�Vgx	���2�ʞ�@eS�Ϗ6+Bݴ�-5��9�G�SC呍r��D��z�ze�s�G��M�W#�O8�|D"�!�%B��G��9�����T�����)�6�wn|
�a2�*)�����?g�@MT�H-�M�N=rě���2{!Z��j�����.�gB��<H`2��o�F�	|!�)����v~�S��Q�uQr���f7��{y���lqx�>	�K�D9���|�84#���n�G�)�T�_	H��HTqko�&�Œ{	8����FK���y�p&d�����F�#!E"市[�(,��T��G☵�U:һ���ޘ"��}�)>��u���t��c��E�R�IO� =7���-X�Z��?iէ���jKy�߱m#T.{�6��-R�~��m��8s�YO'�P�]Z�<(��3}L&c�lA:��ď�$IMα�k���<x{��vC�3˝ۥ�V����`�/RUS��1B���$!�7��a��x8Q-J�5w���3�Q�O��\�������5��H[��Q�N�>������!&�n���%ZS�����NC��:!�)6�r�����7��m?xA���b�M��_����\�G�G6�ׅ�cP�-=JE͟�Ge�0y؈�lj�Fs͇�w�r���Jr�;�7�����p���,0����{,?���B��p�>b�	��-@/��8�Lp#�����]P�ֹ_ɴ*���?Wvh�{�`��l�Ndb�P�L�9�>�;�41'C�����l,����[�)	��t�A3�2=y�.tx��(;T��L�q�2�@,ޟC�0r��2x����%�2�L��Q�)�/�:� ���2��#hy4��+�6�dFE{��Í���o��1�`>�<��� �e�H������;;1py7�wǞ�!^0��j���㣯���و��=�ke�%޼YR�E���5M�B��O�A��@_,��Ss]9R�(bVy1��,����n0���~���؜��Ĥ��zs����+g_��Y�d�h�(�|�9]�}��/ڲ�N�����3��l^P##� ��t�������=�t����w��2A���n��̨:?psv��x�e^�^'p/�F*�Ɖߩ��^��%i�hRRM�8�v�����-:��W�� a��u紽_��ڿS�I���X�<H��RW)`�%��D61���1܏���M�7mĮ�	��k/��ì#)|K0�HR'a�fr���
 g��UPȖ:�.%�(���lx��9P�P\�R
Qk�9�����&s��^"��@��@0��旹�Y��2��ڋ]�����]�vT���N����L�>^����hKy�ʋ�3�x~�?��
���g������_G%��pWz�D��-^��qSޞr�KQ��
ǅ7�X�[~��=�@sY.,C��V��2�t<�f��X*���Mtx�ip�ƣ�)ВH����p*��k�ό�A�6�z�r9�Nq�́yoG�L�t9o%�mA]E.e_�c<�T�'��G-�L��ߧ���0	���pW.+>fuͨ�sj�9Q�*�ܧ*r1Zz��J���vAS��_�?`�a*o�󃀘��[a�:��p$$:�J��^�p}�c�!N���K(�?e��ꩥ�tS,�����A�����ql2�L��d�e�+����G��^�D-b�B���΄{�^&`�Cn-�*�͇�A�Z�L�����bd[�F7偵��
Q�F�%v��+�/9���!�O��%9��~p�d�����۶T�h��a�*榧�|4��A��#]%;��2c�z~Չw��T	�TH�dCك�=�>��}[+g+}>(�3 .��}C���}�����( ��� ��VKܶ{w���^rH�tfb���P9�g�I�=�zLE��n@��\��y� .{D�.s��3���R2;�
 (cgD���*�If�#0�T�/L��6!��R�9��n�U�s�0f"SʸIn,t8�Wʞz����2͌�sr>�3�{�{�3�}�X2�"�*/��?i��֓��U�'��ȉ���������o�ܦ��W�4q����g&������5��+�_�GۄJ�	�9'*�^�qs�VW=���+�p�n���"?.Ub�㼟�����I|:��\ŒC�k���Xk�g�-����� ƛ)S!֘��J�7�	��:�A{�E� $4F��<簉&�Q�E7؜!�E���0ز�l�,Ť72��f��8q�x�
5&.������d@����b:7�� ���(q�ʖ�J0��dJ�'���������F+�G�@���a��nc���e
��fJ��I�F�r;s+:e-�(�խs�?	.�Y��8�!��d�FzƁ^�$6��t�:�qۤY�&&�/�jDrRVBa�T��E��Ѣ_-I��mUэȨ* �A���RE��V�8]�2����!DnVvI�;�K�yv��}�'=_��w�J��Ȃ:��X���^*�H�
�)1�u�b�]����(�����tt�b�a^i#~/�*�=)�X�<�/"U˔&y��4+��M�j9���!��p\�W�u�W�w��ĵ&��j�\c�{�KH�7%�s�:�-;��p��ڹN����Qqu����y�����{W��Z���4�/m���^�����[�o�z:�ƈ���k�/�xB��,G'9;,��_wU~��m%0�M�d8 ��i��z���f�A;t�И</ ��Ӊ^�)��V����b���%/<>�ͨ>�U���v��B���N�S���VY��ۨC�H��a��/��t|Op�$�T��,D\���{���#�R�g�2��+\�8�>L�S	_�<�Ԟ��2{�^�{j��*��W�T��4���x����h��_�+�G)�*Ak%P����w��<��Eզ*��J��8�]�|-�F�t%�8|�Mo
�:��KHg?Y��E�;�-���CY��EY�3�7,zY�c�3ĵߋ�p	I7����pQ2��c�N�d�Ѥ��87L��8�*G60�6	����)�u,ڇ�/w.(\�s`��%�x�	���{@�,O|B�ȶ�Lx¯*f�H�}�
Bf�T=����#%�6B����P
�D��{�Uɟ����TH�Q�Y�y�^��L7&���#���.���m��۳����@�ެT9����9_^���C��6|!�J�x%}��Np����4�)���u�r:�(.��$[
)i��!��$��q��RH�
���$�0^&�B�^��F���=Fvp-��4tW�Ͽ����A�V�с�49A�&5��3�j��ni�R���K�\��7�3y #�L �O����S�Y` �9������D���9����|
vGθ�V�l BL�7�@O�Y��4�8��wBňdZ����z�@�'L 5W�G,W���Ł�;w��Qj̬L��J�D�q��VC����2K�+Q����-�#�x$��i��]©u���
��1l�8/��z�&����Ʒ[�N��1w�1��3-�Zݡ�օ U�`X�yq��m���z��g�S���~~�F�X"��U�kn@@UY�����Nq�k���~��B�&}�s�s�B~����m�.7CD6�̀��$|"���.k���gB8��&��>�L�2�ڔ���U�O[k�����~L����i�W24٭�~����e(g�� ��&r]��ͮֆ���b`����ϸc���O1��[`J6[��Ɲ��Bbf^:U� ��}v���(e��� ��>q�����S�RFe�����&�6�~��՗�y��ە���i_�8AZ n�[��m�����Y�2�`ҋǅ P��a��h¬\�� w��l>���P0A=�ɢ�NW��{&��7�$1����jT���݂����|�j��'�-+;��t�/�&�#���U��4�F쇖��秜 M�}�9�?��r�� /G�^?ipԋ5�O��	����$3��/�ݐY~�籕��\0�D8��<��d���1�K&=�ޔM|Z�
�-�es/%j��������^���̮/�]���g�l� '�\������(����� L��=��\�)��j.U���	LEӀ�?R�aW��/��!������v	�Ä\�_�9�tTw^�*N6tg6a�,�[�����cu�Y3x���zʷ�(�Dƚm/1:��H��\3�j�қ}��tp�`�^Z����.?�<}H	s��	�x�@�$��i
X�V���{>������3�bW��z�(Й�T�Ͳ�h��^BLMk���h�+D\k᧸����|�إ�~%�I���
��۝�R����-޻����w�c9�f������	��*�)l�t�������u��﹂W�-�35�~��G��[]W��+�y�G+\�Q�f�j�;�<���^-��i��e9&�C�p�]|�*[od65}�m�t�F�HeS�Bn�%�^ތ����ێK����Gay��-��拏��<���g6?NK��;	g��+�j>6����<�=�����F���P��۪m����j�:�:�!���"b�#������N
�\��x=i&�n����3�������
;>VO�Pg��Y��5F(9J�Ub@]k1����In��������%+L�>n@���Qy0�mq穙���>�TWb�m���E��K(!�U*�l9y����ys��*�p�<��/�b&P(�$�Cz�����fu�^a ��wu\t;c�o%�K�7�����!��1X.�U�|?��/�M�[�^Oэ�!Vbd��//QgKP�		n��m�����k��R9�P�~��K�gH�b���!��2��lE�~�P�,;�0��� �RW\oҮ<ͯd�yњilq���~Q������I$�>]���0z�C���e�ഔ�}��VC�R���X����`q#ϛ�V�Y�<��p*"}�lP;�2e�J��I�A�pt�P.u�aO��}�!����Z��(��j)R���<p/�Y\�/6�xEKqoY-q��%�j=�jj��PȲ�y^#�18�xpW9zl����K�
�| ����_	�$��̯}	s/�Q���x
���װp�<O���K:�5�ݎ-���<�i�|�-���Q�jBKl��j~x�Ra��w�������~	K��F��6���}����q���W���+;p8��1"\��������c����v����y����M��\~�IM���^V�O��e���0��J��6�'�!�^O��G׏�1��	�^�d�t�sQd�Y`���X��� �l�[:�w�T�}���8G�rGV�c���r�~��/�w�?�vg0���!�J�!���ˠ���͇�S��ӑ�@�P�� sb8�!�oY`�b\�dK�J$�]߽	��w�R.jw�?�n��r�j�f�wOA��P��,"8k�6r�gާ,�CŏD�kGU��η
�]����[H��tx7K���J0X�C<#�Ef����)����sכ[;���}���R�a�ό�D7��A��Ut�szP/����"����4Rږ
ώ�m��<�ES6%��
�}7@�����>3��P�CX�VHr	wS�T
=�'&��B�C��+)^��'�v��C���H��&U��J�tD��E��\v���2<w��,�~a����:
)��tX�e2��7}�U�����8�/e���|�Oٶ$NZ��/y��%
���5tr\�:��hm�Ky���:�#Y��n]������~�F�|�^�b��^��S���ۉ2��m�6�TY�+v!�"}�a(tc[}�O�ׂ������jb~� �2|+O3���c+��>*����!7\)�/c�I�a�^�ۊ�IX,��'�kzj#~!U�R#�0i-�N�'���q��o͟�ES�".09z��'��Ą��@�	&�p7pQ7�������)��%���z%e�bܟ�cd�l�:g���%�����ݭ5kt��?�r�� L�����zL���Y���K�/w �e����c:�D/jks.����股��l$F�\��e�����Z�Jx���5����b��was�֙ض��O|u��]X,@
�a}KD_����T�=a����#�YV�*�����fH���6�jZݺ�� �<��T��흎���.�{�{�]���a��j��qL�ʖE�M�8��{�/r\���;�̔��j����y�}qʴkv���'�7��=��k��A!󕺕�{��<H�V�Z4(�J�vV��M��7E�T��^��i�T�[-ӐJ�9	���f���[-��XH��	i�s>>_T䃈A&�O���`�.kj��Te4O1-* ��)HDL��>wp���;�B�=+�+��3�Of ���طh��\�!�
�E��o�tB�Z�2�c�P�/�L���X��<8/H����e��*@�pdõ�Vo&t_O[IsR�i��3��l��w��2O۱�_�N���O1jB]�{�m9������+�3Q?��|��>��6�+S�d�ś�.A���	�υ�v~������,9�Ge(w�/��"ò<�[�o�'R�_vϻ�� �^CS%�2��pG����tTA� 	1u�F�gA� �H�h� %21fo�;���pM���]�Υ+��5Tڻ:�&�b�C\��WѪV�*��r��w2#�O]R�̃|����_�mUM�L���W��MW:~��m؆����'i�gq2e(OlU�$�Q����z��/�>��5���l����2��8DW�M��H��B]���Ͽ��;�T�o�cp�饤v	���H6ӏ��7�Ʉo���z�WO��%'j�1x�o�{���B��``�:B�;�Q����e }o�bĞ�P#�����I�ot�*�������}"�N�� ɬL;50���oD�[��s.�Yq	.ĥ���YQxR0�Ϯ3y�} ��LNQf坦�s���>ҙ	�ٮ���/�)L�F�+���o�N�T�;h�+�����dYU3�5U�ݍ��WxJU�A�T^�\L��*Y}{,�f�Ë�������Uʜ�2��%��I���w��.G]��:�@V+*C�zI�9i|o�m~=
�<"h\�J������S��ݷ>C4H��I�4�6���~�G؝�K�:��I�]�f�}?��c6��F�g����y���tа�z�닶��A�8.�3.�>��&W�d,���9<Qg�̍��{�~ľ��
	n�~G�e�2�� Q{.Q4{��( �a�'��
�O�(��D��.��T����/����J8r��퟽�J[��5iɌ���]6Z��)�W#��q�Q��5�VU� ���˧?*�eC)cS���08Ra�MQʹ�~�7�)r��]Κ�r[}:b�j���uypR��U����蕯��޳ n��#��bZ~�=�I��j|0h�$���/qu�m�_ +I(�sh̢:�Īs������e?󐲅@:뭪?�x�Y����<q�1�s��;+gxcp��� 0h��Oi�l�@O�N�b��H���S�I7��PPZ�(�����g��r�N�n����L��v��x�v��d\���S�2P�a���j=W���<�L������
��N���(iM�
�`���B�Ъ��L΃g#�4� �eߤ��+<x\���X���5`�Q;>3,��2����;��T����IIV�	� ��S��gCXaz�4P��
��t.�Q�)�����j�R�[6\0T�¦L2�����r�-����J�X��j��o��Uq��O��i�5�Z�<�h��l!���%W��ì;9�y��DNe��B
�N��$��EW�[��CU�g莤�A@��*��p�8��ydک����nS�ϥ��%��&9�k�t�W 5��Xw����A1V7P���41{�'"��葢l�$ ?fJ�a0/�rw��7A�|s(y?�/�l4rTS�>_���@�s��S��"��q![�H�`�0NC����;�U}#��PЃp߷GHA%jG=Y�;<�	��"C����F`�f�y᫈e��>`3hVT}?��[e�Z��K�:nF�(,;�pM^�P�#�����\��<�"Y�e+�^.T�SNv���Ñ��7�|�V�����{�86��!����$��un�n0�lk9���w�e�gÏSzދ�r[�Jrzzlǘ6�!O��t�����Ȏ���@����9391���}�KЛt�}�'��?�,qq���
6���R1���0���q$��ыF�̐��]P�������PBs�/;����:���*�J�2�#/�$�˦��M�������X�4�G����,*���_/M�[7
�B�>8���+d�E#�,7u�N&��i�,�:�t�IQf�n��tk��"�o ~�BZ E�ų�R0�c���d%�v|��a���/�Y��4}B"�G��R\�,��_�M�v+��U����^���P�l3�]���O�?,W��ʖc|Y|�>�x�Y{/�,���||�� �Ʀ�ٰYsrO���[e���[�� %��;2VO+��L�I����{���*�-��
�m�c�'Ϙ⮋�t�(@��%h�`z[ ��f�h�}��@�@	ӓ=�&{~B��\��Ɍ��ke�z\Gv&Ý�nf�ݎI/�a��s6c�`�T��
?Az��4�m)�F59}�-<�D����M�ᭆ���:;��?��p�@T�_����$�&��BQKdh���*��֧�l���A�������W�l�،t���_\Aw�"%͙��"���9l�\\�הq��)� �V��ً&��;A��'c��� .�0 r�N��%�·�Y@,]J��?öHw{��H���:;FZ����	�y��R��"q!Q���)����2�i�%`+����J-u�Q͸<bRVOҳ@e\��3�����vm���;!�%�I3j��f���=�v��3J�P%�Bj@��ݑ��w����쐌�:��@�	�X���gyC'�kIR4� ?����X@����	9Q����s\�՘�ar&�1�����P8�Y�l���kz��ynF�Pp�^kM��1���"z�ŭ���<b���&p!�V�<��t�	�?8���@T�+Y���`$aL��\e� ��%d@�x�O(c���k"�Y?��ߞB(j�r\!�h� �9�L�(8I�̩����PM��v�zD�����A�lw��GX�U�THñ��S��wn���Y��{(���K
�κ�;��V���>�S���M���4\�eT�"�}�y?)�u�\��=��B.,����)��qס:��o͍@9�x��g�ӆG���1D�Z����t��Q����9��r��%�}��Sq�u.N��� ���,�&����@I���Xs$�}���3��4��m���_�0�C��5����4\�L��z�0�e�ѐ�h�I	�}��Q�b��侷2Р	��p�!@XM���Đ��L�,��O}%ą�B�Vd���	}U/�Ù~��^f2�����Mml��IA��\KY ����������xIp#���{C��x4YY��x�+�#�mۯ�6�x���L��A,p����l驽��d�mXvU>q��`aܒ��"1�t�A�n���D"!{��d)@��K$Q38w����?4��Ǻl��RG�z;�t�J��õx�qCo�MO�x*	���u�7����6���|��X/�3��Xc��f���x{��=%�Ū.��](��S�q�������譕'�/<��5p�����pn�M����V=X&��e�K{+Z_�"0�������S�`�45�o�-�Ҡ0�<���u��=@�䧴Zݨ��o��Hi�r,t�3LL,mzι�f�	��7+'�wyN��Ǖ�j�83<ږ�6�!����5��
�5�@ڬ��NX��ւ�-��i�����m��#��k��4'Ȩέ5v�گ%�b���D��q�9Gq��ovR?�s@���g��Q���QH�
]�C�s.B-�+׃��FT+A#k��.�d�p�����`�l�$���i��G��o��WM<�㣷v�`3�����[w[+)�<��Xi]wC��U�4���<H�2�ཱ�����DW|��__Q-ܸz���W�R�7��i�g��@H*��6�>D6�x���N�5��U�-������.��uf�:��H���5��l�������G��|���ְpYўuN�,{�|���se���``m�(*C]̩-��ì��LJ^�v/D5�7���7D�2�=v=��.�0�~冫ݺ�+W��<!��e��͗�L�'�E|V��6��*�b�+�����/x��<�	�[��i�[��fd˺�D����W������Djѐ~�r}b�������	R���3{5�y-0x9���p����(��t�{��r
��Yo9Y����,�Ȟv?�к��yVU�m-BQs�	��U �;w����	�k�������dg�E"q�M�qs���ҞPs���V�یS��Y@��A�ʂ!��p�1�����8p?��PӧIiU��EN��#���-	��l���S?+1O�Օ3iڳ��F1t/6yŒK��"�mx��M�B�Ǐ'2�[5��8�I�K��_گe��p .mM�dc�ՠW��$�t��ĝ�Qz��ϡs@��H�&�-��9>|��
����nϟZ ���A�@A�IT�~�Վ5f{�5��[k��Sos�..zs.H�#-6=�\���>�%g�*B�u�?�2W(��I>W1f,�Po+Ou����C}a�gq�	Y?+6������N�z��^�h����q>�l*����R5�c��@P�	 ���Uv���EW³��I�!��4�'ԙ1n���ʈ,'V�A12@Z��ip���
n7l�u��b9�g�f�+�n�5E�c�
w$^C��2ݛ���N]l���'���9���b�J�����v���������מ��LE��V�@��آi\�Zc��j����~h�Mj��5x�CE��b��aL�{�I>�o䪯	�N�l�F�ߩ8������!��>'xN2� �bq�{[ h[�>�|����0�/��K�[�y ��Q[&�%UJ���P�R8�=k<�����S�y;��m"9p7��ߎJOBx#B�B������2!�A��G��i��a� C[��io��",�q�����2���M���BeF����a��I�v��c�Ӻ%U�#)��Z�o���{ew��sY�����t��0��u�w��c�rG��8]�憳���AGMnf�r�uG��M]v����e%�FM��H<�K��c���#@�5����aK��{�F������M,�u��:����с�9Z�%g%<[
�Z"IAY�goD�g��j�:hn�|�ܿu��H�?�lf�	���Aw�I�>0�a�BL5�R��娲MyC)HI����%����d�A��;0�D�m+��̏��bc�wXl^8�9ZK�(fvC�X�Bţ�Ƨ(TE������Q�3f��Y��q�)Y�Z
$�)y�n���B�w���-��#�D�#ma}���!�8�[��ʝh�:��<�Qҿ�B}A�5H9<K�oV����bE���i���g���5U֌ݷ�+�ɰn�@w��m:��cJ�rv�A�P�IB�{�0���
Zb���A�x��m�F!�*�!��3b��=��s�\O��հ�3��Y�}sTMS�~�6D���)}�������Aw"���K�����呎ց����Es�Hp�>�Ɨ�nB6g.��A~~l1G���*�4I�uG����[r��.��)[$L��'���\�Ļ����=�(�gfz5!	��15�2w8*���9��IGx>�8p���醞(���	��T����ӠO��`dǷ�0��E ��16�Y�h8�2�"��?c����m�O��6gAQV�`�;=�םÙ=*"�����E�﷍�`���-�b�G��TU�PU+��9t���z�o�f�`�v쥩s�'/g����֭ 5<���|5]�=���O��O/�.R%�Z��l�?VQ�������\��Z�9R0�L�b�R@��	�Sq3d]�JMU���DA������ ��S�E[3)����R���~�V6Zv~���3B���4 ��b��5؉A\�I���h4�3�O�i��c0���X�LFN��u�t	V�KfC@�D�4�����n�ݡ'��'v���N�OZ�&gb�;�W�92|+�h֗�XR�E�[/t�� ��f�;�)��1��)o�y]��򅢓$ฯ�G@t��h�@�B���gݳ��d̺�Hz��"EcŻ�_��Br��ԉ��\W�z)J`:b���]� @���=��mU���m�:_i�ؿE:5�CW!��{������2�S\j�.Np���<�MJ�\�8�oct\F	�ʪ'F������K�&�-p�,�rff�3�y�X��]y�9�<	��!�}�t�<b%~��{�G3F���'4@3-�_�ct]��O^iF���:<�$�㤴�'wr�K,����B�E+�����cş�|��)3�X���y{��(a֏��K/W�H� x�-1IMc+*���ړ:��M���`�O'N�pp`FU�=��8`Cs���@��p
��ǖG~���;�t�h�xMn0�ׂ��nw�x�6���c��)�N�A�)B	���`��<�oލ�Z��) �6�C3��U���J}�3�J�?�b��d��׊kcp��B�6�RϧN.O����� �I�����."�^�7.�n�L�+9�y��b�e�|_%�`�ZY%��X@��i�Z+�N!*wSo8��(j�E7DO&���}���$jոR����,n��IT�uP���K��x�w. aXg��X�EM7��}���i-���OwF���;��e;�1!�َBIA��:�]�|�Q�z�������M"R6y�]DE��x��i�W�,�����""ݾ��JA�#���H;�����+yo����ɿ1�K����bVHZ[5��熈�#���RV���019�S.N4�����tK�·����Q(��8���0�ܸ��a�  ��8]t���fp�[2-d��W��)qnP<=��ڃ�ڲ,\4xޜ9
�P)��ء(�Wg�	\�4����Dd����ưLă�
}qI��z'G��y���d(�B�pi��~����0�*st�#f����J��D����L�'�����t��v��Ҽ8k�x"�2��lc8�������늒40A�Am��Y��,Rz��p��fm��.�'I��}���m�2�{�f�a��?L#h�4ה"��.�&o�h�������d��1��Wq��\rM��-�A������f�o|C�Ò܍˰7U�}�QW�hm��g���l ����au�(�2�-����q��X�T�4��4e�$"�����3����YX� t:T��7<*�bU%K9��ek(��1;�!���C5
�b,qƘhCǎ��ׯ�bfI��#0�����`��n�|����a9��3xf��llv2�EN~xa3�}o�ɬ��ts��/��`�M�N��G�e�����@����c4��#������͔n��ك���W�ŷ3��� y��OdVo�ʿ��.�D��O>h��R����x�P���	�7��8�d"{S���=C�Myk���Ȟ��H͚8nFL��J.�+����BO�8hK��;-m8���քK)o�!��TR�t�>;غ�W�VE�F�:��b>cfh��;��*t���Du����*��z���6���Hb�1Gk���f(�I{�l�
���z)���2[��A�Y�J�!���O�bz�u��	���J,�QE�j;�1�Q� ����ǡ��RګQ�˶y^�������=����t����hU~���Rsr�u�Yd��b�1�Z��7��I�iS��IO��,�b��)�"v�6�6ͱ��VUp���$��R�cI&�~�w��!r��F84�tZ=�����R\����|�FK��H��˦ݷ�[�1�aA�
�m�� ~�@�ʆ��ʩ�v���ZEU�5@�p���9(�v!*�u���)���ii=�+GF�؂��u=%�Qн {!� �M�"�Y<d �q4Y��=��;Ϗ����vw�?�͂��,Q��5�=8�Ғ�7�e5��Mx���[u�^��݆�k%)�F�����?ܣ���L�Wpq"Z��M����������D�x��M����GRm����ԫ�R��Ȁmؗ"_bCu{3ڔ�g
Pܲ�U� ���m�3�ef5��^�曹������l���p�T��ǯ�Ћ�c�,�b<|�Fc���Λ;R�t��Ʒr�4[�k"��fV(��������ep�nH��R+)�ѣ�uP{6��0d�+�rfX�n�L6V�cUٳ��*���\�Nͯ�ɍ�@�d�M�Wdg��r��.$�%	|�� K��C�t��;'G˺���A\��Ď��b9~4�S%�v�j)nB��=����ш)���/�' ��봅Ru���{������ @Pz��ݔ&�zb8v�'2�L�<��B�5E�P��̅��\^���x`eRf��YYަ�߽��fw��S*W)�ȟT�u���L���on�z6.{uY0Ǵ��q�)	5љ)�d�<�)�C��F(V{GB�$"��֤����x��?V�O�ZdLL�z�aSi��lz��͝ҘRf5\j~v}�����X��+��Y���<̿��UUX,�͵/y�В�c�������o��}�^��ߛ*a
���B�Q���U�"V�_�ϝ�v���I~�mnF<>"��H�Vh�?s(�x"�� ����T\mL(�?(_[ݤ\���5���T�|Z+v�1��]�"�=�gm�-ԊV��)"��b+����1���bWj���ޫ����8��E�G���(��I��!�d\�l�	ևIO"�:��5(�WW�Ow�7�굠g^�w���,�!��F`0NP�ǩ��߱4�.\}����*:����B�`�^n�dU�\�<�X�C�%\�[rޭ�����ٔ�8�U�h h�9l.�� ��x^yyY�"�Tf�p���Z+Z��z���W�m7ܖ�B�h�Y��
v�3Xc��N��:�B���*e՘`�^�Jrq�KL���	��q�)]��/cEC��'=�B4�������[�:���IY"�b�|�4��8#�|+9�-�D���]MMO^�P���m���^g�Q�G�ގ�3J_�N��
-MJ1��c������B�I�~�D��]��gB��(��	��vx�g%�2���vצ�ObE��F��X�Y���*�c�fv9'�D�Y�M�ktr�����^{�EY�Y�E���5<
M�f�)�vM�ࠔT"���Q���Yo��A�zip!pZj���~�}%��+d�#���]��Ts�#��-I
Y���o��9-%��5<7���
z�O++�,˨�ύ��Z���K�Y�qS�wEk��`G0������K����F
f��}�����X�Bj�7���R[�i��ې��eɼs�򔁜X|�wW+�e���pD̩��uLV��~����Q?l�g%?�qXF��ӧ7b��i���� <���E'�?�T�n�ɀ�ܵ���N��R]� ��,��#v~$A\�-��되-��''A�[�y���u%it���|�@۷h|�qS�a���F�(���r�Kv���?>�;Y�I����]�s���6G'/KK:<5I�T޿z��uc^�p�H��lƵNoz\���=^���]����*w���j��X�;пnS{n�,%v�:q̨�<��8�<]�������Be��䮽��_��)l�Ü�C��>ϰ��U�:�,�<<�
�y�a� �&w	�6�?�r���g�A&Hb��F�ǎ�=\
�Z�*���m�o�_�Ř����|9�\�D���YR$l��9N�v1�o.ՔB�l������:;�jht�i���Z�r~R�ǎ!Z���H\0��g��m��bOhGbG������-e�|D-'��nBϫ��~#�[�?�1�KVѴ���\���N���ӺD�7(Y�D8uk;�Oճ!
�� �\�B��R8��3ǵ�nT:L�*�F�e��i��9||s7�˶�Ox����&�9U�� �J�q+B���	2l�$�s;�[cc�LJ���6&�_t��x���a*��1�����BK�+������d
Ԯ��@=[�लm͎j���?���Ƹβ*��uz�ˎP�m#X�Q��8�K�^�n��mZ��4le ��i�z~��$�,�iU���C�bu��+k"�dEcGF.K��ǝ�vL�?��{�ݛ�Q�9��.��o��b06�np1p��r�"V�7暒Y�-����i���u���)d�vJ��]�aiUHY�&t''����\쫟/���6q���a��W7M+u���=�_�d1&��՞׋S�����뵅�6eۍ���Q���8F.��,�Ҥuw���j7O��+�V��y�U��n��KP��L� Q�8T1vǖ���F��?��P���Uxĳ^~�0��(��̟�7Q~[c��S�`u�!c1��S�\�����kE��z�ꃁ0�8գV'����W(���a)N��0G��dԡ���������$�1oX��[��d0b T&T�[��H��̘813[�O�
�n_Q>�Ɨa�+�,iMM�J��G���Ե�����8/\��2�m"��â�ĩ��K�ԢF?�Q- �t��Ra=��ֹk�l�6��!u���9�*D�q?���B�V'Щ5�#j�"AgZ��^-�����
 .�?uoH�[�1\W�w#�1���f�tB��$mr�]��>nn��O��_8�03�:0�[�s��Dw�'�9Y�7][S0�����n3�`8��n:�����+��ĸ�Jm,�H������&�<��|�V�@,sV��y��C��P�+��jÊHlD'�v���4��Nɽ�UK���>P��`��z�
�⏘?������+�Y����1=����'X͊D%�3���'C�@i�G�5�㭒k�5�����:^�����-n�����@�,�b���P�S���ҫ���<�	��iBŪ=���O*�o�U8|B6`���oe�T��4:b��p�x�1�׹Y-o�a[��� �m��5R����@g�mv�/���1��5��a�B����	�{�{#�$$#�p�F��#��|���^�_B��::Բ1�p�3�Lv�h�`D�ɇ�^q�5�ay�IP
����|jh���%��g�y2�D*�Xc����!*Tx��w1���[Iz�e�Ww�3�l��&���R����T��B(%� w���ǃ���j�?` ��^A@n�~�v�~l�>:I(�94�>���AW��J�ɕ�Ou�Q�����H�[��N��V��x��'u
�Tvxƈ�	L���_�Ua��y�Ȱ=�<�%_�X�7�˜"�ߐ�{+4�~?�9��r	z���C�?ʴ���e�QS�"'�h��4N��w=t�+��M��:	L���%��;Ϫ�#��rԥ�|ǽ����I�wіh��	��C��V���9�	p� Z��Fú����p%��/rv���2Ჟ�=4l�7��\�(����ֈ�y�(=��T�����!��xW&�FcRx�RR*�]���Q��$tf6�@e6*D�n�����h1�t#?�X�h�fy_��g_5��]�1�f�p��;!�!��0:�-�k����8iP.j�)r�:�Z�Ȉ��u+�2ћڽ�n�H�2�{�>��m�ZQt��D��/���N�ݮ�^��.L]>�t8P��q� 	���4z1��E�|֪H���	2}7�,�̦��J�*��[�޴�� �4+�9�@�;�!	H��::��_�eT鉸w:�g�?�3Twt�)�)ЌTP���DRl��=��:��<C�" N�^������{V�q�um?��+Ӵy��Ұ+OY��J�?�4�y�T���,mH��ٜԦo��\OTj�E�Pp��f|�C�ݤ�+]f0G�� ��G�j�'�}h�%m�7D�({tg@�Y�d�����ѡ&b��Ƹ8��4(pO�������I�:'Cg�!׶���[J�VN��=���UM;BT���̽YM*�T%�8�?���f�J1r���ͦ�(�;b��o�-�+^*�K�ߒ�����0Q�����$���UV��[�y59/��ۇG,
������`uftg���(`��8�È� �w�;��}��Ơ͛��$V>l+��p OQ��nώAC�S0��8������z��6��a������ϼ�o1/T�+�

Wv��z$`6�C	����3 �K"�E�y3W��#��gE>��$5	��5�`�m�Sd򼖩�  �qV�/�Tb<�q?���e��~�~���b(OLa���j�c�.��h�lin���Y� �mxۙ�t�&��y��!l�����س�/��gS��G�0�Tv�ڙʾ)~sL���Ź{���\i[LZLe��/�����͵5���;
M85�����ղ�j&�m�=�;��zDE���R�=���gn��{ ��������4�X��P��$O���h>�aK�F�p�%I�D.��Xً������J�.V� ,�W��5p���!��^�d�Z��>�Y\0��ٔ��}Ʋ����/b�L�A٠�ӡ�C_0`im�9����2+Omc�hzaF;G�?+㷴��?����'�z����J��7�����t�7<��S��)�����7���vxA�B�~W�Fq��ڜ�5ْ�:D�H0	��i�5�����cD�>w2�z����/1�p�_nt�,
��d�j���P_�	�Z:�~�QA�-z��/ovy�p�3�n����
�7�o�G~[4je��yP�}�����jn�hR.� ���ᬔ���^��ao�
���N	EK%/��~��m~d��q��j�|Gm:�M<�MBoN�A{�.���}�Xªfß�ݧ�^��$�����i�6�̝Q�c����tn�
k ���ew����D�|���5s�F�R�i
�yXc}��E�-�LEI�;n9˴ |!��/Z�-�g�ݜ(H9v����p��?C�$�c<��dL�L5_���p���y�t�<,@� �96%$4u�,fEO��6�5��*E,��ȭB�$\�m���{�]Ջ+�,m[ps���W�1��C�Zf���\+QK:�4g��gA*������1���N.�}��T�F�3�YgP=�	*��y!��D<�����7yS4�� z�9p-���`�r�*�T6@�i�_��Q�	`�d���
"�r0��L��.g���l��vSm���(Z8c��մ��S��:�~�=��%�T�s� Y�!�DA�5mS���5[��#u�BD�ů6ݻ��Hɑ�~��-�cٹ�����8����U��V���4ȫh��91f/T"�e�*p]�ݵ�QV�~�Q+��:]��[�(�5���(w�{T�s�6M��0�}A��!���&� 6��;�}JD6G��.�+��.�%3b`Bs� �k�fN��rG�{VZ�"W���[�Ĵ��G�u�0�9p%3�6;l���
۾�A����<(�����-Θe6��Kl���"of���Sz�)E���KƠ�~���N�6�Sh/2��\D��/i�����(BY���N�)<ͮe&`>S���/��/V�� ���:ZM�/�"�$�2����J �O!-��ȉ�;~��J-R9�|�����#F^	r"�F$6�8�`G�ґ���4���Q�A��I~��+�t���;�� \,�@T7(d:��RMZ`�t){g(���e���f�l�U�Y��t����]$1���+��LrI2 �I��WfYn�n��=�ԏ�u��fY9�D�>�Ց}����D��8�/%`�� �՟�z�
�)���Z��L��U�4����h`�	:��r<�⟥~q� Gw�(o{.N3�9Z& ��S[����e=5�\��)~PN���C�abdJ��2d4�7��U�K���Us;�zy�&���r�j��/��d��w"}�l�����3�u�Z�hdj!�[��qʄ{�&g�wDz]YvZU��0Y	��8�D�V.	����|����{��V����T'��A������fgA:]���`VU�|�*_$u�`#�>a��uX&t��-��N���� !30#g���8�)��(���6m�\Z�հ��A�e�R�������%D\NA � ƍ��+��/�vz�!�������U�ᤞ8�X 8�C��'�7�5��u�(�"	��&���q.��?K1V��2�K$Y(U��O�y�cJ3	��64�,kx��;����${=�z ��w�ڤ�	��p���A�qWJ"�Pb��д��u���Ag=��7�,|9&�����5�A��2�S�<��Z��O�0N�.�M�W�:���k�z��}�VX5�z���M>���Vb�|}��m��c�^�5�׆��{��`I
Q�D+�v"�~Bu`[>��½���AvH�o����0�������Җq��W]��~1�
�d���u9m���z@tD `�DɌ��ӤӅ�~�5�Lq,aC�"��͗�P�,M�cyAO��i�?H]��c�0� ��λ������v�i�\#W]U��H�?VǶy�������8�/�!sn$�6^L8,e�1�l��//: �!1��*&4���g<�2# �`<�ʿS��O�1c���ow���P~u������~�C��w)j��n�6y���u(>�Al&�ƴ�,���i#�9_�vpp�`�F����U�MP���6ƴ��\��3�-�I�y5�0��6��<$0&��}>�+��U_=bcr_c�_V�EooR�R���*�._ײHV�5�"y�̄�H����~�.Na�x?q`��NA3�%0�D����וǺA�J�IҮ+��XO'1+���-���eMz����2��a�i��s���0-��,����ςY}�(�O|�'��N�'��\#6��(#	�(�kc+�a�l�8P�oX��dcƖ���|6{Ǻ�ِ��S:'dl16`q-�&�yWZE|[�1A�V���k��4�u='磦ZN�7�c�6F?��S��^
�ܝ)����2J5"_ok>e���{��X0�R�h��i�$�������_�u�D�A��o`�[V�����=l��G�@�^��a��5���Jۈ���.o�H�8wzi�׶R���j~:�����50�}+���cs���+g��-o}
H�8�ސ��(.�a_{���L���e��.�-L'��?��E��g.���q��=���H���k�^z����J�:��q"�w�{#�������a�m}����!1���=<蠂���Um�(��0n����'�2vh��Ғb9%w�m�ߘ��N�Q�0#� ��ݺA@X�RJ�����5�nWIۙ��g����?����.m�����|lp2nx�(�B�[a�;s2�7VC|���H�9�T�S�?nh��+j+�gڵ,����J��殥�6�X�G-i$L��x;��N.� ���i P[|���D���d�!����%��P����{T� ٮ�u��K�$�O89	TH�3�oWpP�\!�t�Y�5'(u[�fD%'*~���΢f}}��-�&f|��|T	}�?@�?^��,�]l�D�	ԅ��h?$k"�F"�=#�(
'V\|�@M���q�i�)e[�{;��yT�#P*+8�\���$��x�.R�/�� `�:|u|�ҷ��W�Y��޹�5��vcP����	 ���}��c-W��+�=kp͠����0K\�9��OͨV#87<v��[S�|)��!���e�XӋv��B4n���7���^_��{�!)(����h�dw=\S)M1���i���ydĂ�ig`���0�pB�[�S{0���6������o��Pd=(�m�~�0�ﾌaU#O@Rk������ǉ�o@iJ(�hӖ�(�[E�O�=�<	�<��d�����V����4Q���%4�#`JJy8r��c��C��66S��? '�14|!�z�墰�,KB&]s��p�$����U�{��Ҫ�Ć�������M�u������J�:64jJ����������D���u���X4d�C���f�#�����~ڇZQ�
��mR����z �����f���<��Xcs4u��p�#LU�FZ7��w<��k��Re��/��:�@��t���w�>"c@�㶇&IpNoKp�w�g�*Ha���֨< ����������U5�Im;�ܧF�ۣ��ø��'����Ъ�w�����AF��X� D�;�4l7����6�c����E�I=mC:�x;��}c0����;P�l����S�H�{�b�,�	!#�G���m�aX3$_�9��9��+�"��#�+��y�9P���S);�Θn�������@L���fТ##ײ���|"���Y��C9����j��ت�ζ��$[�K<F�٤[#�Ac�0��k�x�B6�<��ap�<���vfELٰL@B��]L�v{r�A�e��;�&�nn)��`Z�
7uŪ�Շ�aB3��#f���Aށccr+�U�r�/����Du>$8�e��k�NBR��X��A&qgr��i��߹g۶]��5�Z� ���$�-ir5��Wޔ���h�~���.s�ɧ�p����l1B2�z�	�@�dd���m��(��J��j�c}�6�g{
�H�ӭ0 {Vc!U҇��)��Q���9���RgBJ���'�D[<V����~z�UΕ;#�Q٦��f� ���������V��F�$xr���ɔvqui��,�]�)�c��G���3�%���d��w���Ԍj*!��a�*p`e����A��h$��������HT���1�ᤙ���8U����2v�a�̟a:X��_��y�.��7XB�_CY&g���D@1%3w��-�ǌ� _�HK7��z�-�9�ā�h{dYz�g�+z��3��#��b��r`j�C`�1���q&�" }LO~��)���x��o�N;c���j=��@Ä,�?�٢���V1�F��zw������򼈎"�u��F� ɤ��]˗z��O��+w ����Q�7�v��U�6ԅٍ0���9��N����>�|�p9��7�'�{<ǡ��>�c��z�'%�<�2^3s�a+:�Br��	?Μ�߱Qy�nL�$l;{��q��S�;�R������BDD�*|�t���W�ǘ7�^�IN�J�F��}�@د�\�A&#v[un�dSr�0��[N�|��+b�2e?�!j��uV7hD���}��ҫ�+Y�3�, g��"u��Ҹ!��m��M�M:�'�Ƞ�Uq�E����m��g�<�ɿ/�p������3h����>��Q1��#s#��yⳍ�rz�LWh��^��{��y@P.�*|�]։�@��e?<4��藲�	�k��ĚQ����tmn�� �E�����.����κ��~�ww�CS���t��U�<��d�aQ�
�oI�����,@׈�R���������&�ݣ\M���U�.?����\�TTx���Md��Y� twȌ�}�Jr�G��ܫ�<b����Ky/�p����	����P�F��	�R��y�uRd,ʇ���MR��i3�����pզ���w��n��Tu��P�d(��X��C:�Ɲ���%Eu�"���Ǒ��;�<�� 4�-�<����$d��T��B_��gކ'0`3/bZZY;y��H��(.��<�	6��/UL�v�.�}c��>e���n�y���=	�	TZ:��F%s��C��gI�CW 19��{�Z�,	3��T<�@tk������Cz�|t��<�J�k����0Cɏ���L}*6:����5���iQ}�;��mrΑ��u���a�z��R��p�JB�e9��u�Md�^2eW����,#�q�@��F�v@a'�y/. w쾨���#5��/����F�*`#�0��률�j�L&6gI��E�t�S̟�j\�y�S�q��f�/��`Ÿ�����]l.�&Y(*��l�K�'5;�K@b���Q�t-�����6]f��:�����}K�!�r+�2������\1S2�.��h�vuހ�͕º$C�Dm�J
$܉�mCyd�.
=�kc U��nF;�*�1�2�
d�K~�Ø����jj���g��d�r�>[K�QGx{�i�و
�Yx0"n������vQv6>�gp#�<O��E8�RdG��j�\'Ú�!u n��"�o�ڙ�/�o�^���|�*>�7��!OG��6�Vv�Κs����^Ր­�g�yhfN	f��(��Rp�Ń]s�t�pBG����b:U{HD6٨�~�-�dm���sV���}B�$Y�W>���Z��E�^�:��ftpn���ş�"��^F�c%�fF����z�������$\�c���~.�q����И=L���`�|Ҩ9_�7�/gӷOd)oU��kw�}<�� ��{�g�h��3gC��֛(�lsWt�')5O��1�ob��~�R�G)9`��e@S����m�bѤq�O�]����j���gzU�2>��79�W�Ȓ%��2���e�o'��>��{��r�S��y�X��=�Nh�����$�S�Qn#N�e ���#9����b�ӓ����nJA6�����
#�,��H	�[������2mqO
�Ƹns� ���S�
t�����0�m��ԑ�;�ҹt5Ę�T�1��Eڙ��r�����L���B;��a�g{�cFp�e{�������IU6w�GC��X��������L��X������tQ�ދԆH3�d��/�y�|��TJBFo�9�є/���q���
�uA(���F"��5Qi[�~�-��v���+��7�dH&~�!� 	�Rul�	�f��Ų����!C�z�����U���O`��x]W2�(���.�]E|��L�k����y�����/�§����I��ݣ�	�^�q�1Ge�_�<Dv�ę��	�C�q�dL��>�̸>�!��J�j�n�-4@��e��Q��=�MdZ.��T�J2���8X�m�/+�sc�s�$p<Q�I ��K:�p_A��RT�x���Tff���������@U���NvMc�e���WY�$���	�^k�[�[����ͮm~D�t�?�@��bk�*&C�nC�?������+c���go���zf������uw�כ�ɳ�lE�#����F:ȥ���%�>���Y8�l�ͻNP,:1�����X"��*FBj�s��ʭ~����8ޯ�h R7�a�#����l�"�B;���yW7��[	���m?CC�N`��§BY|�O�!f�K��1��7���?ϝ߭Y�س��{��V���4��# X);� ��aD��0F�[�[�<�q 6Y����D���>��6�>0b�AH�F��M1%j��/��4f_��������'���L�u�RЩK���	-�AʸC>���b�DxҢ�� j�;�y�{�y�*�矮Y�I�3�Vd�{�tM.}��$�mwL�o��Ջ�nǦ���;h8��ܱ���������{��MX�zٱ)����Y�z���g壪�HL:���B�O�,�m�f��"H�\P�{���2��b>��&M��m�z��7��d;P����!�c�4q-�Gh_�'�����@�Vd��Z-�����^Uk�?#�`��}c���#�<��0�r*��8 .Q8�����*�4S�����(:4.uQ׋q��K�D.l�`��רP��Mi�*yH�a70ٸ�<���Hӷ���t�ZQR,��|����ڧ��g6��N�(3�Xء�w!m�ꂈ0W��rT�rNV�t�I��n�C��c%���o]6d�<�#5#AJ9�,�l����S��"�ܮ����CB����}����c(�>�4�K�Cv��_-]���lQ_����F�F�o4`y�o���4�+�g���p�R^E�kA(Z���zt�k�t+@����FJ�5��,�[M ����@�4�_"�Z�ȑ�7�=kP�)*42�s���7ޜ�����v7�/�H{�u�/� -.Lm�r�������?p�1P�r�f�7� ��ŉ��+���mh6�d���LdSL^��U�j�HW�e,ZFve9騧P3�TF��޶o*��a,��m��^Y�2��[{Tx��V�ESg���oL��f�1���Z�D�j]!��@wזQiH��6�v�q����E���z�W
~�pͽ�32/v2��z��r�^��L�+ci� |HN�)��~�[U�T� A6�j��3�,�π�����.c ��,�2D�3�����Y�	pf|Pt�Xr�o/~�R,���0�����6�.��Ֆ�Rc?sπ3`Ŷt��J����㐜0y2cj�k~*N-���� 4����� ���FR���x�)��#�׊I�U������k�&� ڧ�ss)���R���OS�R�J�q�h8nꌾ(D��$�?���O&��^rjׯ��m{�><�0�.�T��}�a�e�щ�.|� T��d>�Ր�J�e��`��G�h,T(*k��<�f�QlY������of�e�Kل�����|�=���I���)�Y~� ��Ffʷ��v�|�O
�{-���f�9��y��{q�`��DzL�. !b�EA*K��l׍"��.W��XH=����ؕ�u��Y�I]9�2�����f�-�,+e�{�xEq)�)ū�uf����:�Hې��Ű�my[�q?����N�#*@�~+�����E28�w\Մd%�B	Z�$�3@xXθ+Yj(����Q櫱��R[r�K\�V22h	��+���+���*KC":�D�(Ч��X3%0�UX:�L�dd�Nnw�2�����&#�x��q^kDE��F���KQ�se��O!�Q���^�.�'�p=�d�~�9q����19F�	��N��"�9��n�,�<<5w�F�2����n�t�	����X��=�wF�b�Ah�����/2��d�	��<D�����=@�`eki ���5��?`��k��c���|�K���Ќ�#;��'�7�������$$�v,f�&ݕ|Ǉ����!�
�����#��M��NS����$aHɺ�O�궳zHӓ��ƩJ'D��Sj�֯�Y��G����S�Eݭ6�Xa�!��͖Um�a�nv��r���E��Aq����'c2��ڙ���t׫FxoH'�u�=&�i�ᲛbV�t)$��om:L��X��cA�˴T���ȩ�7Lu8"�Ư
LJ{�PJ��	�pnQ��Qj��2�T$rɖ�j�Op��v�rP�p�Rp<�)���?�G�䩥C��'��.P�;K>��ۆ���/�q��J�)�C���UPM��Oa�Ry!*�O.:	��f��$-^� R���9���ȸʀ�T{)qi8r�04��Ow��g�bZ�2�+T`��3��E�J���ZA@��+M4���7 ���W���κD�(��)m�i����	�y��9x?�� .x�A�����TS��A�@F��#^ڥ��r�͒\� ;g�>��u��?(�a�O� �bjG�`����} zR�0����"P����)ϛ��SC�k�H���a���tM��~�#g��.1�����(��)�B���
�h�,�
��l+���]��սy�.|�t�`�M�B�.��M�3�p��Fkz���v��pС��
Ea�T��x$�Ș��t���<F?I�X�H����#F��7w�=
��Q�#?�{'%��2ȃg�� 2G�]���z]��ЩsR��Ě��݄.t��O��O-�&Ѥ.���N��}����Ex��G��������\�^�%vؖ�B05��01��E�i�5����	�����}�8 ��fsOS��RzM�[�g��:Dڂ)�>=�H��iZSO����`S�E�Ӎ}a|�=_~���wP�h�_��؄��S�_|� 8�����|�����ڧ^�dIõ%�5�f�b�vQ_J�����"��=��'j�g�����B���ڔ��㧏���/I]0�u]�MOpc�7�5��y]%��k���2�3Yv9��7�q:ڎФ�a>�!�jlJl%�t�[�(��.�#�8�J�%�C�%3kT�h�!j���彞I���� �ܴ2�ِ�%}p�V��Y��e�4?�C�f�M�Ƀ6a�v��ۍav��{��1���f%�r������^E�]S��̸��	z�p��r'ݒ��cn"�
�?� j
���m}����䇥x:���
>�9(���ITv�d���
�r?n�24}��o��G�Rw3��iB�e����U):�7��dW��:)����m�3:xά&�W��o7((�V%MU��uv?�]Bf�Ns�^���A+�3z��R�{��z
�**@h�&�ܱ�8���G[ma����H�oɊ\҅4 )���(Ϲ��Y�=�j���nDݎ�.�z��^|]U���""�j�5����O�[N�awLL���.N�<z���!��Y�[W���!�a��dQ�V.N�DN&q��|���Ņ ��7��r��\0ef�C���J1��3���A(�J5��$�5���9���:g�G���ı��q&��\�Gs�����k�U�����1�\��(U]�֫ ��wu���	��o'l?��s�q�'�h�;�r�
�#���yϵ��X<u��I�dNӫLB�R�~�]�.(��$۾��]^Bs4�y�̤�mB�߻n���_r���a��6529K+�������mH�ePW��;�;$���%���;I�V1ߨ�GV�B4��(M^��<�D���_~D0��@���A�����w/���ҒF�6V�n�S�g���������0����M�TL�'袽9�����P����;u�R�"ՃpB.��N�S�H	��E���م������K��Im�f
`��l_�H��E�V�~�����#��ᷱ�����9�]�`��+�[�(���ϯ���ɦ�'��*� �����m��SR�9�ĈX�GBV����k��!V%|�`�[�=-��N�:�) ���S]7-�x�,��,nj���e����w%Ձ�B��b�Hg�')(s��t[�b�a�;2�|�� ZȳX����8����iu"��>�\k9»�����ӣ)z���-�R�|�5<���ŵ>&;��Z?_@�^O�qm"������v 2���|���WL$L�IC���En�pp�9�h!�.觤�Mc��8��v�u�Ô��=�C/���KW��B?�/?%UD����?h�.�?����~�TP¤�ۣV�������@��LH��a�t�׀�y6e�F��Jt��Y�B��2�a�&K+��>J"�;�<�v�LbҁXy����8��{��A�s:'d�V�<@,�}�}��6u{6o�R`���J����c��R�P��a?Ջ��Jƞ�JM��S�������U��Z&03z�o��������o�*�qj#�����jo�2���P�^������պ�f�UHf���l��❟��YE	�}�e}�^Z����e|mr�j��o�[���t��B^�ť����kC�!/ &+��p��ą�0ߩ��z�L�:�S����z]��1�Q�G�?6��*��l9���
��少�9�܉�/ހM ��Kby�Q@�6:�� -7�m��?=���	��\40"�T��Fq����_eO�h}��4<��{](2�_�{Dh#�����PgIF{^/��p}�Ë�E�x�A��k��C�[�O��4�n-�Cm��QG\�����g�ﺹ�>�*����P��Ř���"(������C�=��~�������v<.9m�QeF��)��	� ЎH�w��ˇq4l׺~�CU�>�o
��ړl5>����8�I��i��1d�6�x��n�6�+�D���2�߆ Cū\]Q���!��^̔���D����᷑�\�4�M�j{8���H����Xs�*��u�Dw���-#q)��������:zXߨ��^j�vヂբ�M��`i�\K��r��� �>���AXj�2Q�ACB�4�陦l���]��X�Wg� Zf�A��h�!�L�|&f�����.��yq��'[����UQj�I��6}v)�<�3���J|�-�{��J��!�)WE������5)�R�&nI��s�AK���9��	y���fh~��]���	��mF�b�-��}z2/�(-�B�|�ʽ3��/Z��!�d+�P�l�[�QD������ ,����W���I����.E+��J��V��+p��3m���ټ��Vȕ��d+��6��=��k־��U�{�z���,��|�o�Ky�4��Q���Z�&N��b�@'&�x_r�	�����LHe1c�#?�gW_3g��M�J�ׁIf�r��ÿ��
�Į�69G�;���Z4������>���|^tY)lS�x�C�]"����e�������o�/L�����C��!�yO·�;��I�08�Ƈ��qf��Fh���MM�M�6�J��?��v��{[�z��E�hP�U�Kq�2� n�{Ym�cka�B" �ߴѪ��}�:����?L�+Q���SƶSu�8��0�bv�T)���	r~H�S!�@�s�L�}i��0N�y�{{!,<{�<�� pW��#ڶ¸p{'f'�3�c��������U��n5�Ȧ���F @R���d>]�NkX��{��c�Z;c�#�j�s��+�]$�~���cS��=����.��b���|4ؘi(��
�.��$�e�lX�����#/�����.h� ��[=���0��.��[��,���Yev:D
T,��|$����Ǟ�m"]���I6ݡ�s�t�z-} y�#r��ѧS�؜� H��b��vZ�����۵:�����M�������8M�������M�a�Ӥ9s��W�v�q��TYγm�칈�4�o�/��I9��R˛�ϟ��2�׿T�Dąg���d��[�iC��Pz�vpޞk�ش��/ i5���&	�1���x��iħ��Ru��j&�葶r�P�^��DC�u�`��`�{����(0��䥰�ۨ\Oǭ�i���z��n���$}JȤ�8K�_��B9�p-���*���mA,�@E��w�tk[����g�r�"=_ۈ٣1xnupO2�K?s��K �sE1g���K�ܢ# B�&#�%����,�����o�����7$n[7zː
��d*�>��8�(�"���O0%mը&����iF�f�ƌ{`����I���͛������ҏaL�(��w?Qfz��r^1�I�2�*����4�Sf/�1�Ͻ��Xl��J's&}g��Vu�
>�3��
BطوI N_��X.^љ�^ɏ�%��3�%�%/����c٨���_R,����۔��V�6`^tk��a���9`�����Jt3$��h������бP�����@$ٸ�{�����q}-����������s��v�� ���:m�d���#�T�kA��t���Z�cx� ��P������xT�Zԃ��! �X�/�@��%�4e!SA1��)>Gi�{��!�X���9���Gd�RWC8��H�����*�ꢅjT����p
r�2c����l�=� �4cz#ty&���bSV��*��W�Q������U��~�+��e9X�3OuS Ο�NB��W���4�#ϽY���/���v[o]Ø�	���ܬ�8�^�5�ŭ�� ��q���< �����م ��H�֓L��uy��S�ҷ���a���.F��2HB�N
��R��rl���P��0Fz�� !5��	R�}�N���e[z���H��?�HdWl�ι"�L��/ݍ-̙6T�k��%�k0e,���:�X��Ŝ�Jҳ���Øڢ��q�2�?z�����"v�wƠ�@��Z�廹�X|���R{�n߆��	�h�5��3�O�22�w:��Uj�)PTi&�(���b���A��!�����Þ�,Z�s���F�X/��8��&�w�1t:�܏��{�}�L�4�Q�k�"�Pr*'�����H�/S��1i��J���*!N�]u|���� ;�]���V��9��v����|-Ж?�� &���!B���#P"���S�0���p�39�k42�U���w�?�eZq#�!��=�d��}�ҳ�>���W��d%���/2�s���Ɂ����w��!]�p�O��-���E�r1,Ճs�A�<`��%G�7��״�
�xbC����W��M=� >UJk�L�h��`<����w��Ux��-���[�.�ې�O�O;=���e�=eeO�6V~?����s�n�_�W`HmX��z�u\k�љff�	W�6L�.��ƞ0� ��Ȯf/Bੁ���j~�dk������\U�H���\k���6�%�1Y�P �JPi����
4<�����.l\O��C�������m�8(N�Ib�P�	>�-�t�T����Y���dF#��@�#�=�j��3 8؊�����T��%t�V*�l�qп%�3́6�H� ��D����n��VxE�B]��ޢS�����L��p�j�����蝫	����+���	jw�/uO�}�;2$��pN��"�.x~�j�/_��?O�Q�[&����}���{����c�z�����Nq6n�[��
A<LTG��Vd�!��0ny/4�Q9�p��@�ϼ<&oq�S��$��ݧ�v��j27�r���;X�[��L�+��&�W0��t�cWfQ"��O�tz�����Dq�CL���"�s�Ղ��'0^���k�7l���H'�"�ǯ�`�����r��?�[}�~���8�tnD�ޟ5k��y�B ܲ���rAv�S����+�i�r�S#E��j旒�1�-��hz���[a�[�&_���C�Bt/�~cUf��N��[Ȼ����:�X����Ʊ�����#���N�hO��9��ƛ�'��M�w�:����ŢJa.3�Ѯcd����7X}���g�wR*v���`_���Kk�y@�[z$6�;%�I�I�]R����C$:�=�m϶Z��o'��È�5�C�H��*tf98���W�O2ލ���K��*('�'�ћ�oY�P�����E=G��nɁ���2���T��-��SR���	�^l@=�d�T�y�S��/��d��{d��Xf[��Zx}�<��WN�O�ăp�>�C:Zz���9�{<*^�Mr���#U���e�8�n7~��[ѤR�Y!�����),��� ��AX.�L,
f;.{E��f��+}��m��|C1{� <�8��[9����e�
�Ʈf�3~p}�Yl5�(��#O��_�k�]f�΅��h�������>�w�)$���Se`��{�*�T%�>|O�V�T-.}�<�4P$i;ve���	�h������Yw���q�Z�e6i�逺x��`q��)�z{'GJ�VE�<���'�͆ʿ^� �58�0/)wن�.	���u���"a%y[ �{��3M�!�K.�f����M���Plg�ST���X2�`_/9�U��
lE.:Bab7Jx���F��YR�Xt��k�]�����!�<��ƚ��e��'�7�&ó�����3�=�n�W��i��Te���M�#��	:�|8�8^p��ۿP������{�����a�Z3��?Tw�F%K��7�rPc���N�p)S��
�ʨ������B#��N�����k<<�?=|�'��[8��{%�'p�z){*�"������+}ۑ���A�����&�AQѢ�F3٘]�~/����Gӽ��ϓ�Ҟ���"��>Y1���L�1�nh���S����4�����MPHI4En��Vw�H�Pu�6G`����T�@����`o�l�����W���j=fȄ1z��}�P1������X�^�Z"C�*�t����V][�M�ɇq���Y��P�ڪ/�"��r�Y�?yH�MP_�ȓ>��pV[�w_�bt���y��k�*�r��=��1F�)}:Z�#=Sݺ�ĥ;��)�k�?'���l�&����r]���,i� (xh�Tp�]���9٧.4f�z=dgQNz�&E?��9���Q����y��Ε.��g�Ͷ�lD
��y�����T}?W�*���*��O��	B��*���צWB���V�������Xy� �k�7G�7��^��W�>�<�"��)%}��*�ws����G';ӮW �֎(	6���Հ+�a�P6Y��n��^�Z2>���Z��$x���I�d�����|d
��6W�ׁ�D�Z���P���@Á�U��]�����y`HFmC�$���ch^*ݤ@��!������=2`�f�*%�F�;��E
������]'�ps��vǺG(�g��6_�Lw�z��ECL�|� ��ۼ��;'�>|\�:g͊������DٱO�+�J���f����U�l�����/j`mj�x��X̿�$�lT��gWM1���*8�m �-���+tՙ�Gʐ����O>u�ƝE~s��:�b�������/���*2�]��Z�t%P���n��YvS�n�6�X�Td�A���k�%��vb�]Μ�����sj��Y�RJC`�`����l@C�;Z�r��
`��c+����l��6�·����EI�u3!��ҟ� o�a�u���AUE�om��(��f	� ��h:̶*[���J
㝵yrn´W���i�����p��:���q������܀%`��0m��z�+���`"1��f7S���(�%4Z�)3���.1���3��7��Q�C��Tt����!�
�h�y�kk�aS���MqF�kq� :���t�I�I�WX���L����yV\���MD�D�<�ڦ�W�Y��nh5�U������W'W�@�Y6�J��;����UM���mf��{\��N=�#�Ҹ�b\h�Q�?�<$�M/K�x��A3A�g��6�H�n�Z���X���>8��e4��M4�h��9*A������w?&>��s��Zג�;Y\Z�4d;
\��{*��m��ܦ+F�ɵ=��)���	���ST:��S���{�z����b�Τ��a�и���:Ǆ
����`� 
���,rx��Q��Q	x7W�կ��,C�}��&�\�ϭ���H��.�+U~7�F*�C��de��R�ۉ���ʒ�[kI=CY�><������g�:)l���m1gK�`�S�P�{��@f�F�U|D�mBT��X�>aۇ�Uj�}'w��JZ4�>(o�Л_����`�r��
�@��N�JTݫ6��y���%�����Y
s̈c�ɓq��X� ����*d��`�}�h�&�Uf#�lh�qu-^nGЀ1-�t���-n3�F���S�2S�E��Vtf�/x;��:'�]b���	��俹;*�+:����ɻA��}���
��իجU	h��8�����YU.2�%���ʶ�m��RL�\���H�S3uOp�b�$�U��	,�!�֔�P�g�:���PJ��\]�Bats�Y]UcN-*�s�%5~�/y�s�c�w��ΠBNU��4�W��H��Z><�\K���7^�����J*{����A��:��	eP"��I�i�A�>
lTJ���Te�7��� ��S��Ӫ����竆θ��g5�=Zp��,�����o'f<h4gEH}{�WsQ�p[*z�ͤ8��o��9��B���D�F�6��N�Ԇ|1�AǸ�]��쌼xu�6E���jN��Se����V��?Yu�@]Qij�~��;�>@�-��NV���T���s��
���(q�\x�]S��8Z�8&�����w��HU�oO%d{X�e��h9�+!&���Qu��)Wu4���������3F������>u=y��wi�
����#I����&�+P�HVH<��������"�D�)f��?oY�&��$�\��c� ��q�.���k��
�n�������޻�8̭����g���@���2nx��=fkv���}�D�!�JB��.�¬@Z(FE��(ޒl��f���šE�F0�B�c#.��)��9 =?(vSD��_]�E�\ �ܮ��Ӯ&Nh������Q����}��~����mu��W������ʞ�Y�F��{�̀u;ۮK�ߔ�P��l�����1��������M<&K�3JSl�1�Q�Zȏ���3ipH�G���[�O�#�ZV/�'�I~0J�EKS�q�~L�/��(��`P��Y������6"�KБ�q����b�|�QC1U矏�h��)򄙙��������;�>Q,C�#R��r��zZ�B�V#]`�;���nJxoez9?ךx�U���]�@�����̩== ˪��v��6�-�x���߳�Jʵ�.$z����:��6Dq�ƹ�VF���BD�t6X���h�3T��9J�i�2.
$�h�odd�7a��WR����a7� �ۄ�f�a��#pd2�����`D]�*��{�����5�����gA����6)ݗ	�ɻ2��!Y�BY;z�����Q�;��/.��b��F̖����v�p����G���������&�`�K+{mFwx�a)�����["�Q�8<��;h#��Ѽ�d9��</:��2f�%�Y��Ƌ��ǯ>D�