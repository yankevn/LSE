��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�3��G?�P� ������R:$=��7�x`|һ����@����g2g���W2�I�~��0���w�W�u`r��ȱ�4^�/���1����)�V��΃�����ɡ���@��j_/Ѽ'�N�y��`�� Q?e��&���H߇�ἁGܻ��e�%�ŝ����01�TU�s~�{�d%]ǀ�+�BX�G�"e�;Ìb������{K.l��^�>Ȯ�snࡇ .�I�z�B�3��mq��Li (�
���)H�R�t@"��G{Qmj�j	0�͌�V��o��Ê��DѤS�IЂ&�)����"�B	��3��}�jcl������5�4 E�
�����8J��Ju�L�Z#���6;�f������%{���c*��9$�Qv�-x�P'�����x�Z��oX>�C�>���g���ݡv�!�e�=�S�~�+�8q���Z�[7k����z6-q�Ƞ�����{'B��5�������M'v��:B�!G!���Yq j�(�O���,{�Lٳ�5c�S[-,��e�*ł\�n`Q�C�?_���vTh�"����5z(w���S��3iЕ���Aeo�XF��uJ��|29xZU  ��f}�/
a�E�&�B����٬{���Y�l5����ʴ�k��U�x]F>��tG�<2��O8�;�?�Ņ�w�[O�V���^qُj�}��Pju)x5J���y���M�5��([ț��=�7�4.x���1��9���p�xe�( 
�����eA�9�8��MT<��d���3���Zk�7C�!�Q���g'۠]
g�$������r=T��.�7��G݀���H;_���g�ж&L�i��f#��	B��`!F�#�qQ�)'F/$�;��m�LE�i����Y�����lJ�q��O�tр1�=#s,�:��W~ ��`��:��C���4��O�p
�Rߣ�	���CK�� u>1����g�݆��p,��O�:(��W�@�C��|���;�r����P�����CQ?����Fɕk���C�+׷�@5y�]�r���?��bp�����0�A/;����8� "��_�ZSD,T�w�6H�I��K����nIZ/W4��n]��S'�{0&���W���b܂X �&��`PJi�	�q���4�4�A!y�U�ݾr
(;:�.�O�R�/�.���>T�'�����y���q@�H�b`�Y���Ï"��pwIR�:vIq6���(���UI= "���q��Bd[VV����qs�;�SZά)(D5&˳�=��Y7a����H�VE]�hZF�rdd�m%���z;�Zk[	�MQ����19|WѲ�5&�E#MM���@y�%��r��]�U�ï���5�#5wO�2я`�}��pz)�76�Sp�u$@�a�kGU��K����'zV�/�0l	��k	���Y�/�%�&���85�z��}+]Zz��s��� BE�n(�׈aD ]�m���+�~?�n���3z���Y�p�[����n��ݮ�F���0��,��@���������by��
��^SYa���\�O=�b���N1�U�`>_����3���R8H�Ssq+j�ܱ##E��z�f}�SF��6'���1�C�U(�ssY|�����z[^<K�N��B�%"M�c����ڭ���z5ͭZD����*��Bfg|�n^0�P���x��bI~��Q{ڐ�mڿW5OΓt����<6���P(s(�6X��MSgk�*��@S��LB]#>��ݹ��8E`�h���2��%z�Xy�X��MR��{D�z����K��L�
y�լ<o<Y�7\U��+i�=Zv��[i�fXG�wڭo������>�-�l�c�����B�C����L������7``���?9PrN_��y�&��k7�K��[��(z�h �~ېa8�+����=-�Z�������z����PEB�'�7̈�6Q��P޼T���Waa�gù/6�����ƞ�?\�ĩ�\ɝ;�x���x᫐�wճtFBLЀ�V1�FkP3��e�p��+�zN�����hjdlzUQ����R:A ���b�&��xt͔�@���iF����:;L��O�t����SW��#�-Y����s�Z1���0\L��Cg����4NH���	8�Y����!��(��l�^�y����U6$PX5��8�T�3��]�e=�h��%�����` �S��EX���.�5������a����@��G~���n�֞	��S	g��L��x��`�H7(V�<���X��[�U�B���]���Y�<}��62���z���PN]���K>3eK���"�K����[�!�t�v"�W$��M��m��B/?��Ҝ�y��?�� l�>��%C��k1�S%1Ӊ]�_���W�s^|�$w����'���LÛ-�xb]�7&q#�t.כ��D��js�Ah:������v�!�s�oq�dG V��ubȃ������'�ߊ���EjF$�-��}�Y��V��2����!�-^�h����
��]�-�a� T}���n�5��6���N��B�#�1�G��NE��fDdU�^�5��bj�Khf��'ؤZ��cljPO�G�oi ��K���?��z�e�������1�wƭK����B�Uŧ�w�+y̢IP.|&�[�ݰ��iEvOC�m/��PI�]�]ZŐM�-���-��?d����NǜQX�,}��KA���f8�%֏�|�|y�c*ei����m��i��w+�g:Ā蒅~�<�>� ����_N��� B���X�m� ���9م����4BEVk��-,%E�?�J|�BL��4wi��R��	��h��:Ɇ왅���²[�z�ʿ�H���Lza�,�#4T�R��&_��yixt���YHs@�O�4�=Z��p�]f\���ث�0�d�6�a�� ����|@�>�xbc�R���.3m�%�boT� ���̈́F+�0�)hT�-��s+��䬾���ƗP�"�j4;�({�HQO�{��E�����(ɡ�%�f�����E��n�h�hJ'�fc�����(�p�E^�8P�Q*��+�UA�p��É��`E��;�����'��q�� ����E,�9^�g����A�'r�!a*��2�2�'Bҵ�"dm��vs��]��5"9�0]�.��*k��Ig7⿨�hh�/Op�{��`}����+�[�/�K������IP�pN���q�t"�7��������,��\����'��	�_I���0fz�w�BHg0Tz�܏��'���ҏ[L�SL+J�c��J�|�n��!s�(��E�m%�\25�M���NE#�z=�S����d�Ka�>}�oop�\3����^n���WL!`�9�0H�~h'�1jbx�`���q���NC�D�>�r��۞����tq!�慩jF�fb�(T����r��:�Q���jY��sB����B(fX&�x���>W�{�����C�:��l���{3��@�#��gP����d�.r�{K�4�d��&V|�W���[<H��^E�TH|��ep%�<�@��w���n�)�v���j�n�~+�J~�@���l�\#���S�A�;��h5r��y��/��A��������h6?��g�8���@��������0�0"����{��2�ۚ�<������9�E����]��r�^T�E��A�3vWPr��D�}J�T�����_�+�S��bcD�&o����×���	H�Z0�B���K"!v��Q-�R��t۪p�
��Ԇ�G؟{�Ai�|V��ť��3;�uq�]k����(*��� �2�N���	��w�D��������D>� �XW4�9-6�M�� ܊`��z��_�JMB9��o9��t��Mo8�{(���KQI��M�*I�j���������'e.�(�BZ�ܼf��RΕ����m�.��b��!�M�T�g_��m;5�o�nS��q�c/��D���qRۙI��|Z���?�����t���+b���|*6aqD��}a�/D>�SO9rq9nPC��<�m5c0됌�������0<�EH�t���JH`,Ƞ�<?߄�����=\d�p��[a�����Eao�Uk���uģ�����>9sc;����h���|1����thA�̸���6�v�w�b��oV)�c7����L�LS29;c%a���m�R1EEWSLh��s�՘��d�z�2��ɤ�r���j�']���������K2�Mb���Cd��d4���X��vC���ݝH��3��=�+�]�I�=б�/lP���f^���6�΋�!�1P�	.��|no�h�a�s�L��n�����5p��X�=�{����"���䞇��=~�"�x8��b�X��>�������vq���gn�{_K�ܰ��%!�Qh�S7�=���L��a�w���&&m<������ �Pā(f�Ɇ<��HͰ~!�C�=p���͑��´��i��/��Ŧ ����?�m��Cw/������7�E�'��B'�/��2��lp2#>,�,	R�謅	��4�U~���0���#�jrM�DIV7
�Ak����%�OS�/�n.�@!q����H �c�*:�;X!%� K���!�h'<2���e]=�B�x�HzU���Ѕ��&<3��EgU	㡣ٗ�ຟ,�sP+kJe�:m� �L9��4JfV�j�����ڸ�v(=_��W��d�I�8j�s�p�O��H�8T�:��/� �P���bL�?�jU|�s$�A�
�����@���-���Ѷ%l5�*�ZT�k�y�5+!�TD�O�$���Ң)&P:�*��E����q�>'���K&��a�aO	��O���VF;�����Z�6�^�u���N.�[� ����"uު8U�ߩ�Y1_�&����� ϭ^l��5���Q�`>'�+�zc�#�d���	w��e��戯#�r�Ъ���y��`�2�z�撦t� rE1�ѵ:0�)4뤪�� r�F��+w�렧;G��=v?�ԢƆ$鐐�����@�db ag6���&��n�i�q!�i2|W� K�g�+d���d`A�y[LQ*%9t+L�6��,qo��#���l����U�+�.pBqyȟ@��28~���4�$�t�`*���s|,ݼ�4�����ޜ�g�N��:�6Ie �D|r�y�~ȸlI�H��_��ؠd:hT��˝� �$�O���PM|�\�]
:�>H��[E^�`?_N�d��KH��ka�s0>u����P�JL0���7p�mMf�^,@���Iځĉ�F�Okg�#n��oc�C������yg�q����J���W�"�?��\i��H�e�
\g /Ĵdj����bf%\'�����t��h�����cb"�5<P��G��r!�-���
�P��;p����?h��i8Հ�v׿�HC�c��4�\OFD��L�3EP�H�Z�g� ��O卻�9�OACKܗ�.N��8%��[Q�`�'+�?��x���>&9�mHZ8���g5�j�����]���ve^����j7�H���z�z�6&.`�+<��7����~��>� �1T�_�8��W��z5��ީ�p�����]��o�W���r�Z\I)*	�p�H�:��^S����ѿ�ړ�oU.R�^2T���3l`�݃sy9n����6��5bΜ;j|m\8�(�?�����h�@�Q֨�v���m��G:Ba4��18�I�H�i�� ���	Z�\�0�� =۸Q��GQ\��]w/�u�Ɉ������Opr\�%�/�@@��������7p�b��&��T4
�|��d�n��.0��g?���5�G!s�`ʴ>�ԋ�;��~�(�ID�Xp+�n����2�LE��'\�+p���b��-��f�3o����	+w~�e�w��H�u��7�^�:��RL����
@]/2�ww���HW�MyRQ�g�I������z-]�2&��S���/�}�\.8�iy;05������4pF�)oV�NHw���S�s�.Z����FƳ�ȧ�zg'����&�[5�H��/wnܨ��q����A:�JT��u��\ﳔS^d#�ؼ7�^����+�<�ߦ-��-Y�π@��P?2��4XO�f�G����̖�f�&e�g��b��!�g�|Y֯��x��XI"0�o���_x;=&�C��k�?l2��,��񦃃υ{�2��;�(�ՋL�-��2�a{�V	N�9*Kvi�%/�:�_"Cҷb�%o�7\$����Uh	(﷡���z� a�W���f�[A+LF٠��A\��Q�i6H��[�mELf�k �̒�lC�v%�HU��V�r�����!�B�Vҙ�e@�EO�Nų�D�a�A5D��zI1Ї�SH{��y�`#G3�ژ^I;i��'yC����/��N�acT�sN�Fm;����z��aoD���I&�H���lic����꒧�u+��e2P�X�j��%*��A8�����OB~5L�Pktj���Vs�0�N�M��u�W̖���r���ϥ��=���������]Ӛ�%4RY��
�QN&6���>{r���n�����fi��T_@J��JIS���O����l��h]űY���aq�;,>�D��@`�����u�g��D��"ި����J�(���J��Q�*ci�,+�2k� &"�7x���u�I�s��b1�r�\��d�y���FWJ��Y�`$�y`P�^�:���wj��^$91���C��Y��|��u'��IE�P�8�7�0�wS&�"Ƹ������s��L�N͗n�s��5
N�Y��j_�%/g����Ұj�3dHEb��=\�F���D#����#z�W�>������'�lmx�ҡ^Nx���~��]U��Փ���Tq�Ƚp����1C���,·��,ѧAcׄ�/jQ�dq�yp�� *�A�z���'��tԶ�DOr��}���%����z09�QD�:b"����%���pk�(T/�͙�좀�F&����q|�~�pg�	u�N�Ħ<i
��`��sZ��W�����M'�����A�/.�B4�����s��J�hT�%c��@X���j�@�Vy�Gr�+��.��U�����M���J��A�d�a/=~���kݗ��'������Y��1�qJõt�W�;+0�Ch\ZN�A;}�X�w�."i�>9�22��k�� ���i��Ȓ����Er�Нn.2�]�9��w̹L?�^��d�!�ϮB���0���O�(&,B���\r�-�.:�V������Jz*���ڧ#�5��տXgeÍT--�r�%)�ʃ��~�FF` ��aT�it(����%�vfE�7�h�!"�p7_s&E`ڐG�\��!��IJ�`�r�7�ӌ�9Igh޵�[gH?.N.cI�b��r���/�xQ������}��+R��� q?DzÐ@���z��&� �=-�Yc����㐖�{��<Y��b�'�P/u�w����7H�X��\��unC�5��[�� Q��j���}��x�m��6���x�G�b��X#실�)��^�y��8�����:�QP��[���������IӍү 1��΃��⍘���Ye3�޶��2D��D��\1#�Av�\�I!v%/�t�]`kt�M�7��q����g?]�ŋ���)@��1z��dr쨁dcc})aDF���룂�>�����f]�ŀd���l���yНrmo�u�*�����9�s��fA����Ŧ1�|�����<&SI�
W�I�S��}v~zX�&�,��*ѷ��W���U3��_ �Gd�!��79f�@�T5����Q�aj�61v0,�sH��o� S�Ƚ��s�� }����73���V�'��!U����Et5����Ԓ��*�\�~����sr�"g�n�7%ʣ���<!�c{�T۠U' �>u�#}��P�ܵ����-�2���l��B��yׁ�O�!0���r"���TM)3����|~鉸Е�s�I/���jk�E�]0�=�	3n�B0p;��7��q�mqA��_��꪿�ɛ����dyv���RC��Ο�[�sB��|gM�˒����	4��ƀ�½�Ռi��_��} 7�/���o^"D���������O4]����&]����چd�^k~&B�k�_0��V�k��+���Q������=��(��>a�gc������Z��3\?|G4�Hy^]�l�IpG�\dGr�Qq%?�-UT<�9{��|���s���'Lg"����E0@%�Tzr�u��iCG���S� H�Fd�����a�yt0G�C�Q����N��1�b���VS����O�����P�Pe�A�V����*����B���$��kV7ɛP�NU�I��Xk��j���°->��lif΢��%�����sz�2���٧��@x'0��¬�>��c�nj�0s��/�'�O�/��f�WCS:J��;4ϟ�	������y7�dAA��t�W��Csa߭^��pn�7E������\�C���0����
���	�G��:�
�����y�p�F�!�����J��z?�iSR`6�[��r�*���56�YX�:��	gڤ��� r�޽�)1P?Z6q�z����erBY]��!2�s�<�0��cC�zI�X:�X�����_l�+���&N�����(��px}��l�����J9��aN��������y�;if�L��E��oVã7��0m��TwM��̛�E����z��jz�����YpQ���`�7��q�ԨLs�u�����A��6��js�{X��/)Tk���Y'�'�K�Â�ߔ�_��qa	l�L�b��a�v+����a*(�H4�@?fd��� �M����y*�'- �݅�p���J�����C%>��bOs�Ы���uB��	�C�Zh]18G�}7�J�|��`(���8���}iJ�^9�S���$�qU ��˗����pCxM�=/n��-��j��f����v�}�1Vz6T��{v��K����y�C8&�f\�� �+�k��1�D.�]��K����",:yW�Ln_u�A���y;�Mrb��{�US�|��k�>���d�����-&�|;� 	Z/i�x��}�Լ�9��9N�#�^��4�3�Zʈ?ҏ��)������̱K�����dK'i㮔]�υQ���j�y=^+4�'�-s�G4Ւ&*�J2�0��oҟ1j��H��~Q'Z�����d���SnA)��"J��nYr��^��e�hv�6Q�jb��ea��fs 	�8=��E�������'S
=����8n�S(�\��=�<�8胂~y��w��z�*����Y�:��r	��`�i�f�5~>�g���D���*������nMޢ�:=�_�|
`ޑ���\���7"�� ��j�S=�9���Su���B��7�Y��0ݱ�h��b�nk�b���t��hʡ;��tr�TW�Ivo/M%�n �4�������~;�/�����r����w����XS�zQ�xJ�f�Nv^�';����`D�yK�"���H�r9��\�ٯj$�K@W���LE�Si��5.���4�s4�ʡ.]�����T�'jǕ�5 _�{���]� ��l^��K�2�U��Z��Iq�����B|�{�:�l�����2A�0M������@���,�ӕe���h6��2OAJ�X�,	���;�Yz�TdO���(��]��GC�K8w���A�Dh:��1c�J��ۨ���m�g�����~Z\o��1��c�F}!c+�L5��,q��ư�rx���"}
��q�W|�+��q�|��|pt��x�8c�r���=�t�B&��u�
��Fuf�OX�Y�v�_�bL0d	�e�5*B��RUDم5z%He�kNJ���4P�Q$�HElT���#����	��f^�(�z��E\���4V�C�dw����z��S��b�8��Pd$�M�maΡꙩ�����o�A��W�<�� ^�d2���B��=I��*M���xɛ�a�1,"�̏�:}�vf �G�~�Ph�ϧY��m����z;%�9~+^u��n�H⫚r�;�j���Xwsj	l���u0:�7�����#����֖y�D�[�3?�!��b��4a����:/��%��_U}׭Ȣ� k�$��i�|O����;�k#PM�b�5̛	UH��5���I��vdı���mzeT70ٻ#(V·?.?!���W
ʍ�L�a�5͹��d�YH[ (@�\U%��a�6���d�مM����Dh�l�#E%��K'$B]RR%l�^vv�����~t򬕿�$�<�!y;$�[���5�wf�d�o��ޝPMY�#�m�uc
�҄jv������d)K#�H�։R���*,�Һ9@�T^4���ڛ�Q�D&�MM����Myz�-��R82�^�8�y�M�U�R�����~r.t�W�]�OL��|���HQ9�7<�m:�s��������/�O��t�mh`D!�[_�>�����ZFe�Ox
W�ځ�� �TGD��ߊ�*\��A-���Z��E.�Y��Ő"��z|5��鹼6j�5��/�*�L�!�;�3��[����%E�3y�-��9(H���D�a�нؽ��Ъ̭���/'�4I�+����_���1�	�d腦=~����b��(v|�d����{���"fE�ƻ;"�t�m�3X��#�2p���y��j
��Dh��7��S���ײ�i~n�H�ϊ��Ǿʆ�K��M��g����1FS���`������"��vs�3�����dK��%� �̖x�xM�Ò:|�):���dU6�,��M�܍�	���IT����:���ƧA�n�=8�R��,m�}!k����Mέ_��he���Ѽ������qc�2S�뢥Y��_c��T��*>p6����D!��� ��!0"��'��^yPt�|���Lh���9���>n3�r�~S�P�e�~��M��<T�B��.���������i�'?A�>�а�$4ȲW��`��nUݲM�2��k/�����CC�EO��&4�K�t�Īt��(��-k�F�E���b)�u����'}`�����ZU��ǚ��˪��JcEw��Ztذ�RQ1Ӌ^]�l	�}�2~����XZN����Mj3�zr��l��}x����iS�{�F��w�}�����+躔���^=s�b����~]1�2��f�������~	YF/ao�pf�`��d�ӫ�fE�����S/?�`�w���C:����=#�.J�P��GҬ0��g��J�1�z�� �?��G�|n����ￗ�(F�88�i�
���D6*_��w����C�|G[;�獍7j��^O��X�+;��G�S�:= |j� ��CiI��憿���kE���f�1T�>|��޽����E�#8�Hr$�e���J���QȎWB"Om&9��o�����>���$��&�c�86�"q#���ǖ����hF�Ҍ���,���.:|R�sE��K�Ʌ�e�w���gRb
Mٜ��zs�kV�`n��A$��\�t�c{S��m�I�����oOҖ��Q!�J����8yQ���9a�W�>Q��'+��gks_�PQe�����a�� �����>�&I##�l��;������$�ydӑ���4-�-h�f���� ���6����HQ�l���J�7L,QY��c���B��e��o@��),��{�a`6_���iǧI	R7�$�\�_��tv�H��Q�\��4��_��9�h�$���N�x���/Ƭ���Y��k�Z3υ!�u�\h��L��X'��)�IZ��w��U��n0-�!z��A( �2ʪ�= 鵱���Sv��-8m�����o!��@/Jf�Q���Ҫ�5��2������|�A��ƶ<��C����U��uO&�D�O�T]Q0�WXFh����T��]�&!~�O,�=��O�Æ�~փ��oQr�VA\a��p��U��h�t_!��J��Ol5��h���&��ɗR�&`��ׯ��.��L"ۃ��|m�E_7�EH�hU��눴@��SVnXL/���6u�8�i��7����T	�[+@�f��%U+$.8_�-��H����C�ڱ|~��W�"�=�v��p��f��y�Ƕ��T��G0V�\tXj��� �\������f�P��H��=m�%mn�f㦶���;�9wB�FI�;&E�xL�L��]���Z��+�.(�0<"G�;�����r��a���Զ9��o��r�N�t锜�q6�y|䜣�������q�:t��=����h7��j&]/A���Vv"�~��v��[�q_zsa� ���`��C6���麟�i/���Jk/:A�"3tT6�d�0Ze���/��H=a�{y�6�B�P��n��;=���m{�0��ۻ��鐅e�a`�=f�*���
B�F\vx�(�/ڙ�~�2�<A�/��(Q�\�2��}�X�q��kj�����ƌ�⑱�轛�yZA��#>�6�X�~sWA�r9D�SN0�C�{e�iS}V.��D��sb(9�N�碸�X��\9��S�.�>%�H_!�����AHv���}��KRָ�-~�M�	�����8v�y���ǈ5y�h'���U��]��}��t;�Ԗ����z0�>�Q�9ipE:��s�=�2흊5R�NTF/�$�8A�*�/cUkJ*x�|��,�<���ӽc?[��]���q���-mU7�M&Z��p�u속�Ǆ�!y��5��*b&~��,$S��ܡ��Z`�W��x
�0��Ԕ�s�1�8�5 s���8_�p�@��0�ϊ��#$i��*����uZ�D���V9�)���(%���I��r"Cnd֏I�l����g �l}5�#-�|[>�>��"�!��DZ�	����S��G���!>����8�P��<}�m��%�LZ�Ϻ��=�
�b<h��!d��n5�\|�#l_�X��Q�C��b1ǚPm9��걖|q&��f��xu�*w|�;1���e����]_���������ґ��2���!eʗ���%����%��/�>͸���E�{O��Jh�
7@��8�`^'�F=�/�<{�	,-����W'�6���)�MT�������K�\��O1T�H������w���1�ot�T�����QBr�)<d{	87�qx�(�\��7۶�W����ڗ3���i��;��i��oB	���r�PM�SB����An�s�����Ū�RFc�	�F�	�����K�U���ޑ��b�9q���fy�1,�<�m^� �og�s0�����_@=N����&C*,��A�
��?7���"�6wP�=��ݐ�A�,O
b� �>V4�FQ}����/��"2�eO�_=�m?�Y�l��=���(�9%N�m�X_��&������B��2��t�=�vz+nB����"20�TƇ�\6ƴb��ݐ#�2O粠�-
�9*�ϱ�g)�L]��0�y���ݐ.s�Y�Q����� XQaК4��K������_o+��H���N�+N��f���x�������BT���\�Tz��z�hE�js�� �K[4��@0q~���$�8PhN�̏��:B���,�k�h����T����D��I�Z����f�����)+�'JJw)H�]��'�ϰ��*�\.�Ŷ�V!:�`��o�b��n=��#�_>+�:�� �f�&A�.��?G�O���l��pC���l�ܖr����Dn`96��dyK�ܨ�G3K���M�wE\t?yo�3��k�h%	�8�B���|5皑�Htٹ�>�r!O ]I�w��CϺ�"�F�����J��%JՉ�]�����E�AY ��t@F�p�d.�����0N�f$�Ǎ}rs3:����3�&�'���Wp�b6��!��F��ք��D�������Мy��8.���
m�����������A�~E?Ȁ��,��(��#�Lv��#`O��K�E�Y𝈒j�Y�%FT�^.#�g��l�22	X�m9>ID)E�1+�u9u�n9`����	�YQ6rAP�p,-��C��HVQ^�2��V��5��������Lj)8M�A}=��a~{�4���ǰGS8��ؾ�_.X��Jb���c�!vi~��1+�EKЧ���*}�=�=^%�F肁3=��np%�����l��2�}%����\��Z5��8s�x^F��0�?h1|N���V��_�D�@�O����h�-T��5&����cp�ے�)��93l�I�?�D�A�'m��CV�o�OtH��P�!��8��1&�Qq+nws����#q8[�ʙ?�	~���X�:���$z�k�����+�#����
k�0��ð�F�*w��4��7v�4BZ]����i#r�|�f��"�eX��~W�)լ'�?�oSn�%ԡD��g���!)jT���4�����rW4��|V�	����
o<�K3C<J�Ϋڟ�w�����T��՜]����x�;��O�&"j\��/qP��|��?O��Q��s5Vg��ϙD|��+�qi�G�@��zK��k����z2y�vو��^��v�ԑ	���׈�%z��$*�M\���M:�3��0