��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���!����hlC�9����?8�`��d9q.X�(�L��U�$hZ�Skw�'ĥ�%�0��Uo)��c�{
�#�`i[���o^i���<�)�w*)�\�/��!h`���0�N�6C��?�k{rB?��p�(��F��p��U�-�aq�F.	�Ӿ�L��_t�����y��7\.D`�}����;��9y�����n�f)�=g���������$�>H��^
�#Mї�B HKg	��P*�ϛ�)��H�JMo���򸈔�0�jS9$p`ސ����v�R�%�J2H�$�S��TY���~+c�&:�@b(����(�O|X�K��N��l/��XH2-O��|lŅ�k[�Y���^b�c"��9��Z"�P�n��.b�Q;.�GQL���k7����t�>��D�U���T$s9��`٧rn����?��8�U�n$�B�>����	Aixs�f�Xf{�P��Z�����N�W�,�&�w�aJJ��1[�%�0/�yt8�4�]55-�n��2�r��zG���խ�c7o���m�$?⪿����*}��ж�A�����7 �aZ�|�:��Im�)ãI���=�L�BS*r��1�'<�����\>ko��Nӈ��Z���[�1�*���)Њ��I�>�&����HJ�O}t!e���5�y��^cq�Ò��a$1����)�짋���~�Ng?.?I�:
�FM�rK�x"&T>q ٬��'!���#���=8��GK��K�U �L.�Q�X|��]d0C&���wo�wu�Z���4K2<��D��?�Dm���pX4�NqG����Z�wq3O�^ -�熫۴Јes�^P��Y�Y�m�Ӕ	����������''1��!,��Cj:��݅���l�*6�Y⹨͟=ɶ����aW�����>�F�gZ�("���T��(˽��'R|ztgHˊ��i1'�cW�߈�(*��Ӥka�a|c�f�r��ƛN+��]W4�b$�m��g�>�ݩ�ZT��8ҽ����OI�,_���*a"s>�!�4����Dt�h���]W0�����t�S\������pU�, ��I��ŭ_��������fK��ă5��T�5�_H_����i�M�I
P��׷�k���
[�2�f���d��
R���[�tA��<{���5�f~1����U�ܤ�bdr�̃I��r���V��Na:�?x%M�wf���<g��Ƅ�0�z�|	 j3���G%9̠�PI8���)/B��dpO��~1�G�V^���+G�'JV��:�A-,a4�,�vg\