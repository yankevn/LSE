��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S��-P�${G���X@�������P�IA\�涰�o]����u��	$L� ����Y�NC>i�l~��5���G�q�����;�3�(#�G�����0��Q�U�<�@�O�xzx���@n�5�CYX���O�h����5A�)\^�M�(-���Y�\ �ᩦ|&P�+�'�����=[��Z���3o��[��+��9���V2)f��q�n�-ߏ��(�]{�WF�G,���x���p=Ny@�mT�9>Ha��i�����^�j��]�9J�ڭ
!�W}M"���&����s (�i�*��A�-��"�p��.ݱR��I����\������F�)R�%�?5K9�� K4C�1�d���؉���z��7�1y1��0B,�ZC�B���{n����osʙ���ԭ���l
��n��K�E�"���E��t�iO�崕��\_T��e2?�72�L�r���0�ќ�Yt�S#�<'���]r�i.�e_*a�k�K�9/�ڏ�1�nGV�Y|�d`����X���YV��[MUG�����BD@7U�H�ռ��ޡ���K�������@�kZ8�m)m�Ƿ�"p�������V�6��N�e§�:�:V&���a�K2^��7���,�_N�7����1�:�8�'6�"�N��ʲ[_h�h����<p�L@���Q�$!S뀾�`�4�����N��?���v	�盬�:��2���#�u1��;Z�o*7)��O���60����١<�DKޔ�0`�x���*V	''rC�/B�TK&����{�a׮�8�͘�S��V}����+ ��F����$��ӄ`I�\����S�Dx���AgK�E���D���Ww��QG;�;S-�Kո�'�(VB�LE��,wI6[K�6���I�6	��8�IX���R@Tþ�x�Q�Z��gl��/���M�� �Q�;�]��8B�m��q��=m�q��R�	_&�	�x&��=~�"��E�_Pi��O����C��m��Auے�W�$�����vR���P��n?��n��	��^�)�t�ҋ�\	s7�8m�uǴ䚗�W�������9���8X���V�U<��G͍�q�?p�������#��=)�ʶW�.tv��*�(�6:�ˇW�5����ݓ�ǩ;�YV�rYC��*�� ��9/)�Y��bph`Mz���K��[�Ҭ@���g���9\��Y-���n#����"B&,��l��ms�2Xl)3�[�e]�\Z��Ѵ��:ɎL�X��S3�!�tnx/K���4��|HOvJ�KZMh��躗��;��A)��Zm��<��r
��-�Y�J4����7�k>U�1ڢ�)�ớLK,��|���3�}�Z�+�S�ц}P^��%�/�(�k��L�KF����;�����*�2$�͸=#b�����X�e ������Z��5��l���rOIW��sR���L���a=��ѐ�Tw�^Z����e+�_�t+��@��Q'\92��:�����Ŷ>�;�:z�X�R:yj��ī�%Q�`��h�AfDV�;��^+�s�w}��%�1Ŗ�#]ɹ9}A�*�h���`'$�ĵ59b��&�Ɯ
�h���-�Xx[��w͢4ǳD�X��|K�/\��לc�l(F���=̖t��c���*(yw�H�[�/��jF�i�����;�M���d̸:��f����U������J�jE��C�M�5��b���4:;8��U���U�lZ�iL�NBT1�6d��Ŷ��CP�.��ܖ��5?�Z����na����)� �c��s�{��G���Vf���7�]�f!�ö�œ���yiX�j����7�Vs�l �p����"��I�?���R�v.'o LmG�P^��JFA����n����2�n�a�cj���X���
9�Lt6U�ğu�wN@�V��6�MG�������3�xRN�8h��n�����ǡ"�a��gF�1������-�f���qyMM�/T2�uJ��|�grg��㧥��׬r=CVMJVl���]���X�WRʤ�����0�k��M.4��rq����>tu��߲gf)�� ��Ap�\
��*���0Ks�>�l�B����]λy]\�J���ݧn����i��8dB��/}�ޤ`��Z�9��~��G�>홧�2_/N��ɣ��A?\����M��?�I�vE��n���W��O�ߪ���ko�TZ��[�V��&�x@�����ye@��Qx�«�c&&)Y��o�>U�/�f��ax�S�x�9�"��%�$j�E�a�(�U5�=g�zkz��V{��se"�{�k���h�7T��5���eD��LL�JpN|�a�r'i&�5�Hnoʈ�YQ�����$�b�ߑ7_���'��c%u�
���,`��A�$�&�-���a�����k�!�+=ԸS�<���mf�h��,�������V�@�����1��q�W��$I.�����������Ϸ���e�M����~1���:��ii�~���]L�0X!5�<ԧ�z|�,^"��Z�)G�N�����'W�U��s���:�y8�!�q��������][,����?�gET�gV�!HȐ��T��@E�6�hɬ�lW�A>��T�˒��4����Jj����ob�dD��lg4���I�������3Q��m~f�p��լ�Q�e��Y�Mf�v*���2�X�ʺ���U��F�Csu`��bwA�7�C�NG�<iҷ#��9�x��Bד��X�=���K���]��X9�⒝c�oM�7k��P��^H�*�ײ\g��Q��*�������ڤN=�M�q�m
���[��;�@N��W.�
���wJu�������T���ؑ�9([� g�A$�]�,��\�8��ԽtIiC�I������@K%�M�P�� ���_J���{΅�,T�7���!7p��yލ��$��h[��J@� ���:2��g��r1���||r�]j��
ʸ@]�n�Q<�O���fF��?d.�8�� �G|@@qi�z�_k��F�q�>P��A�||iU��hlG7�����׈'g ��K� ���l������j���[.ӯ��q���L1��%�-;��	z���_�O0/�</�
L0T��%I��V���d���IPW��*������_����#�O
�8[H�,l�g�"��H�O��"�8��Ԍn�*�w�y.���;�1	�І�&��q���\�-J3p#K��6K$o�su��u����+�M�$�P�u�.Z����b
�SN����[ȼ��4�L�?���nģB�S4h�
�����U�L��p�q�:iY��b�F� V�isXm�޴V��Lb/|�Z��b�@�Ү]��;�L곂�7qb�N4���w_���&�j�|�v�����QO%*WʴOhj��җT�V��DN��x � � ��L2�ק#��'��#�Zz����������{�ģ!�������~-a*��`cmQD����b�I��
��U摿jX���~P tC���
�.�֪(z�u�WB����G93��g��!�o̘j�{h#�	����)�r��������ht�����ۡ�������7B/�S�{�\br�u/W��hʎ0b4�}�������]��C-N���'Y9m�ܻ�ʍ�g#Y(N.�4=]��z7� h|o�X�!�a6��x�ĝgp�"�v���|Y~��b��:�5��jL�BA�c��mZw���W�ׄ*����Z��#��E藖k��4�(fq4"w��eҰ�=D��X]d��l"�@4�WHZ�|T�"=������q���>+�	���6H?V��Wek�j�>�D�p'�=�V��
��a���U>��{���%�#��q�ꔖʜnҾ��$�~ô*;�M���"�%����oׁ�����m�"1�YQ���Z']�8���A���9�M0��뮁0�G*� ���\��}���ѧY���TC������4�����7��{�g�� �W��c=�K�����M�����cE�Ϗ���+�NS��k����D��d�!%�i��	-�&4����*@��-�;�"�g��\�,v�6(0)���4�-�5h ;�'|rtvM�(.�U�2���=���:T��A*�4�E�٬�f^�P:�=���YpH	�@��[�C�C7�`�J�_n����>�3�_j����}�.;��F<��Q/Q��>��x�`�J�o�E� � ؑ���u��٪#�_��\�3jU|a^��g]��k?P�e��?&���PYB��WE% E(E �'�H��
�����.u�a{G0=�cȀm��hG*��z�����(T��ש� �5��wkҧ���w��0S"�ܳ`�s@�me��dP�?��^���\x�O�{
;J!ö����]����M�K�h�0�w���!���{Bv[4�&�- ?AX�WA��r������hI���;�\s�m�A�x���H�/K<IvQ�B���Q�14hT�N~�)�Ԥ�8���� �`y��מo�iD+YA������\���D���1鵩�f�~�V�"��>���C���)0?����e�
��ha�wh�]�a+�cX-���*!�+�8�t�x��\��;vl�i���qD���w/�_�N����q͖E���5z�c�v��K�3�!�L$�Nb�9jX�Z#��&�C!��!�lr������o�3��h�8�ho�5ʳ�gʿ�{b ?33쮸I��^��H����LE��(��Q�GA�,�#&U�Y�M�͉{
�#s#0����q������G�;N��/�qy�����*�ŝ�[N�n������3�)��"C���I���X�q�g��!hk�c�9����e���e���ܪ�t���������HVSW���\�$.@����,�tiv���r����r��m46Ɗ/HGp�|�4�GУ;	j�7�"`8�v�aE MtJTUo�3���ȐBa��/��/K|�e���ȁ��
�,����tk:��Z*=�_=���7y�P<.L�{����CI�!����9�/(H��^e�_`ݐa��ӀgE�c�I�ڠ5[WNx��&�K��tnjގO���^q�b�U��<O����8>(����-q�xXA_����H�rǓ;�>��\ ��L����l ����3��B.�`�{^萮��$�(ȳ��m���l�Dw���#���>@v�ɼi8����2�&�����d��=&�u&�~�;�L'�D��"ˑj+E�b�uYbfp��{#+�ES^����O��/TY�0��~p��@�{
50_�1ȵ�T8H��>j{�'=�l"a��1*}s�OӃ2D�2��=�B�W�o)0I���ŗ:���o�s�T����]G�{���vp\k1������IFhv6]d��}
!c���b��]��y6���M���VY&ɧDD�E@��.�v�R�&w��za꓅)�3�A��ԏ��Z�\��[M�"_
6���%���y6j��G�!��v� �~�K��P�1k��HJ�� �cA��w&-���ws�,۲[!�9N�v��+��%���}�u�7$�@�-�æ���]rM�I��ҵi=Gf*2�Ky�^a�뮘��f�\�sc>�Q,�"a�{c&��K�X卫��z�gP��mOI�Q���Ɏ�'b��N���{o�_��3��(�I0�[�l$���.�A�Jp�2���/���I���	��x�8o
�[Z_�	���7{n�_n�b�h��b}���'�O�l����I{/���QUM4��1Y�� ����*�^(K�99;6��$������d���SBpY`%2�K�<m�RC��kVR��G����;s����ˠ���"�cN��&v�E��� $�^#H7����W⢄+>F�������d��}e�����SQX�A��� _&�Z���u�:E��U�ue'�r�싨�Iji��'9D��E����$VP������˼�����&DҚ	0����W71��⋀�޺ɵ�VC;�����J��IFͽ3�����j#I�2@Gl�� �,ˀs&_sy�8�ٯ~�H��s��ͯ��oM����~���b�?�U��8�K�H�QQ��d�[����d�ݺ`�z�����`D	<m|�J��R^3v�w�GJ��e�ބ��)1�t����!��5��m��)'��&i��T|�q[�{N�D_�qa��1d��}'M,Z����|�S�-,r
�W`c�L]f:���c���la<�����5$L�R�}�h�m�M���+Go-��םf�a�/b@zϮ��{츜
��h[q	�R��%!JO���?C�KT� 䯸xa1����\ � �b'cO䟔�a�]�y�JRk�saRq�x�<����8�����5~�Oj���[�;6�����KW%mQ�$�!<G�� Pک���4H�:ı("�>��o�eD<��z�eＣE�����)��n�Hg�#\ �p��>}�R�=[��'�
`��
̝����ެ���]l�9�����*�t�Wn�� #.ۈ��^���`Q`��T�����H�G�-n/��)�^���������k��=�a�ÉH�����k  q6��.R�x�x��@eq����ge� 6��n�^d1��პ�[�8<�a�t+/b!��8�U��!v��8�+�a�ޕz �b���.�jѐ����Tؙb�ڨCO� �Ư͇�5AG{�t$��d�\O,���N� ���Lf���Ȭ|/����9�SP��9'"e��,�yq�(��"����ZI��^�;��.��7�M,��LvM^ǌ ������jh"���]ti$+"���c	���d�k>lq���,��S;=�KV�i�L8��5y~+l����e6���D2J�V�6_���
	M�����#��:8%R�E�BHa�\x����f�yQn�O�z�D��n�w�ά�c���ڪ���e���N�ľ�s��>�uRZ�5���|w;���򩜝,Z��Ç_4J��k���Pc�*oz5�DRI��$<���dW�՝�C�:7���BoG�1��u$�FӜB�M�d�':2�ǹHz��;)�sį�|��C��l�	���w�.\�0w�ў�%���H��<���T����� >�f��{C�%E2c�>��)�-k22P���M(L�����Vй��X��'�#���2;�����؟��ۦ{�G�ju���|�6}F ,)/�O���x��,V2jH	d��7�H<kQ�����%�`���u����|8{F�7DЪ����buY僒�X/�;0��"�@C���P:���!.(�����M�."1�5��6Ѻ�~;Ϝ��B5Pk�����zӥ�6@��x�D N�4~��JLM���-{Ce	Bڹ�LZ\�5KE�y}a�YE�L�2ؠQ�s&��e��d5g�1��c����u� a̵p�r����e�ώ��:-�� �[Z���Kd���O9<F��+5P�c��W� B��e��G&<r��^P�7���&���n��H��Lz"g�m�X�S	nQ���e��N#2�oC�|�&_�@lŖ(_E��˂��o�ke�u;l�J�p�Y�[����V���R"�_�d>��T��71y�U��p��]	�m(���¯a*7�s*j��]��S�YEQ�ɂ�IP艦������*ͤ���b�;���^�X��w'6��t�մh���v�]�� @�o�jk��F�����Ja��S=şl�N��@�YG����������-Zw�ˈ_����qu��"��q��y�Z�=n����35�9I�9�Tx�a�]��i�ؖ�>F�t8�8�p��t<H�
J���G{ML��-/Q��������2�� +빭�Jv�f��-R�
�3_�K\��{_մ]:�Tm�R�V�U>�l��;�@��'�>�fC��y�{�m����������)³���C�L*���-K��A+�0|�n�J�nZ�8{�
�����q���}ԡ��q�RV=u�`��(��߸ι���#�)�i��Yj��`�SE2�!:�ƶy�N�[�G����u��@Z�.4W�g��\��	�/_��c��/�f�#��b�Ħ�䖵������b�3zڧXz��Rh:�;�%	�SL��kY��}���C�d��6G�0�T��#�Bܔ�,N8V?Ww$�̩�e��I�'��՘aa��O���eg��ńJ˳���S��zV:���\z��c��[��}v������O���S���\��j��j�I�[G�ഌ��]����V�v�����	�.��&�z�2����e�ͫ�E0.�8F���{q�ib4�!'���J��R���E���=#%آDдJ'{�*`�w�k����~�9ÏV#�Z<����UD�]*R��\��9Z�H�����9�B�U#q�v��铛j��p��_�a@`�(1��P�����QױU+%\2��'�v
��)�6�&7Q�D44�A�y�V��\��ׇ�N��m�'�;���5���-����k���I�0K���xO	� �s{״R�'� �K�q�**���C�7�S[��R�k�;j3J���sRw�H��@J� ��3w��%ň5���	3V�;%8i��~�����=1gJS��u�f9~�q��j��)����	k���D��8�<i2���t$�x_��s�$�heJ;��;ϰ#��7�:��&�r��\�2��'Hf\71����.�`@�`cŋ�,�-ޢ<�.�a�C�	���?ܡ1g�?2�a��ǟXѕ]�1��I�p�JY0u�s���#k�mH��Z������F��NBf�f�0+>ե,Z�|��y���K��@ں��8`6��d��l�=�c�D�z�Q�4����'*ю�ŋ �'�劶/'���j��sBܒ��� �K��e[-g�T*6t1�V�Fg��C)�k��ݝ���C�����YJ��YE���W�2�k9�Joȱ��1�Xn�}����5�]{��J��lo4�����6�,}���|��Ei�vX��>�`�̉a ���x"���_�6 2�cqN��+��x�q�)�%{���5g	2Ť�V�>���b�
��!�f��m�`����<��u�0�qP]G�;K�|��=q� PG�clT �%Gw��I;Xs]HH�ϭV�:D���bO�e�d�haz>�3D�Km����`]">R���n�Cc2AL�Q�-к�%�t�\��_3q��?��8y7�eq��.��ٔ/7�9��h��J���~�kv7���Y�]���Q/X�TiA*�B'�	�R��7,|�9�aO�Wp���
�o�g�R�ś�G`��R�<��] �k^\��U��s�Ѧ��
�DL<f2/�ݣ�d_�ܯ_ђ'Z1@z��C�
�����K
k��,����]h��SYI��T
�:���$l⪵BF����c�\�*4_�i5�y��t�����?,�l�n�8K6��z�Y�ٌ=3p+4��#BLt�b#8�
|ksƝFN���**N�I�t��4)�$�]������"����t�{m`g/����2�ߤr�=k!9�s%��G4=��{��W"��x+G�m�������G���B���pOH$��]A��?&��S���]V��j�0��mMIQ��Fd����`j|���rC�3V^ԉ�QU<b�ly�+�W�i�s���l���)n���sі���e�P����#�����9�!74s�O���7�O#;�OST����:G ��X��D��!#+t��d�2�:(�6�y��������Չ
\�9�G�U�\@��*�k�La;�Szt�$ߤ���Vn���ᗒ�>cn0��aa��[��7Z�8JG���;[$��O��7]>�l)���*��Ǔ�&�w7_� Fn�����U�E�"����O��۫	��]`� ��*1Q� `�� OBUp��C�e,�l��K���&�P�}��o}�/�im�$��ۛK�VO�O�J�o�L�/F.6ĭ4ย�jy�K��d�ؓOw���BJ4����)Ӊ��Bt1aw��� Jj�_{[x!_�����HG��*Zl��Kj�oW�I�O����d����:��%�~ ��]e͛};��|}����<�۰�Ҙ���^��D���q2�dYAJ��c���)[C>�-'��})�'`�;u_�3ǈR`�:J��Qoq֎������@���vp�w�FS��O��������y/L��O�L6P�{^�Wx�8q�rM����[�����.u�faF�9V��1�>?]N{���	˪]�{rae�'B8���%�*"�FWMg�1A7cĥ�i��R�o)>a.�l��9Dbǻ�MoT`�F�eRyˎ�?F�?�z���u=�E#�\���c��j�-�	a��q��N����{��MNwΪ+d�*k�W�2�3�V��Q��#Np>��m�Lw(�)�&�6%х�c�w���]�`��f,$���0���Z�[�)+-:�(��R�씿h�)��4m�y��&�'�Q쓗��^�vL� �����-�0;�QA�����wӖ	
m�����㏓��������猤̝�m�Uֺ�z�
�&D����`�-�F-T��5��e�S��r��X�D��3�JYuI Z�0y��`��=�/�F�B���FF��^��q�����[D�K�f��Z�f-��f��w@���݀*�>tl�6�痖د+���m�TB yɔ!�P�)T�G,-��\�dK�I�k(^�J>A��P:x�d���%��<��7�?���#��b�Bf�9x�&�'�����)�Ey��/� J��Y�awb��F��u.�!��$�Q�����^9�N����mGO�/ղkۧ�����ߔ�L�.�"�m9I߽���ء+�ݙ�јW�r������� 5qZ}����o�7�b7L/�J�L�D���b����tߠ<��b5f��P��Jc�i^���R�	�v�#;} �8Udg����f<�A�qc�"V�w�7���g���� ���C�I�(�V��j��alA�C'4�:��d��2�t�$y�?B�y���n��W݋�%�|J3:��$�i��c'n~��6U�G7�?�z��jss�x��2�� )T>�Z���b��>z��w�|�Eag`փu��R���e��'����n�F�C����
�p	���ײv��}��!���<C=�!rVA��ҋJ*cr}'���d���֯?ߧ)1�$a�O�����'<3[ $r<�}H�Ib���(�b��t:~��oEm����w�5��qXd�j���Q��Þ��<@��������,���.��O�:�8��(W,To��dYU�` �-��bg� �5����DB��m���x���%�t?!�T���=^����.�/�s���(;l��jXa�S����,[�2?=X��I�J��+U9�|�C�����oe�o/�:�Вyd��/���X\ۛ���,wˌ��NR&_}zt�q~���LL�j��[����4��Z=>^��x������B�;ո���no�{�=��M��(�1}
�69�������{S6�%,�������<�Z�J��a��>0����)���ݰ���c��a��啿nK�؂XrX%�]t;51]0��R�<^�2�7�8T>T$P��"�wK>[[邏1�_p����*�K�������ɒ�uX^�FxO�H�� ����࢝�mml|w��'Ct�� ���4Ic�97D���E�� �o���Aܠ���P�0?�̏c�'��ۅT8#��eT���q�6��Ȇb!���
�/$A�_���5�0ⶎfoe�� �U	��63���tƺ$i�U�-n���{������u"o��h�	a�`�WTklG甼��;��·>���gO�^�Hٷ~�80�,\��2ѱ׀���l�`'�Vb�c�-gȌz9���%�����-o�J���!&�e�����8ƙrN��GLGw��9z� � ں�3��\+��z,�u� Dˮ��~F�83^T,/G�3G�aBJ�8�jZ�������kKv�!�6�nڢ�aV��p�����w�4���
;�h�7��ڸ��C�r���^g2�f����g�#Z�F�{Sak����3�����S�*%if�\�&T�y��/q�W�9iHn7c��T�L'&V��Esw�>�U>��(D��_;ifC�Zסɝ;�z#"2�W��n����y������� D�2Q}��3���ƙ$�y=p���d���P`
��!��JK$%��
{�3�>��R5[�;~`}����əSO�iNf9�IJ�	��#���.q�B��K���S��f �1�3Po�M�͇�F6����iC���7� ������qn��q��@yi�9IQ�6�"���̰
?�`�ڷ`w,XRv�JN5n�)"%3��@�
�`��ðr��=�\
�܈G�f���P�ec����:qCx�w��}���x~��'��
1ߵ�[��
#D���-唱��"^�
�c��D��,��7A�P��^)^l�{�H~��r�-��{�lPYd &�[���3���u�zl5�3Y/S�R �D�o��Y��^D����U�P���N�ϴ�tcQ�r������c�6
�E�Q]ҫcȖf��h�B0���[Dp��m,���~}M��4�T��c�+?gAeI�D^�Y�V{y�S1�0�h��1|yB+��G�N��e�J�^5k����=!:�h����p=<��v¼j |&�i�����*��	kz���P�6��f�(*�O�"� ۹'��=w �$��(֯�)�%��+�A�ђ��+��0�8+I�[�Fk��c��6* ��(R��Z�e�~���_�IT�N�3���R:�R�g���E-��Bb��ڐ"�l"ȅ��|��R�6�KL�Q�o��q�?��Ӿӹre�."�U.*](�H����˖wW�*�M�5y�����|�-���5&i��=���'��i��Kȉ�'��uCLt�E0 ��\#�����ws�����h�c+��1�meHN���ȫ���Is�D�����Y�^�r��������p���g�G����Jw̎^,�����D��/Z&������}�AK�����T�AYH�D�,f�=6�m�ց���� 	b'N6��-Q��0G��X'��4��$t�o!�-f�B��+L�//A�������z9'3ʀ�ȅ��@DuY�k!�`۰p���<mO �G�������x���{h��S9����X��\1�/B�}_dL'	���Z���~U�W����8[Z��gD+u
_�ym��./�HU�������0�2��l�M�� �HT������`���/�9e�W��#d&i�Q��n� �)�� �rf&;4�D�'�������=$�zL�/���N.��̋!��d�-��
 ;������9ٜ�H跸`��h�H�Y2�� I����E����}������T0�XU�8�T�׷���
oyâ������d|��1!�@�SM9?�F�;��c�՛8*w�0��S��� L��6�_j���M��7a�4*͏u
�#%:����� ��uݰ0�������8�A�K��l���3��E��U��}���)�m�1���AAcg�Ŗ֋�M��0J�O4�QG�����b*,��c�_#fnd��=Z���U�6��qR�>S��s�t����㰝3�lƀW��ѓ@��1�)�/�}���%�TJx�=*k*��-L����)3sS0#�5�ड(����_��jP�/A���[�ܳ5�K�1�T��9^e��,�7)���P�U�5�S��|9�-��h����/s��� �%6�~d�ԛ�t*�:��2��ь$�^$@��7s'�J��M���V�BA�[gV�X��JJHo�?k,*����h�o;�S�
	�n�H	���	}�L��eD���`B@שy�il�2Cwf���j��-�ǯ�ւ��YSB_!^�AW_5�3iA4�L���k%�����Q^?cJ�ɨfm"'��y��#V������yџ�G�c �-�J���ŗ*���(�BM��:��C?t\u�i�J�M��
n�ʜt7�mX	�q.ر����z�M�C�;��I���v�;l��q�����7�pY��ì��b5��~��k��4����zщ6�\��d�T��!�M�~�!��������/�ў�>��f�O���)��z�4=�0
 W콼ճ�Iؗb�%��L��R)��X�(��_�	H��<��	�@<u����2'����fJ��8n�9̫��'�y�k�yO�^O��K?X��>Fd�5��2b�����I��*�Fj��iܣ�njz�]�-lx�k�Rs�(�f�b3>p�N�����B��.�cWb��m!����Jsj�A��҈+m���!h�{���� �C�8t�eC�*1d�Ą"�W�L����*v���"����La��1P���_ﲇ�ӵU�p����
͍:a�ֹ�:��m�֌�ҺjO�n�|9g	�¬&�/��I��q�S�$R�/ŭ�JK���~���
M�;�^��FaJ@,�������ݱX��`N����>�u�����z�����gn���=>�	5����)�[M�҉ke�q�:K�
��4�h�Z���Db�\\�j$�Uk6�d��Ld;����CO��G��xE�ms9����f��-_G2:��E�ڠe����e�-��q%P����)|��y��ܙ\͌�5/��)��\��G�����h��ޚ���.>s<��\�M@��i�����qV#��m��>Z��&M�lSW�TA=�.�]M���*�òY��&סz$ʯo%�6
@���\�vڢ��l����C��)X)�])uk���x�Q��{���+�>Y��	m��J��A� l&�߳��(�B6��5m���(Z�?j�M��n4�C�D��j�}�rb5�W@p���L8J� ���'�*�r���Y�e@��y4f����tKb�rZ9�<F�"��Z�XU�n�1�H�Ǌ1��r��E?������&ԕ�ǎ�e��Q+�4
���P�_Tl��2��Mىi�[��t\|��[�z�b����rW>I^#G�����1�M��xs���t܎�w��mht��{��.��&�?Oi��Mh��'�^Ot|S�_}���u���),�w\`z���js��P�H���x"�L�]f'��x�M8+gvb������s�E��>}9ݟi��ՠ��z�F��A+�W�?��7�`MwA�.���8��gw����B�<M�u�Kj�V���烵ɓ�G:�e��+G��	΂?�]vO��nb�Z0����HL�dQ��n���[m�n,�M_��^k�hm�	K�$o�>�ķ t7E��kL���R�-]D&��;��}1���~D���YX�wl6c�C��-U���Ŭ�"�&����+�
�	�}�1��kq�����ږ4�9����9	4��uB
��:�Wۋ7)H9$Q�s��U��e��$4F}R/��~b��	T�
}5v=4�|z����n�[8��ƧfJ��.��q
�&6��:9g�d�Z��ۜCIV6�ђ�k׮�h�a覼�vV��^U���끦����A�6٪�-3=�r>a��n���.�n%F����[�T�OځT��)�hoM��t�Q�i���p|w����M��eH-<����E�P�� �N
�� ޅ ���k��mT�#�&;C؝Ue�e@���ǖ�	�B�7bʤ�l�썈��3���4_�3E���r䥫���o�h�זl Ķ�ʷ��~b�ES&�����F��hR����VZU&0�����5�	�W�hly��8c��"�=:�2}�f�
SY����91|ܻQ�EܰUd;�G�"h4��4�O/w"�i�\���z��^Љ�+��^��6��u3��d҄\Lg1�Y��>pݻ&[���dG�{o�.��t�����C1cOQ!�I["��ef%^�l3����/0g�#�(�1+��@b���ʣ9�ɬ�EE�����\*	�c��= �����S��~�u*T&-%��0�S;�.�"l��Vg�:����R7��}�2�����CP7V�5�q�R����9��tt@����3胮"��2��2e�<љ���=�������V H}�?Y�����|k`�>���$�e�m�E�Nz���>���<-�O�Pey]?E����֘��C9�+�kJEQ*��x� Ծ�Xꇯ��g�7So��Ӄ��;Ԗ��|�Rw�
����f�ƶ=�g��`3�(a����Rz��A�ZA(\N��'ҝK�����=�t�33^�c��>'��"�5͒��8ɐ#�����I���
����_o;����*��U�/T"2x����J�	
-�e�dp��LC����A���� �U3iG/ժ�� =�ˉ��CHXi�LP���,[�
��	����4VQ48n���S�c�����;؏�+�z�]y���E�CaP�_���:�cǄ;�����YQv��7�<��(r���n!��{6�`l�,���멦��H]����̽h���� H@αΜ3Y�����wTݽxғr�9N��d&  co��;J?��K��,�9t�O-�B4ce/�׼���<���(cGWVg��A�f*�	�|������`����e������r)��� �([��ۄ�Rv'"��Uk�LA��.�[։0d!�RU�N�Q������N��a��^E�>9(˺�4�ƞ�<��b]�����D����6%�M�Y[���EO���ʐ�KA�TW+A ,�z��T��ݫ�"�(���v9���������C��9/E�����!��h�uRנ�O�UE��z��$�uՁ�!�>&j�_�lf��a_.�ҥʾ�-���;�B��˄%XN�Y["PBCS��_yBS��+��p����J���?)[�)��$�id��K^1Y&�J���}X�\���0���P�K���O���b	2���
��]-d�P	M8�l��\b"L�M�ٙl��ܖ��b5dU -e�
l5.p*����������&,��1c� ,���;jG�7�M+��o�/��
DDmjcx�^�Q�������7�w(]�?2$\hpBE�NQ�L@k5��lûC���$��59�����!?�-ҀҢ�\�Ũ��}�dLj�%^�����М.G����|��*���Y�9�t �ݙ�A⏬y�*�vM��ڂ���1+ -�(�`I��9%<a�Z�]�h���*X\E:�5̽A�Lb��2
��J�ꁓ��X�*�'�c����:O���i��z@���,�A؞.%���_k}U/^��s��׶��W���S�$��Y���*Η�s^�W\=�����^�ky�y^)�����ʾ�VZ M�`��e���1.� �ńq��Nr�P�{HY���(���8@�.F����h!�x�,�ɖ�V���T�a/F�DU]O{��6�G~�дx�'H��.���vs�z���,˪k�Ԃ}�M�jyWͲF'"��ޓ@�$~뙽+�S�_�����F}Ļ�D�iMdȔ3����Z���((���)P�گ)��-�&�����s�-���^ìOJ�i(a&�u/�c�fgJ��\$�!	n�����c*M��[w�Yi�U��f�/f�Zk& v%�6d�ʭ�\�P�����M�2 �_O�]i�1�V*ᢷ0n�k[�I�?u�rg�!�u%%�>^Y,̭�{G� ш���Ӵs	��XR;(* �H�2gn���Xg,�����Q4��m1k9�[ԘN*E��ĒB�%f?2���KCm��TC�Ůg�h���1�F;ݱ��XO��\%�v����pB���-C�D{2��v(�� ���a��J1��/�E�q��N����+�`R	�P���ܩw�4܋|�p0�ж���‟�R�
fqg 틵Ѡ��ʭ�i]w����8�/�n.���ԇ��o3�2�4���}��!  ���O��~H�Y�߉����>��#ϯ�03�exb�ɲ�ʋ��Y��Q/C<zMIw ��]�f�c'$��"�b�Z׬�/Y�d�3
3B�dd��[��O�݇��Kތ�%X�V/LGNE7�q���{QYB:F?��kW��ܜ���ƈ'a��r���.��-�H9���)/�gJS��1=o�<(���]$as��`Ep�.
M'T���(���I�v���mx+����9�hJՖ_>�K�I=3a=c���6f<d������я��H:��t���>7�Ze�+ztփe��<Fcn%z"<n��
��$���9݁��qM��Ő��{���<���*�얪��������@����"�N�I�@n���x�=���g�4B��W��ӂ�t���s�w�l�#�?�e2�����g�ON e$k�&n=�x��5@Xn��v�O�:����T��o'���������`���@� s�t�
\FP�R�,7M�Hj"'2W�{��n
��Z .Yl�}��f[�S��9¶f�"�_��T���E
c�V1����{�*{�42=ׄ6!t!Ȋ��|���(��B�:#��h,�9�й���_g�.r9��p�Ϗ�k����������O�$�;T�\$UU��yЎ+���m��ʷ��ǯr,�.��e��R��"++H�
���� ��@�]����~��JqsǨ�*H����#1����~?��`p�_�$���_eC��}��2�uI}M#'<�mP(73�,(->��������4Y\0.{X�\��z��``e��n����)"�S��nˋ�.�M,����f�?,j�[N]Yr=Y���
X޺���}􎳕���A��4���B���s����T��#E�W3GC����*-g�E'kL���ۇ������B�R�k>����`?�R��e3��Ec�9u9W���U�}Se�<Y�IEI�`�'5ZP[���Q|��x�۳��xGr�Ƀ]���ԏ��m�u̒И�'�rT�_U>�'�u!	i�5Ӣ��rt�,��|��e�P�3�ג	�_�o�TǸ&�A��v2ٴ��i��/��n-�<OX"B^n�'�74���;&"��LĮ�O���ٳnۅ�L�ߋ�C}�D���8��J:z��S'h�A=�m��q�|��cn��2�@)$�ҋ������(��n˶�ksd�k�2����fF�c��|�/-cK����@��[g=&\W	�!��*.Z�(	G3���Z)��)ٗ��e�7$�=ع��RiF.�b78�#�ߗ!��Mv˫l3��I\90C�N�3�b  �Z�/4h��v=���F�:��ݲ'��.��B>�I�˺:m����4�=�� |��+��G�
=>M���p���[�r�iN�K�M�\�g��'R}�_#SR��L�7��G�M�6�kh1c�"����CK�i�dE�-cq����q�L+�����l�#꽄wׄ�F�q=^�LU����'Rݳ5�DǼ���B��»IZM�#��o"T��6�g.a ��6ӝ��d���O�k�Aೋֶ�h��=/e�cQ���)B�J��S�ث7���Y����˚5�.�ŉ�7\�M�<x��'s�'�U2�I����SgE����X�233��s��(g`IT��|��<4�[O�"�
b�I���^Rɸ���U���+��F}�e���=�Ey, ,I�2U[6��!����jL����-�]���ܼt.L�}@R�V��2G���=� �-?>'�EV�����U�r(@Hq���nc��!	q���y�z�o��1g��ZE�F��8������8�Q��	9�eK(��w5��~�"���>��Y���Jb18�1K���7)3:�uT�H�>����C�0t"Ro�F�i2����z�y�?Am�x�z�P �_.x�H�Ĝ@��M��4P$�Jo�[�@� -EN��?����O�E2�B����£@���w���˻�抮����^N�6���`�r@8ag����-Uc-´E66�C���
	�!(��tV�*�C��Bi���G��/2�9}3�1����J�(��x���7S2�|�l���9�G#ښ����P_�־g�x+})g��\�S� ���g��� ��|�[�O�wR�>5|��L>J.�P_��w��J�N\h4}*�5�dz��i���&m@�6��PN�(i�P�+���D�ζ�:V�ȥ;�s�ۜp��h�K'f�0�����U"����&�
���"Ҡ���S����F��,'�IY��/�|�+���E0�P��;�5����$e3 ~:�1:J[^n?>��z��V^�Q�t߲8��!cH�F�:,���v�HB&l�_�Ɉ�Q `f�\�_CW�t�R	*�,X}AKӓ��y��z"KU��y�ԳC�R�ِ��UY4������G�f�TM�3�6�mˈ|ˬxe�PV�| h���M�
����/�N��6g����q���+�� 	�N'|�;<@�A�3k�@wf*�5�k�iTe���y�H'�%�׋�1�W�ԊU7��&8����͊d
���ʤ1�!��,�8E���� ��Bv9s�v��֡ #V������.Lx]��=n���,��;�
��8� ��*�C�T��Ƃ>���R������u*�uWѪ���E�J�x,Z����gf]�f��:�[�t��Xكfp��CU�'�*��.}�F��#��s�<#Ҍ.<�>�Kv��g�Upfw�q��~jT�$=��]��fb�n�@�%v�[:��xF���j���'\�&i�6�s�sB�����7�
0ͬ\�(�0F�6�ryԣ�[��<���'.Q��$!l�z��Z�����1�d2���6=D,{���t� .6���"z�<�}.EW�V�a�JnS�åK�xY8ro#� =R�/+�Mq�;�П׈����7�`��28�?�"��-�?��$+i ��%�<R�A�����B�3qm�Z�3V�C�xg�,̘V[�{�y��a�BrI
=$���ƙP/эoo"�*�1�K�u7Ϭ��c�zE�$w�;5O6	�hFPx@����b������r�ٲzR�Ҏ����nd*�*������4���D]��P�|����Q�dAS������9�D��SZ�|�/r�t���_`��;1��͠9 Xƨ��w�����Fj?D9���}>sț8����=W�@��Ƴ�O��ϥ�4t���un����G��t��zn�	G�ۻ�z�RT��?�Ňl�C����!4��qX����Wƅ�T0`~�,������­��&�lcX.i����'!�L=���g�!�p.���W�>�fs�#n�s-��hKr]	�Ф��~aNR��M6�;n��\�O(ڀ���ch���D��0$k�3���C��QS(Ţ`Q�r�����B;��b���P�#c"�n���9 Ct`����M���L���F�h���ƨB����A�8������M�to�ﻻ#E&�ʹ����c�4�~� E�=�ի�p�[�eRV)G�u�@��Q�"��fS�u"�L�
4ٍ_�C��~���wt��C�P�����������[9+
��]�H�tOe��"������7B�ȹq���CF��qf�*��p�B M:Z�ĦH�x�9������v9�ʛ���/G��*T��ݹ����v�@�?��.륙��Z��`�{Q�B'Ѡ�1���8�rٴ?ϟ��2�+�zӖ�n�`+P���/B�辤��Ｐ��H� 2:���0��w�����6����s(g��.�Nlv;�����3����h�����p�A����׻c����t�R(�pϮl[���R��1k�j{z�����%��l���	��8vn�$<Н�_��P@�~xY������rM��{)t�え1��!�+��xz� ��Eg٦[�
ǁ"��Y$�9�uf�t�Y��@P!�Z=�f�.�B�-��lNu��K5%��'.��YA<2�"Vw�
���֓����+��i�?ZV]��S���ס*Qj[�|���AޗqO���T,��S�$��b���\��Q�X��D�2�������^w�'f�u��Ҋ1s��7|�ʉ��(��\R��Q`|( ]�(�"y��[�]����dK���V/�VuU����7��M�a��2��jLp"޸}E�����lc�Y]ۿj���/dʴB�y#��*M���
X��l�h
�,g��D����{�`��*4�-~ub��e6l#*�qL~��*��̤ԣT���Ѵ]�CI�AF�'�T|)F�'�lF�P߲� �b�����!b�v4>��㗉�m�A|#���MJ��g�V�����u����̞㬧�-����skؒ-k�+�.���A'>8K�h�ی/'+"��P��=��0 �j��1�?�*�d�>��/4M��2�4�RW�OxFRy[�e�%��0����='ʳ����^R�0�-κZӆ�g������#�[��Z����,�	�h �E����H'�y��V�W'c��� ���U���S��*x�Yq��E�ڲWfMh�y����'�xwF� I}��tԒrpU�rr�Z՗T�{ݞ��4VQ>�!�c��D/�[Y��+��i��Ɇ��ƙğ-��,�<�iÑ���d`]��s���{���J7��a��j+��)�N��o�u�� #�G���z������!�X�ɳ����ǒ�%1j���V|�βí@��3B<��
�tl�Fsqay�	��:�޶B& ���3�a��u��՟���ˍ`�M�&,�N)�@���f֯ID�|%℟!bF��	��K�@��%�c� �wpߵ��$�h�Eu�=k���V<�������2B+6�*�k.�����:��'�+f�����ؓD�d�f�3^��|��0ɒN�e�z��P�m�TL,&Г��BD�����㫝�h>���1���.��{�ɉ�/�<m+�AS-/^u���a-���`�0��s���~ܑH��I{��L�.�q�����w��,��Vu \��*	����\r��>!�+6�1͇Sh�ED:��"�-c�L�j?���q�����{L�\��E�>DE#hj#��"F����6>��#���R*�
_0���y�w���PF�CO'��x�#?C���A*
^��
{��o��%��n5Y��+֛��hz�X���>�r�2Z�d
�T��MW�-��\���q������ Y���'kN���^ȈD������)W��?����L��'3w]�V�%���6u�(=���Ku�>mT��V6�cRU%��R�?Uv��d�"&2Py���ƌA�ņG ���3��֋u|ǆMi)�E�wRj���%�A�8��ܧ�E>(��S��I��Lk����jtڎp�$�v'������7�� Xz,='�e��ȏ}
�_\k(��P�m��	#�8�9f^[*\����=��L}�vs���L�]��Nj���ӲT�[�fT�/�M��V�Lˬf���:h�+e+~A���|�n43Fm���v�pb����S�F����|?�%����Z�X�����aU�f���ml�=�������t��{��H��H����&Ɍ��������d��\��ѫ��B]�<��P^{��f��]T�j� @�ʦ"~�sWp>����e�S�%"��x�A���Z]����z+&2�ϸ�EV�~�u�x#�a�	����&*�#m6eJOg�H)/MP��t��e7�b�
&>3QK�q��������N�eC�«pW�6���̻��FzF�3�N5��5�2�@�"�[��ˈ/��_�!���9�+�x�C֫���j�]Y�ۂV�t\4�$sUP�Di�p&���Xe!̢̺�'�֠y�`��Aޓ�Y��bG��g�[k�3a�_*Q��k߉��tݝ��٥e�1$���= ���뭘w T��7sN��Zr��,Iv�bל��Y����OD���*�	��.R�q��s�ôއ�r����Ņ��f����Nߢ�~y�$��w)�'Ns���Q�X2UK�۟v�����K�+N�+�ϩ�ԝ�T�p�Z>�4��L-5�F<2���ND8]>蘦Ӛ4�t���/E�'��)��pO� g�:J�D�*�'w���6j{?��?g�Ї��V��j3m6������Oc#�Q�c䁒�"��oh9�O��&<���(��O�����B� ���P鱕o�����o�Y �F gn�䐶\� �
��X"��S���ȩ��N�����j���������WAr:/��-a��/�ˀb�4�L��4?���|T��-�S�rW3;2/2Yծn<���_�䯀I��\r���f���"�+��r�d]�Z�iI{a�{,���L�
���o߆v�޹��5�
�w�����n�yK�,1"b�k�C��~?+�9�k�
��5�#����0��`(Ed)/�0�$�z�q(I߃%��_�3U�r�wM+&e�b���m�F퀹�Z'Prjaj�GJ����^��k �o��qL�ۈ$)� ��{�/Օ�E>ˆ!x���H̎��p��8/���%� n`|������6~|LQɳ0����c?G� ���8�����>C��4*�S*�L�s��.尙xrQ.;��|w�(�V�X9�>E�c�/�ťl�2	.*��)4P�����V2E1����
T�:ONηr.��5�/R�O�n���v@���֬����*�A�QJ�d�!C�8\�[�O��Y��Cjp��^��D�1kzq!\�HE-���D�&H=����"�2���m�����[��,����s-k@���4�]d�H[���������~D��عj6,�Q�$r�Kǜ�!�V�40��>�o��(�2a?M8�	�<�"��z�i	���UѻŘ��I ��d'�"�F>����`��h¥6�ѳ|���
��:XX�mUj��_2.��b�Y%����Lc�zbcH,�i�u{T����"Ms޿�QC�Jy>�_{i���� �B�'H~� _�7u��uc ��_��h²_nܼe 96V�BTS�47f%��I���۪���&ݛ/&s������g�w]�q:�n�\ �=��L���{ժOw�tW�t��h �� EdGЭ��@��$�|���R��T�}�?ƭ�3��M�v��b׀>��j�>u�#�D:�R�bS������Kx��ڸ�C$(u�Zwq�,ƞ��������R�g��~��`��q��3����m��v@���sa��	Yt��IĪ�@O����ngZk��
���OK,�ԸW�z簋P?[�_��
��L=-2vk|��U"hpo4jܾI�y�.�]��1�[� �����)q��X5<	����Q)JY��,� �CW��Zء'm���,0	�-Y�0����C~D*�q|�+y���_�o}L���!��.|�k�h~(s��P`$C{���ȻH����8�bf^����(�?�] r�ǩe�&Q�z������V�;E����7^*Y�(-�If�ˡ]��7F�"�Vs��a����1�	�����j-��C,պ��V��R�SD͇�Rt��x�nV��H5�ūm0�[��<Z����c{�ҋ���M@�������$W(��B�#����6MPr>�~W������|��Δ�3���tN��<,蛦���wx�m୭N��hΝ|r��6]_"'T�=���:b�3o ��9�dc[8�+Q���YJE>����;SN�jr�����Tf��cL+��@�R �����(�0��v�r8u ����=(\k7�6���
�-�7��Oՠ(l����̐}m�5��Ї�R����c���U4Wi[n \*�P�~'+�7�Nһ��*�jAK"r�Y���H��hW:6�۶����`n%*�5]҅~xi�+<٦��ϰ3pL�����gFqm��]v"qUS��[#�b�)!�c�����m��m^cv���ɇD�N�	�,�$I��u�+�kHsE�vJ�](�p���K ��O5ϙ�����Р�U�d<4�#fQC\���C�J$�M@8<i���	��m%�ĳ��
¾N�sS�(���P�֏`h-,�%5䶋ݻ��9bX��K����O5����;��Sؙ3���9���1��zK�P+�;��P��<\g��P#f�y�և��M\��Z�FIW�{l����Y���[����ʿ�C���BJl2��d�ttxD!��������2�vԂ͞x�'e�"����U_�ؿ�d�F���-�g�f[s�Bq����ŗ8�y�B���(O&�j�me��=�"?����U���vQ��n�퉽��陨��DЅbw�����G\��3�ǘG��%�3mo�2���)˸��5�NG����o!�Tp*
�����<���*Yе�&�)LǸ��v�ne�q�J�[��Dp@F���#9�w��C��3����dPL����63W�S(���"x<���+w���%�������l��&?�Ď�s;�f����� �O�h
�d�87FG���~�ޓ�%wG8Uﺗ��o:8mڊ��Q���O�o�+bZ_�����sw��9�ִ챯n�`F��=�P�B<�����ti�}��k��f@Lx��*�I���ҋ���BH`�Vk]|�RQx��#���&�v;x�E�s��3iv�����*0����0�)�+S���Ҁ)2�Z�O�0GIT�@�s�t�C%��.���#[ ��^TmfBΊp���J�8��O�8Qc�e\&�K#���sN��;�E���j���+���$�z�h��b���t@�חk�_��^�:c�#�C��V���4�y;���O=W�N㨱�m#絋 3�H0*��	�Q'�N�ev�a$Ćw�y�?���>��K��\ހ�d�(����KWo:��#]�ttw5�I�F���dZ��[Z!Sܹ�~בBn�Q#z`���
Ll��oI��Y��7ELoK��su� ���֎`�xp���A�_���p��d�6s�������d�?/7���Ŀ8�j��4 "������蕈�(��B� ��a��-��ܔ�_@s���e� �5��\-���G���+͂TM�7gX6\�������7�ѻ6�,w5�H3�U�2�fC��Wy�P��Yq�t�M�$���0�;�� 9��osْ��v�l#�Π�$�͖�5	����uS+zMnB^5��I���͙�h�t���Q�>��p�NJ�����~Ŋ�V�˅ˎ*Z*������Gi�d��&���a�m~_��J�t֙��	��i�  ��5�!�7ϷV j��Yo{Ԩq��4k.��L�w.2�ːjcU)f�Z�꼮�Y�^qt6ڙ4�Ev�Aq�T9�yxu�R�Wf�*.0�X�ԢJ�~{_ā�����J�NM��i� �M@�h_mU��z��EfHt�s�`B�:r��p��<��o}�n���"���Q:�Nb�nq����00�u�������pEԈdw�E�l�,'X����B�7�v�ގw�v��+X���vvi�U����Ηd�wB�`k�m��<M3�|{��q��O߫�w2�
��f��D�_��eOz�����Z������P..>�T�G�#k�G�8��)Oޑƫ�R$i�XE���~�� :"���Љ�'��-��E7F#	$���gC��N���罭��Vo�����ы��&߹D�f�N7%,^ޛS��`[�X�v̑�y�`6��\�
�#�#�Y@���Z�~��'V%b�x�_]���Yb��w�L��Νl���aS�L��e��7�!�����2�A���EJ;��cu��B���'���W�t��x;��j44G
j0�p!������� �{@�w��I�_�mga[R}�Ӌ`L
�Pl7k���(�ꃑrl�b��SNry&'{O�OA+�o6q_�׈���h�n,���d�-&�����I��O��:�'ٲ��t���1{ <�����brO�)��r�!.lRܳZ.�T�QD:�߭�Bm���yhG�j���>ש�?��1�-�m����Rxx"K�a|\ɟ|]����_����C�\��,YS�|F ���emp�5*d[3�+4��'��hD��d��\���|mn�!��렷�?�E3�8�i�/m�jhə�kE�!�}\j|�����y����P���kp�*r.c�L�G���������h���ʟ���=�Onc�=��;ֳWc� �|��Z{���k�<Jہy���0ưCN���/Q�p�:Q�P��Gj _B.dO]��Yy ��%o�>sߥC�yJݾ�h`������hy�TR�&z
ƴ����&� F��3��h�xK �����%ҟg��<���I��2�#� � sm�-~�T����z�Sf���	�&B����|�R���w��$�b��W2�1��5�ZoZ�7)(��W0}Y�B��0�HmS~�<$��c��!�.CV}l+��У�U�-W%��uӨ% \��_�/�-(�ȉŨ�d4e��
��-���k�v���I�������\Qv����{E�O�p���ԫ�J�$��?btʒ�� �E�d�Q�����5t���Q�	�N��*��>�C�zC�2z�.�z��5b��)TY�Vل!�s~�	hY�� i>E��TR@��^�W5��O0s�[U�W_+K�Ӿ�Ȉ����S�D���dA�߷�'����ZL�R������qG)r���W�R5+n0�V�3�1U#%�]0�C1���%�9�7���K~{��h,fA��Cx0J&6�fE���Ӆ���3�0Fu#&U�\) �C	}0ʧI�HG�eW����+�����>�Z��v�һ�m���1��ljw�ߔR��* >�r[�#��_�Z8��~�sW�Ex�^Q�T��8��"�펱�o�n��&�X�3u�Z+_.�*},b�dA�epH#�]	3$	�c���zꁤۡU"�o��Y�7I���{J��{dŲ�ve�Q݇�b�78���&�{��:�d33FEܿ�7��<��)
W�>�B��e&� J(I';��Tv�p�E2�#
���7[��U�MG�T���ׁ�􀞨\������Ks�m��� � �z�Α	v��b�>�5�6�\�RO\��˂|!�Πdg&�\)��0L���?*̚����{��|�x�oO�����ݽD��B�^��-�ma3Naגh�'����hm��K���W/%��[���ۖ��;��¶��u��m;$x�5/8�.��*6�2�dpKy����b��zjw��\��G;��)�$U�� ptc�i�$�;��	)�c#=8��IS��:��;����:0�ּ��8Oy~~�K6&��hT�?��I�YQW
��������0�m�}T)�bT�5`��!��N'��:���~��y�BB��`]G$B����_�ޛL�˗��r����j��h} )E�R?�c|>ۼ8��9�}'�Ϗ��m�a�"^ð+�З�<�W�R���MH�0�ٶT�*�]FH�yy�WS�s{#���0C�y�X�*����'SP�=������.Cr�� �nL)�h6�@{�����l���i��y���NFz�B^��9�{�� 05*�� �3T�����
�C+V/�����6�E4�
��v^@]��R����	Y:���{����熅��KcܻlE1$8@,=�~��e{��a��o�� ��]��1ڇ��Ѝ(v箎>#�}T)@]�=?��J�7�j6��y-+��#�x{({5���de ��mj���j�8�@�F�2��	\�YԶп7�{�'�cd��\�QAsQU�0�����C��3��-�W��0��k����q,���m��2BF6�#Ѕ�����J���-/ȢF
:&O���(_#E��R�y��Ci��Ŝ]x+L� KPF75[x��l�&��d����R��nı�[�P��q���ݕ`�	�/$M�^ӡ��K9�Qs/b0��BD(�J��<1�;H�{�K5r�Ejƾ>�i�����<M)��;�d�At���`�;=f��y��K�����o+lf�{��ܒ(&R���y"�g�	
0���'A崯b�V���Y�%��L_I��v�٫I�ﰅ}!���F�ew���a61��awnR6�3�s��d�*�w#9�^��kt����:�1:,����:�u�d:;e�`i��l���n#8y7t��0.��,ۚ����L >@:Q��3Km��2}+K#��rV���!!s�wM��s�2�Tr�{����H���+<oyC[o���7kF���J4��긐�Y:��\	�V���zv2�C�}�'��&�o�;_��@��А����8.�d뚱�6��v�2�kQ����䞏N�ےB��'�i��O�Y^خCG'���ˉ<g�h�(��Uc�"�li�Ƞ? ~O��*���'��������@����P�Dڋ�Z� b��5�� pEmo��˩�U�K�F'�)/��~�]O6��cRNVY�������*�M2e(�ߩ�!�Ʈ�6�*�騚������E�DТ�]���;v��!��-�/��Uz��v�6���2k߰�쒟�ݡ����|���E�&�}��52�;�E�*h�1JA*�H���ŬP�%��|������w��~����t/�����c�g�C�DB�GҮ�@�n)���c��V�z<�=�g���f<�z���S���_{{n[Z�9j�6 �8�OV4���e���_�p6�� ���I�z�^%~����5�)k-6��g=��Ĺ��	a�$���;.���0����K�U"�Q����]W�m�]�Úȑ�,ք�B��ǯlc-���.����G9�l�R�\Kqi�Fԃj�斕b�U��-��Y�i5O^G�d3Tj
���$��l6@�Z�a��(�'����]>��L��M{��RՎ��,;Oԅ����z?	)K�8")C��A�a� p�4x���m=QXZ|��FP��@��V�Vؠ��I!Y�$ut�W���r��C��z��.�5d �v-?���F��%��|avm;%+�S�<N�<ް�<�������ش(|O��YY�p]���%�fwS�������a�!9�|��ٷ�]zʨso��\*<_�sXR3��eR:R<Y�Z�"���-�bt�+���>����0��Y�?�	Vfs�a����l��Z������K�3H*������($�|�ϱ���@�|(�&IW"Q��'����n�A:��r�~0F�4���f�lS1T��%G= �V���-���oF�x�es�<��;]�-�?�BYM��Mv
>3n sy�uat¾}��^���e2I�aA�'��&��n��٣ke�R����˞�HJl��Ā�Yx���zb)�����\�o�P )dsظ��e*�= ~� [ַ��?�l�D9�A|�´T��snoqt�ѵ;Wt2���
���6��Ț�<������7>����r{�H�gP��.�/sa�~��e[����2��c��ӌ?�׮���B=�&���$�8W�37�h��"Tz(OZ����k����8���|�P/��Ǩ����� ]�yq����x��9����$�	�|~��p��r(����'��vՄ]S�c��E�}/刪0^ᄮiZ+�|�5-����(i|)����"��?�q3i���5%�����',AXCE;���Or��f��˳�7$�T�M}s2��)�`��\�;Y��Jͩ�
d?����8 �1���0�1�j��S�P�����b#������Dd�Ga��QIo�i����Lm�9B���(�����:�9�9FĖ�A�e��},]�[����x�̅�1q�$�P��rk�՜��21-�TV6�D�ܬrH֮�]׳x�^�9X2@sɞ�=��enu��E�ǨLV��[�^Z`�'I8 ׸��<y���cq12�?5�T����e=���d��
�-%�� �HqN��_
΍�y<
�� JǙG�S?ÂS�>��9@�|���ˋ�2	#�4'�xTΚ�;�HK�ʗ��8LT��p�>d����K����w�` �ƥ2�߫V ���J�ފ��q*`,�oU�h����x+?𙍕V�DU�!
s��Ə;N���m���*+B�{�	F}���d;'$�p&�Y��e$�i	��F���a�W��q#My��c&�?�Yn�E�����Z���Fp �t�����8(vLx?��0ǟ'��$�r�,��"K�Ҧ��`�7͡�Q�����kE]C+qQW,��u���9wMs<� �e���Cu��Y	}9��F��T�@�=@�MաA�M-�W_N�+Ԙ	�L!Uk`G�f�e��¼�Y���V�'�И=��T�B�<�3m� B����;���/+�cn�'4鈩[I��=&|����%�����o��h��(�1�OJ��ۦc=�3T��2����� 7UG�1���=yr��j��|�ܭ
��
�C�̟d��LA���T�mCܫ�|�L����[�N��c|��Gv}j��EWZ���.D�T���a�S��wB�E��Ŭ��k�!�b�LOH�*�&�~l�z O��ɻ>�St���1�����믃�f!�g����{u4�:Fh.�\:��Wn�I�<���q�
�ii����3xm5ѴO\l.��;��l,�ԟ �~�޶=����������rEa;����A�M�B�)ud���`��܎V-In}q#�k?��ƐuAz�·p3�&q�E(Bƹuv������#I3�`I9��9�a�j���"?G���qV��CQ9�T�zR�!]�����
姓25��	�H]`'OJ�)�W$�5����������NԘ=@�������P���r���쉘Q���Tv��R]B��q�{�O��p%�*�8 3��4�.�K泖����P4��,��MIy�6�>�;�p���/Fp�EY��Z6�n���T���"�{�Ę�m.��\$�Q ��r��<Y}��������Qa��tn��g;��r�Ȏ��6I$� ��">!�p�o������L��\v;�ST�C�Q��QE5˒ߩ^a<����s�M�Z��ڞ���?������r���ɦ��-A�)Y�GB�_��2�ԡ�qE��8�O�zU��>�լh[�F�5��3��K�fC��݁.�ۀ�zd����������a����׎E�W|2+c�S�Z�`��m�0Q��33z���� q��a���(��T��������ʻm���{W�z.��5Lv�8��1�ن�(�_/����e�[�~���%�pjJF� !�Z����4��rS�i>�����N�h! �x-��u��&�l�����PK%+2%AL �Ѯ���DO�j��Gc�s�Τ3M?��+�� �g�91���� �a$ ��I�q�	��N/_۱�`��>��f�!��4�����`�񊴅.���9eB:46�f��=����t�x-Z��&Z2�:����p��	f�i���.�h%���ܛ�*m�q�d����b��ٗFԻ%�o����Z�#��?7���p �WUd�dj�D.�K~F��#���k(y"�юϬ?>��G�V ��.�B狺�T�0ȶù;(��]���WCWVh�H?�#�t�d�7	��n�����!Z��O���3xZ�gҸ�u�I�7���`٤�c�1��3��h���κ�����S��
��(^*kx2��twh�_3�n��$�T5��a���20�KD~������)WN�/f|�}�}�ޓ�S#(�f�
e֞�~���c��e �9����(�hXm���)%�R�K����h{ ���b�ȼg.��`�«$D�^��Y�@~`)�1}0�&M��p�&�pl���_�$][��FK�\G�Mga
�pO�D&�;u�������bJ�GHw�d�]�l��11a��i�r��h�1�TPQS�v�@,R[;����s�=�HF�=�zF�����vO[%�P�����V_��k��f�8��/�C��D�9h���*H/�Y���4��"�Vh�Wg�(��81,�]��0)�`���їg$���2ү;�nV����A]h�=H��DUl7�v`5��1�'8(CaUEȺ#��?�������9E*�W���(/`�|wr�@[�$-h|'P�Nu�KEty!J���|���0:��$G�o&ЋNY?N��lܶ�DE;+��*�E����x��6f��h(�2Kw	aI*�>^�wF�S弽:�/e<D �L�`1����������H�E w�oG:��3w�fb\��E�s�/8Uq~�J\~��YȂ�9U���Lv �J���l6���p始��w���?�~��+��P���*�4a�D�2��ê��x/�l��9�e��9AT�T�L_p��Ѯ�
�[q�g�Rf�[�E���]�$���$����=8��#*���4�(���J*%�/�����Q�N�1s�.�wL+�ԣ��������\�Zg��fXKcm���I7�sda�vp�=��M��4���[,
����$ݮ���/|�Y������sv\b{�����an���܍��#~�~`�/�'ml��혚d��R0${����T��B餪�����
f�HCD"U�!wċg�^�#@!7B�ʍM,�v�gY`% Z�˩k�bA�,�.w�U��?Bd+�b�Wg̖ �!��n���R���&2��&���g3�m$��"jI����p.������\Φb\G�mR�s\K�x}��q�t��תU}�
 �$�׶+^@�� �ssQ0��=����ClS��u�Rzq�N�z��7g�XJ�� �#���h盏ɿ��&U,�$��$;δ�������(�W&y��?�-4���awj�:sU:Yu?�$�~"ə�SŊ�A��0�x]��g[��<��d\#	��Q�E���N��:��S!����������2�Lj#��m�:`ʹ�UW�Յ�D��1��M_�R�~���b�@���Gth��k�v{q�����#�Do�� QYHv����<˲<f�:e����B����p���hb�񊓤��m�
�刭��2)��3�u�7c�,�q�o��5�5�����S�৊5�H@u�u��YQ�H����*j࠯��P|�R�]�nmpmH�K��lS��Z�
Р�6�U�Ҕe���x�O��Da�^H�40��PK�KnR��0�U�o3�O��F�[f���ͫ�Οu�W'W�-�?���X��ϰ������84���SgY>Σ�s��x��t�de6$�.s|f�����+��h��P�ۛ���F�4�=���m�������[5Yb�	#����1�z	rI)T���]�3�t�Eڃ��؀тjG�zo
w�g�D{�S뫸+�q��[�1ތ2=�E���8��@*���S�nm¾����AD���H�-ɕ��̬�/�d��:/�퍫�7�)�)�� E�Ś�w��i"X�#�Haæ�����I�d�\�߿��)�X:$)�l� k�0�Bd+>H)o���y�wM�\2`��\T#��B����歲
���8�3hrU�;���y��d%.�PT�]�qmn��)�i� ?$�x��~�+9.,]7��?��m&G!D��A�J�����<��+r�i���J�)��qyL%u�r�������=��1Zך�}:>�h�B����:�������s�]I���b��pӴ�D���#���Ԋa���/&��D8����A��ٟ��1xKDp"� ��6�~�TerB��7E�PI��HT���5�\�s��0�"[�`�_��@8J�O��38WK�ULaO���N���~���K�_�T��t¿������u��2>־N�q��W ѭU��m~ʀ�������ԫ�4��D���r��w�) R�?�I���bS�V��%XuýJ�}�L6�3�vG��yN�Ȃa3L���PmL�B �Y�߸3)ӏ�)^r��bq�^�'�qL���5z�B��ѹ��X�e���8A���>o�v.���Vh�)�'�M�{8p������b�!�E�_���}�����*eO�}j����&�5�TE�ޗ[>މ����u��N=%��ZM:S���M��ws�T�f�	��)�>��#i� Z��M��l�Gx}���B^hC�;�_41D���3#g���̱狰����N��0�-�ݨO�!IHSQM��j����o}x��ڻ�D}�1&�%���˛Q�r!n�H�nP�`]n�7"���/�������J�VpeRM��L50 -�~�%~���s�����I}�p��?n�VU�B]�e�Wj![q�!���曽ͺ��E�O�v�d)q�����|65r
g��X��^ԴؖU���<�p<K���d2�W1��[C���\ �9&�X2|�3��7i�+x]�w���9wq�]�-�0���Z��0qy�W��l!�k��BK��&]l�g烠>m���V�.�Z��y���F���<��40���ޘ������%��Bk��La�6�2�x��c)�.����)"���R��^X�>�T�����g��CU��=����&�Ҍx⾘0�W���<v%�Gr��˾�c�u��gI�1�˾17���I؛$�:HrԹ�%��E��+F�jM�!�]�y5�tm�<�5,�� �X氐��y��D8ص���&��oj�T�q��9��80��� P�#4����,O�iN{-A7��d���k�,��er%x��,JfV	�@vq�R ���_�)��Z��5I�I���lw���l�c�9r�Op����-t8��6�Z}Y���D��k��ʑ�(��W:� tΑ�-t��w�Q�V�M���;���)gO?����z�)(�nm�C2>|k�z/2��CZ�!Y\����2A�l�7LZ�!)���d���Wth�fv�P�:r�[�1zAGB\R�l,��-Y�S�@�oz��E��u��Bs*�)����0yh��\} ���-��MY��`���9i��8�w�����gz�b�WE�L�{V�76n�u.��G��a~�����mu�6�5�|�?��m+�Z����ܴTZO���O(�%"@I���{?PvܴۨF;�`����'[h�60��a�'�hV@�V���ay�@�E�wrk蒆n��K�s!��\ :AV_b!o7w��K���`Մj�҆F�ĵ���گ}=4R�������ӏ�gL�eE��|A��m>V��b����{V9�g��.�ψ�8��2MmKڈݫ#��gʟt�`�m� q����/ �;G54���ʆ�<:c;�5E�H� ���k�~|1Y�J;��o�t��M˜ʁ#�������YP�u��w.YO�qZ&�f�C䌣�����C�l#ڞw.R��|�Y�Ã��ޥD��G`�����bEd���[J_�%��
��,5Q�o�µ�(�=���ڸ��S<'Z������R��Ǣ��yuY(/��N[�"��kVæG��w`��2ۯ���Iһ� ����J���8��Ħ���#@ueޙ���;R�hk��|w5 �Ħ���cbum�5܋YқŢ�nʬ.4��̇�T����_@�	a��F�HG�=V,�]��6h�;���� gځe��0�'Ưg�������@-bx
�[9���F����pl��_��6�)�8��m�\W�S�C@ͨ��<u��J/#*�[�H�n_�7�7?�
p����З<I��+<7��eǫ7n�y������M��E _8�4����s����%���]��)v���X�ڲ�&R&�o�:�����ւhN���#Nog�η��h�M��D����L����|�6�xճD:�z�.�VEEcB-y�<
m);�$v'QO�e% �&'،��|2�ez8xL
��@5�� M
�����F�~���?n�cb�Aʀ�^^�x�������|R�0�Rb��%�����uKeD�b�9*4T�(��Q�=\):d���DV���
��8��ۘ�&e����/��ŜxJ�~�R�8<sz��%8
2-^�lۀ��)p̣@u�*^��.�2����b}n{f@�/x���0��d ���͠9`$*����s���f��|h�πly��p��b`U3�2�9�v��9�F��񙋬H��pU�󀲀6�X�^�/����ok�vڟ��"�+���^BtnP�,sF��1�%t�|IapG�)�j�eʐ;)E�Ԋ�6�ju.�n+��4萤-�������b�ڣw�qL��j�Ɇt ��V�Z��_ꆃm��*��㪀���M�;�z%'
�!�X�1Rs׺�z���޿~���:s��:�H�I��=��jtonׂ)8�.�!N��"\!/>��~�����H�|�rv�����w/r6U~� T��KSъܛ������l((,����9� �����j���� �{���|�86�wٗ?S����s���;-��~%�t���{��L�B`�+���p���R ɚw!��f�����_l�?�i\��iop�	��J��_9P�Q\�,��'��"�K��Q�/\�gF.��:Hcx�%��E����Kd�55]�v�% ~*�s�^sS�O p7e�c	��x=���O��� <��A�k�G��iTB�V������c�	H7�9�HסoHʤ!4����}\�&c0݃	5��KX �[޿]�0��O�y���\5�5H')��v%� �����Q����4s�*�#~or�lU�7�.N�
H)mHǌ� +�G��J��٢H[�ж�H?!mYÇ7����D��,\�!U�=���y�Sz��w%m��.�Ci�W2��ǭ�ѾǕUD����S���E���iKH���x)@Q����k�S�NDq�r�}=� �g}D������H�:�FG)�Qת��&@%��)��)���8,/�23��%τ��z=$���L���`�I�u
���m+9d�wş��;Ȣ�E�L%Q%�P����7t��~l����d�^�ʤ
��(�ptj3/d~�u#a
H���Rr�\�Q�ۈ�|<����j�J(y����z��a�C��+4jm?
jL��M]�$�:�Q���PfEOjt��[���BE��-�tl6:�r8[�S������k�x�P3"t�g�� u���j� y�?������ �T!�_ yW�G pMz�x7 �D��@t����;Ӻ"� �������e0�p�	��b��HX�)�.�B��0���W�g��q�7I�a�z%�0H,%]�G�ɉxB�.rY9���w��&eZ�s��T �g�a#����
�����+��	L`	7�ə�N1y.S��}��Y���?��)24_��jNR#D@v����I�Y��Z�6K�
��13��Sc��<|v��ķ�&�o��*�*p�[CC�.�N���;�W�[l��b����
f� �5zP�-�)v����z�<3�Nƽ�nYO��	�XB� �bq./��;��ӻ�^�n,�ns�z�t���h����A�,Uy#��L=���,��ত� �,�� Bk�-��e�Y;[����	>�-�p~��C�F������m���J=�8�^a@?���	�ڦ�q�{��"���Ҁ��Ed.��������Iι�TۑS��VI���04VNx�����Z�?X���?�$!�4��`U>��ezR��L}�r����<s�x�(�qs.��լ{�>���'�Cv�s���cO� �>�EM�mK2���E�H-�0	GA�?@���>/2[ڋ���M:���k�lH��ن���0ڀ�Ģvn�����;���t�lj��K��@ܼ��?}*OU� �����2n,��f�6�rq=lъ�u���|{��o���Ya9zp��ȸh��(�.��n�Q��p����~4�Op+w�'?�%�z�)d{���`�<^�G�k������hGKJ�
����?S���\�'A��O�f ��<}U&7,��Û,��?�P"@�F��-g�-]7
���j�*#?6��I���:G>�\8�ɠ�$��}i9PU�8X����
F����*�ԃ��nڧOz�՗�H�1�#\���>�|���i���n��<{-R�A�[ZD�3a\��# 7A�>T�A���4P��M��� =����cݸB��L�"�9��c&#�"��Շ��뜶3Qln3�1g��R n$��''��w�l[$P�-����U2~�5������g|�**����]��m)�g"���w���:�9T�&���lO^i/Gǘ�ݝ?��9ܗ�͵������@ۏ�Ƙ�;G{��Ѷ�z�Ub���WG�����6y�(^����(�%$'�C�p��u1U�d��5Y�0�/m`�b!o���%V����jf@
y�p;����F���?��G��2�8�Ip�~��B�$�K�5u�؇���8Ȏ��4K��z�V ax��#ەۑ�R7fe��tj�	1�X�IJ�%���}�˒����5=(�� ŅM��](?l������}B�i�Z�4�ϸ0�[��_&#�ꭾ�����أ�(h�r(��Ν�	�U�/%��v	���#�R ��
pr��U��`�������vL��pR�[ץE���!��f)�:��t'�}�,��P&z�}:�.�g�g�����6+���P1� ^^2W�y��hE�k����{y4��k��̶�ԋPV�s��g���AZ�@�m�$�v^��f�1k��v����J0�寇7��ۖ��̥��F ���A jTd����C�<
*#�]�5Z�Qza�I/�c�^���,�:gyu.1%+k1��r���wF�[�W$�������\�j����S���OƁ��F\	��������b�C5�t����?��&uR"I:r�ڮ��{�W��{�����E
���Bx�[Xn��ZH	'/�%�P��Q�˦����,U�˄��'��#�SWf�$�xN�ʬ���+�j2=�/�-S���vf��pK� ���@{ X�p0�0c���K�g{K�ε�P��t	���o4]��$�V$ �u���I
L�|�(�aNi���CN���l�+|_;��I8�``;	���$�ʺ���:��ӇK-R	��p&�9�Vo4nU�a�y��Z)�$S ���t�
���C7"����t��/-[��Dν,U�|Ȇ�TAPV�=�O���?Tէ�����N���3�M�?pD�z#"JF�2�8��=�oR�kc��r��2��l}뻭{��(-dlvP;1F���mI�z7�W��V���'�V��o��'3�f"]e��7��z��U>�[��
������{��Z�7m~��S��m�,�^;ˢpkY��[o���Rg��@�֞��k"�	i-JT�~�C+``� �ɜ+)���I2�3��	�����MyCX���hu�N�ސ�ㄒ��2_�u�#.D�� ���\���,}��Р�Á=�䛻1��{2�^w-%i���:���E#�R���4%��R��!ݭC��܋�TQ�|a�~)����Vꗤ�И�&`��S�fe/ ����%�h�O�xᡬ���/��G�`�{oTOcl�\Vfʜ�g�%rFHV������1�\1q��V}z��åE�9oq��⧀�����H��$i3?��6�(_E�(Ȣ���Ew7ή�Qy�
�tDO]��C5�/	�Fܐ����_j�+��|�� �q��$�H*6��*�E7��m�ֳގ��$8G�+����`?�@	/���>��~7c���[B?�X脹�x�z�&<_���b�D���9��Kǫ�u�Q�jD�<��g�N�dPT*��8����<��`�� �i��"NNpލ�>�����i�4a�#��X��4;?�q-���,�9��x������H��F��$���z�<�&�H �@��þ�*SQ �wJ}���Sz�����!��t+;�y�3��F��|�VΈ�*��|S�W^Z@��CNK)Ҹ�9|m7O0�;fw��0	��	�Q}�ki���P2٧��5Eh
�i�/ؼ\W�Ψ(�l�L�[v��p�!T����&m��XC���O���C������p=}+�c���]��w�}�|���j��.Os��Qp3��P���}��&H���M
?H։�U�{���ǰ���(_��t<�	߮ǐ���U!���j:�����@7S4C�\� ��nu�в��Ui��ϧi�3h��I�\�u6�)LK��2�L�� ����oZ�z4x
����d������aVZqh����F9d���tb4�(��[�څ5:c��ꖀ2���zg�������f��#�q^N�����ɏ[�s�C?��x@�p���+�����Vݲ}��C1���;�����k�H�ô���ͅ���`�2Xv�����hk���l�Zn)�ឰ��?��1A�ď�3�#���^H2C�g���p��TE�WD��;q���3}�NL��(ZX�(��I��;����S҇� �6��t��8Չ�p^��v2�Q�ɶ�	������F�7�2|e�X;Ͼ������9��awrZU�f�y\���nH��zW��]���Hs��!����G� _v�X��������ߵ������	k2 �ߦ�\���^�/��LAR��_�ܜjO$HM���g�0�4��:j~ܭ_��|���u�+��0(H�Q��!&������b�EG ���B@�᳐5ݩ��2��WT��^%Iw3�"鄜������`�B3©�:��TH��J<+Y<�Er����@}x�:�g�˕jS��q$k�����ǘO����&s�ps٘�pIL������~'�w�����\���K(�p���1l������vm� �.��F�a�Rf�ʟ]E�T�f��	�+�5�z�uj�/��Ax�}�L풇�"ʾ�i�����F��^v/=u��*2�̳nd�ՠ�r��[�O����ɾ!������?_�P�V��~��,�$.j�E�4�]ޤTk�qL��@��9�!4���h5��&�nڻE�EW��B�8ں�[��2�� ���Z`1U���z�q��M�1����Z���IB���4r��G�"�û���%6Se���Y?��5ad���&�΃^����;CSp�L��@�,�"ϲt� �g�W �ca�0!%<�io��������evB�l�����^Z��GH�9Aa���jzZ��	�V�Zj�
%	���b%���W�m?a�)���J5�EE\r+���d���S�����v���I%�K7k��hQ[�`����I!S��h��s���ccb����
�K���U���䃀�0E�+6�K��]Q�s�����nγ��Qe��J�ڬ5I����n6�0��͹�	��d`ʂ��i__�R�XN��l=��P�e�(2���Ŕz�D��d&n��V�Y���&j踑T�U���U(�w�w�Yo���Ȅ�#��=��1a�/G��.��cU�A�t��+&������ڏk^4�	V�Vɶ����w���.�B��8h��[$�,�"�������K��;Z^�EvgW9kň�N�w0���k͚�׃��^)z#�p�X�D.��%�Ef''&�|���פUO�5�,C�s��L����	ݟ�;�M�{��JBGo�++Z=��k�"���jڨ엇�.4��`]��~x�Z��κB�U�'����L�B)���&�Ct��)�_Rk$�i�9��31����Vu�Q�5U����/!����Xͦ�,��0�
�K�ҙ��Ց�a_Wi�o]�{t��.Lh��#���'Ѕ+,��B��vJ�
�.��p���{�v��k�>����$���z
�2���}�?M�ζ$AA�sNg�����Y%���] ��O��"8�gM�RUR>�F����`�s+P�e�ہu�n�� ��~�����}��W�݆�?�����A�3��fX��h($�����&��V����b��ޗ��Xq�RL�WOOmS>ͫ������X�86�D+V��POaL������o�O K���+�_������,���կ�:�����<>G0���Ա�D�Tܨ��A��O@�E���c��c>?���";	?����+�&0���ӂ3�u7��[2x��ͼ~����2p�	�5��Cs`g�� ���F��Ƀ&�?��cN��n���-����0x�P+!��y&�n��[���t�ن�'�PruC�۞���B�lp՝���e�欇��8�=�E��i�F����ѹ͇ݕP� G�����nn����;���S�}���-$����eo��㣉_��YO�i;�Q5+���Ew��V&��&��-m�A�=�>������{d�
{�@Ғ�U������,�����ya#SY�c�
�+9"v�.�R��������
E+=�V��o9u����̢s�T�c�Sk*z��"�9r�/��2�������Q�Y���?�����	�Ca��}�^�W/�h}㑪<��^��"^*NE�=D�T��YH]�Q<:�6�<�)�� r0P���*2B���^�N�<�ð"uW]Tz4��;�:�P'�<��O�~���Q�~$8N��'�8w���.���#ۦ�@�e�N�!*���z;�������V��-%��m�	T��f>:�v]CbYO2��&��܎���A<D@c�PW�jT���fz�1�cj�Qw�T4���s��([Ƣ�&),o�{1D��O{|�\�����T�/ƚ`��Y�J��-|WWvm�|iKwߗ�T��|���WM��#��+����ꜰW�~�q^@�];�P{כ���%P��v�6b�2}�O.Q�af��\A�QфY��!���C�Wf�� !��K�}��lm@�����uh5w�t.J�����:�K��?�2��)�u��8�YBt$�6Ē�s�� ��.}�23��!о��cs�� V�Bdm���!{���&ή�J1k���/�^�-��|FT��9�B�f���D�Gz��OP�P?�K�E�O]�%����2������':�i��ga�jes��]o!�uX$�NX\��U�\�.F�'�"�D��.�(�[E��	�����)N�ګۜ�U���&�s<� q6MzΦ#�J薼U�؛M���Jp���?�w�|����M���[���XZW8�5������\8�m=>���	�V�UG�o��ly'>�"L���ɇ7��ŵ�f-s�M�\�R�D�ɲ�L�3ڿo=��I����Y��"ob�@���.�>c-I�}� �L�3�^!�{�ϔ�M��{%�:���4��g�縰滤'pǭ��`/���*�אfEbcuI!6�B��z"�� ����=߈F�סW�R�4�1� ���	\�&Nc)"�Ę&��R��N���� �N��'+~ =�
�u%m�qީ����c�%�����$r� ;�����Sԡ!֫p7��7�]�1�#
��k�g�@���:��>��JF��R��2h�q㍒�� t�rD�g�㩮-/08��-���< ����Qs�2�H���*�1`*9����]��N���Wes9y[�����m=F���R�4��4�Hٍx������06%�a��K���p����)�~,Rk�Ev�Ǫ9 �}�s+囔�ղd/��q4&���C	���=�li���k	�/���u�'r�f܃ۑp�\h8MO&��%࿋�
�_��"���� �a�T$�P�~y��"rmۀ�`��I�6��K�.�aYE�˸�*�c��`P}����'�����c��w��$I�w�ڲ���ɹ�}�n4��F����Qɽ�|o�;�/.RXc`� f��$fJ�*j���g	��l1ﵫ�{�>�6~��a�ǹQ����X�H�����l�����Y���u���I�MP�G��Kwe���6�(�в�pJ��0�
ڬԥ����a�)6"W8�t���N�w�f�������>��	i'���5�Oh�2o
`BK��3���$��:D�p�u�v.5��G0���$���"�#�КE���fE>-٨���%Ew����tu�^�)�lJ��ޕ�g���L�P�s���46�����mG�8jM���Z����޲t?�V�,&8�����{:� Y�Q$I����$|v���$z�
���l�X���d��%���Ȝ���R_jep�NbqQ�BK)�UFon\bB�����b6[uۯ�s�L��}����5|H�+�?#�>#�-�e*̲Eе�BiW�@��
��y+��x��.�fr����!�foOb�&�������c�3�H8���&�Y�CE�Puk������f����-먾�ZRL�A��Uh���k� V�9����!���\�f��K�*��X_�9}���iC��6�QP�X�J9h��V\���ȉ��Yr��D'�)}l����Rքd�P�jD	j?�OD����Uu���2h?9��Q5O7vՒQ=Е�;��f��33��E^��޸4Q��P���'/DI~Dm�s�ɉ9`�z;��' 	"8�C�#"�-!#K��	�<�֯��Rq�$,���������ku���E$�L+�_8��&$mSF ^�T�]w�-331���6^0y��N�wc����KJ��r�����G?��]1�rJv��p@���,ᶽ�(��|4�Mߔ4� �Z�M�f���fFz�ч��'[����O^9]in0�j�!��S]��V�� U�S��O�������p4��8�&n�m�_NO��(�h���Rq�*E��lbu��tN���!T�t���e���Z�GPs��;�1��a���I���!�`��!|G`��o&Iʾϋa?�hB!���n���i�iEx0p�O��)E���iRїգy��qNɗn/c�17k�.�c�v2�Gl��D_�Dl[?���q9Ld�c8����|la�k ��H`MJ�c�)ny�K�ho+s�8�X��	R�7�27�\$
���`Μ�/hu���x�E6��s?\�Ѡ�+�j��Qd#�Ey�Thխ[��?�~���X�k/zvxMLq�N-���\��p[����uS�����8ы���;���ҫS�ѡ;rE�f4�́��Q�Q8�j��0�W��6M�0���i@�.�,o-��H�]���?z
8)��TZj�tJ��/U?�Z�wK"	��������=ŁKf��y�l�����oaf�8�'L�M�g��
�a�6����`_6�yER6j|}m)�Z�\m��3%ddJ;.)��>���B+���[K�3��'8R�<f���K+�N�O���Nހ2�甎�3��vx�/�4|(A�����V��@Ȋ	n�� �o���H��͕e���#�>�Ё�R����ؙ��;VԬ�)K!���]4E�y��9�����l�u�z�����aQ�y�3o���O���:\��$���8�<B�8���+_��c=���� &�-G0&jS�̴){`�)�hI�3b��$��/�\�J^Z�>�K�;C��q�n�zq��0 -Kߪ�����[�c3��E1Zws�;��F�g��̻M�i�Z���9���7�!R��H��gץ�/�T�ח3��0�2\�tI�Fvq���
iJZ��=6x����Άˊ��[WUS}�Q>)�j���dQ,����e�=��X�m�64��F�vM�;���lQ+��_�B��j"eގ��1��gގ��0�hW���4명5�)2���~����ت�%�M&�j)���߶(cᡢT�����Z���u�]�� �֚����t��|ՍU,_�U�g>	/�ML���^�>�x��撦���G�D�{�lp��H���^io��4��яL>�%V23����	�0l�Ԇ`�O���ր>�������}�۹�}��"ҵQ��C�3�l��<�pZ���^Lx��K���f���ys�q�@��ǻ�-˴I�ȥB�qIļ�1vkӶ�M<�'��3�oq�õ���;��3��껂�]��F�\VN��q@	)չ	����M�<X�2$�z����tF��Ӭ�7��.�1���H�!�Q�Kvޕv��U�'�m��v�cn � 1}z��ɥQݓ-Q#��\��Ez<��݇C}�~����.e��|G*چ���Ool��~���g��[����� ��+���n=��+�i)�ڳ}kN�E��`�D��Ű��0o� ��as'?��K6����U�:�-�����<X���N�+V�EV,��Ru/��V�at��g��r�R�v��w�<��;�]E���Nb���Xj"�ɬ�[>/�Z�S�m��1��ƣG����:���R�C� �燌]Bu�wİ��Y���6�-���zcp�x��2�僘�.�X�2�0�Z�ӊ+.�-�o��X�S9�`�/�z��z�I�wvG� oђ���H?Wa߳�˝��'�8{����i2X�k,W�/�	��#T�5щ�� �b���z�ֺ*�6Kk�_�f�������)�q������
L���8�Oҡ�-�5���Ό����T��u��|��.-d�A��������d'�n��	>ᏹ��;q����A���1@>����Y3Z���^��C4��G\�sY��2݂ޟ�$t;
m��fXp��"�Er[y�uV3���TT\��W-Gs4�ę�g���1.^_]Fv�c�v��c��z�u�r�a�N Dd�A��o%FMX��ܿ�Q��h	-~ݽ��@��~�NK� h�9�@��(�xb���~D�y���7J(9�"�]M-wh��s$dj�9L=�pŨ�?j^W��m��2�ƪ��\ݰ���u�^�Ip �/����q�nT�.�y0��s��d1:�9����&X(��Z[�n���_�+�����"�
�yo^�I�� �\���nz��^��6�����E�Ƙ��k��w>���1��k��I-�~���2���4nx�t�PG|_
���\vr�d�#���d�u�V��Y:MӠr��e�� 	�,����&�V�w�x�Bs�`��jU2k=�yP�8�`*�X��G�<2���vq��x�3�����t_k��Jݨ>�����A�`��tSi����{Qk�h^��UŔh΂w��f�i%p���U~RV�K����:�ٳ���mUkMm�5�w�7�� ����_�z�C�"�6^�DTqRU�q��>S�WW9e���q��r
�(�� h�d^����=���s��C�[ᶎ�s����_��v�Z,�_Q����F��]��-�%��n����:T�秛h޾�\��K^�m��\�S��ŚV����c�V�~�������\�4�_��i�&s5ؙ�Tt��-E �_���`V%�e�e��O�|&�M���3�p�H��tj��}GI����[�d"ꍙ>ѐ�*M�ࢷ:�8@DF��������o�!�DH)��O� .���	>bo��i�Y�a���Α+�x>�j�q�G{nK�<,��Tr�]�I�������5U��8X`zs9"#QFF3��VO��)������BFi>�����Y�]��]��z�,u�rc�����0�V.��>�H�04>Q$Z�zO�A��X�:�v�tF# �E�	��<�(�������ri������H�\]�+UQlĂ�#&	�y�������]��0e�=sN7�qEn�疹��6%��~�,@L,B_�Z����G��[=&��^>�?��yI�6~L�~��[;�.O���um!�乿��-����ꢞ����:�;�����,�.��~��f�m8O���{��qf��7��뛿���S���4)�	,(@������yfhCX�I�L���GE�\Nu�!®�j��mv�����m>Wf0ƈq��ݪ	k�Ě,���VV F�
�\#j.�* )چ:g����H�[�4rc��饙�Z�GQ&j_���l6��e������ ᣨ�|��VPҁL�g&�).��AAstH��~�ͬ��~��НXV0G%X�{���!H�m�'wI�pP�o|wNI����jt�Lc|h[����
��F�����}�Р�[1��>٥���f+XoX1��Aӑ��\\L��d�߁i�]xD1�iVu4��F`��;sx)�)��ָ�����`	ZlJ�����a�l���H�G#��y2N�p�|����/.�;�J�$��]\4�|��I�X�ބZ����9r�
T^�B%T��+���$�X���V���$����0X� >�� qO�����-E��n*����T3�.�@��C��`��ڋ�Kkr𩶙w)(`����Դӏ��C�l�J�	��ޮb�b�`�0x"�i���2�`u�F��2OSf�XG*�jE��U �O�����x�k}�{�N���r�j�v��|�9�n�85
�y-��,Nj,�y�����ԕMA^����?lE�����l6�眨;l����Sb� ����~��K�sd�XAU3,���9Ǣ�߸C�0s��]�����`tE�tR�˦�iP��sM���-a�әHK�ͫL�r1	�W�g��D���޹�k.q�zl�����pb��VJ*ɽ�-a��K_saerc��E����Y�)�TFf�0�t��Ibui�^2�tJ�`�[�,ֹ��Г���bo��6���Jdopb��A��G��:��AlI��a5W���s����hUߙ�2�;�j�19� ��B�C��^��	@����`���YoO���k~�.��/�qJ���J�2�ٕS�ջ�ݚؓ�%��qs���E�U����bI��0rF;!5�oi�֐��
�0�i󁬃�ET��L��omڎ����u΅�D��UWc��
�h�2L�0M]�|�QAOm�uRQ&��җgM��8����l�T8�E��.2	��i��\R9۞^E��W�X�-G���PW�!��?{�&�y4����2&�s���ݛ�5J�Q��;��U��R�Ґ�C�vv�V@ibqf'���$��,��Bt�!�����ݒ����k�g���`�8�_Hƌ"X�����>OӝW��ܼ�~z���?�pT����aӶ�gk}Me�Sy�B�*��tGN����i���:��^h�D�?���IǸ������b�uj*�D@��N���܁�Lt�T]����}�#t~���̕#~�'R}�^�W/緫p߈�:�����tg杫���A
�;����F錚���i+�i��Bnv�U�ՋE���%oЃ��<��yː����!P!�q*�@���y �Ps1]t����UlK⤶n.���(� �������D~��`��Q�-6z\+{�4�F���m�h<TF��Jk��<�ʑ����UW�V\������Y�����x��Geg��;�d?���sҲ�n����6��m��g$�-YdE��o��.P��E�p�����.��q(���T�#�Q� �K]F��R���T:-��S��b���y T�Ho^Ĭ�ºō�Eo�����"��^B�$�NXu���j�r@!�^���ӌ�&ii=fp�I.�	U��<x�u��O7�A���K:fW�+�#�� ۣ=JC�L��8 �v�����?�Y5��囥�K��*V��K��{�vY�?PG��C�E���y���5��'����sa��R�ĝ��nA1��G�ZL�a;ax�/���)eS\��A�	#�q����ŷ֍X�������gf|q��HF�
[��9�9���%%[Ѭ;�Mi��Ҽ�3�p�j`����	���8ݖT�$�"�͆fqB{���Y�;0���~��+�-:���U��4PR�	XLoh'Dr���m�w[+�D�����E�;��/�(���V�E�K�a��ĖC䑳�C�yx�� ��RQRT��!ߟr�V9�����G�،������לi����2rm�Ua:�բ�����*�B�'[8t�,��|��Q��L��ozYa��[/��E�)Db�l.�����z��b_�����mߑ��$�0��/u�4vK1����xq��+�ڲ>/��Lǆ�H��^�4"Q���T��7i/��>���/N���O2��Y-�ǻ�o��z��-#ί�ܪIh���Pl ,Q�F�k��Á�%��D�y���b�ʑN�&=�$7�B$��de��h�WaLo(MwS���M�24G�K�!��Z��Y�쿛��m�5 zؼ}� X�%#4�i�	x�ж�Z�R��S�����?�o*	��cո	�\p��T� ����7Ȇ�rV�E��3��p��Y��<3^�/褶�ӌf��؎�z%���y��Ex�=7��,�ʝF��N˼���
_�f�-y{�@av���x�[��Ÿ�` +��>�4��팗�u_w���)M܇P�Iz\� >����:m�3�쓹Dj0�	#b��۶E�އ�H���.���?
3�@�&$����7�|�D5����m��,�;f�x�u���m�2(E��c�x��P�ܙl�}�v�U�CO��H'} �A)�)����,$��Dش�oX�U�I.��%{<�`�`g6ial���u��h��$Z`bX���|Up)�,�R���"u	�\D�;��5��,�q+W��UR«'DJe�9e5�$�r�<�>�J��Ǎ�Wg�Zː������Ai9�Л1ǫ[]�i�%�Q"I�9�~cǞ�I�ݹ7<�~X'��_����P����=_3�Ǣ.�y��&߻(Y��ɕ�`�}�\ p��<�E�`T�6��@t�X����gj"� ����?���ɬ�ׂ)���P1<�zBtw�q/�����/.({\��)�|#�^�6*�JX�S�����]Ǧg�Yߺ�O�(H 1�KlSj7�K�g�_+�IyA�La�8�-�C�Ng�^�ϲ�61�o���s+c�ܕF�]����]L�D�&�j�ʘ+��p�8O�����R�79�@�t��os����ݕb�B=S������N��s-C IR��ͭ�5Һ@Vw餅!�Wi��Ė��p2�>e��"��'li�_jIA�����
�c��_��X�+hS�@����}-F��\�_U��UI����,a;	�A)j��e:��ր��+w�V>��Y����Qr0��lOH�� �*�|؈��1�Z���)"�RZ��H|T�!���	��e{�v��lD���΂,H���칧p���u߹���0^����}�<N��;˩(}:DJ��\��1�s��b Q.�<����l���aI�}a�4��@:��y��F}�l��#�4��(e�[�ԪzK3
�j�z��s�_�u����>�@��ԅF<̃w������W�蚮ܯ�SZ�������J��|f���� ��z*S��;���d�zw��Y�O?Ff>�#�Yr�����]�F��{�5XXl��A��\���&�<�G]n<Q���11���C��k���z�{����Kno�΃Bᄑ́���@�W,�����=O�����."��#�xN7��!���?�4�ie��J."��e>�#���<O�"�WG%�n�õ�(�2ض��V�U��� �KW䦱�p�� �+\h����O��%�0��2�n	&�9�b �+M
�`^`��5�m����\`s
��I��?�������Rg>��wn~sz����ݠ(����5�b[�Ѓd��M!��xp j/��珚���/_4����xy�6�p&��p�+'pF�'xE5�ܲaM��jl��uFkFO�f��ԅaPC��{�H���
�3��.bup�$m`� �����Y�bÜ��"�K���h���0��и5X#�e���1�1�aI%����R�M<��bT@��?~�#BŴ���xG�WCNF�$"�V���f�-�D9��g��{T����社>n�د��	����ŵ~�}i\A.�,�-�0����]^JB"�m!��֑3M8�>b7�_���i$o!_�I��ڟH�U���9翋�p	S�����тӴn�[-���̣��D�|���
�lMp2�B��\�<��왉)F�1�5�%6�w����?)��j�0!������а��v.|��܏�Y|�ݾu,+pgPB���[ȀLq]��j��w��:W�|a�1�Z2s���Q���&��Ő]��4�UW�+�l~tJZJ��y��~G��(��bF� ��*��Em�k���,�,ZX#K��;2��i�.0*����)�?N�R�t�����C�!(G
wdĿ�<��o3uv��E�����a]_�b�֍��-��f[�Ep.`N����Ug�A�E�	=7��^_�_�#JJ�L@i�?�B[�Z�Xl�`@��I����0�K��$d7�\$><md�˔�g���������n���{{\��z;����c=#��2H�-7'�TLd�g��e^�ܲ9:^�c����F��ƌ/jK2�ϊ������L�|��`�!�
>/���j�AN=�w�w��("gCJ=s���?�&�	�=�'eLmߴXK�>P���	A�+Ԇ��Q���Z��:�0�Yu�ry[�4�ÄS߂]邵�O�Ϟ '׹k&lÖ��*��%T�D4̯�0�Y��j�UF14��j�����S(����(��7۴��F"RL��V�u�������z����$�[���%@A���������Z�y�l�wO�5�-�  �����{""�w�&�h�<ꃃ��E�!��Տb}��v��2�$�I�1�PCC�F+J�ý�����4��N&��曃Գ�k��?�������@,?���G�0n�b~'��J�(oB�hB)���5�4cG�����nǌZ&V+�#AX�P�mp&t�u���}���Qn9�%�����F�	�pg��9VG�"מ�Jl�*�,��$h��!����&L��*Jg�=���|a/h�P�R@�x [%���B������氙�_ʻ�tK��q�Ggl�V9����
}�,�>Gk� M0}� f@�w�Ȣ�mJ,4ʻ��I�֏ï�^��sUI֎ �6@}#��� !T�&-Ņ��.���x�^���'툺	�9���ڠ��Q#���/gE��FvB|�7����G�F�뙔bŁRs�&��z�le3逶�+��C���HgN*�yf��G"�c+�)�u��B��\���l�n���D��Չ���~$��;����"�"?UM\Z��m�k��犊2���
���A?C�����Z��=%i��l�s־���bYY?i��j�D�M�����j٘h������K_�|�Z'֤?�T�y��-;�m����B�>R{˔4TBz`?�j*V�
�fcJ>��<��5w���Z����&��%H��+$�s�Q`�00�>�xB��N�Ԥ����!�� 4S7�a��*ЭkV�J�$��H�=\О�-gL#M���U��y�1�E�{���"�h1D��c�� ��5��Uw�?��Xd5��c�9;�12E7��2i�س��N�(	[�g0L�4��2�����xQɅ��;徎����R�蝀w+��8%�4�#f/e�!ڙ�X�CE�K/@F��ҡ<V�!/��ގD�E��i-�+�q�F9�T��3K�-�~��,���|�.����4U�-#��9�Z/�ɀ���+[!\5^B��K���q��f��~l舶��ޞ@�IM�r}��O��o�	��v]����gx�>t�l�Ue!��c#��(����c�r�l�L5�~�t�HY���G4!`V�������Abt���A��������d�N2<:ʪ���	��NP۲,�t�p�^&��&iП<V ���{��j˜��*Hq� ���v)��9�d��qM�*�@D�����O�Rgp��x�`Q�:�C������"�[��S���22��?���Z���T�1Ǉv���j��ک�ѱ%n*#Ɓ?�Hx�K��3'+�lx��;=���M|g�� {;}�k�v�q�n>D.E&Mw�3	����0�@�.]K���aC�<��կ�K�K,��d+���F��ȱ����b��U~7����>_5�/�T�m�a2�/���Y�e�&voN�Ӛs=$�oދ�~^V�D��Z��T�/ǟ�?)>M'�\jT�eF!��r
=p���n�ǉ�o�~T���h~���5��쑺R_1�Օu�.� �׏sʇ�(��Kv�BC��	M~k����aex�e���!J|̥HeR�����>�gl�nrح���I��M}�(���xLfy���(q�R+�Ѽ���g��7�~���P0�R��	� ���%J�/q'g�0���.�P���h��3ҋ�����q�vK=绍�u;���%4	��
nԲ�$vQ�B�)��!�\����<��}���R�H��/b��!��~`��,�b�5z�4>6�*4�Ml}�-˥�^��a��/�|��N;���Y#�����퉗 ��%i�����Θ��9my��~�:�Y�Ƀ7��tm�zlU[�Hk#��BO�xo��A�p�Y�8Q��AK4K���j*R|�$��8�hdc����r[�8�`�P4����<����>[h��e�|��N@>p���I��~����R/JW�<z�V�k6��1,鄃�u�J}��?����:�҃S��>"D�ƣ��_ۏn��ts�D>F���#��6�Ώ��T�0��ʙ�f�
juzoC�<�rP���_���Eڬ���}Լ�:���ɽ��	�P�u���2�E�Z}��� X�?����q���6+x�J!����� W���\�A���۰[{�N����	������8Ҹ
Ԃ�� A���m���K#��H���Y7�[��G!��!65�[�ȕ�H�%W�Z-�fȽO��i7�����&�?���5�����<�w�E9�oL������8/��l�5����m+p���'��S��d�zl�-�݁k��S�Z��V�HvԺW>$<l��ښ�s�B��b����tLs_M�O��}?vT�VDS� ��7�dv��kR(z�^\��1��mz�^�K�
���K�B=s������ ��Y9<c� {,�J���q���I
 �����@R?�)���[�,�C#X>z=�lZ��P)�5ef�:y]M	��d�~��t*������ \ZH2�r
�/�aG��M��*�8���[*�� U?�D�L�iN�̰ҔL���	ۀ�%�|R�|ȸ��Ym����? غ��(����!�� T�0�raX��k{�C"IvZ?GmX����2�r�aY'��&C��)��P6KC�N���+��Y9?����ҟ���m_G�])uW`����Wqm-���d.���KPE׾۵�Qﲡ�������Z�.�b��ruj�E��$�?�f10���Ǭ���M<�������a�+����o�vq���%^��`�/t�x�xKV�m�l�+ ��Ľ��r+Q�j�C���O������v�+�P�觟Mի�=}Ӄ═ ai��w��=k)i��IXeP��%�ϙ�/H����D��EI�� +�)���R]�1��JR���wPy+�Mmˀ��zک�7��o��R���5����Y�lί�jD��]�� [�AuyK��DZ�}�֧ʗ�.Y�H�`��;=��f�"8' ��z��I�I��j�D��qyMז]:���������Չrm�k����30�u+4	�́�;ش�IVӚ�뇙{3-X��Y8������s���F����G*��* x[[��y�b$���Q,4i�a8eI{2�3rfsÆ��,�x��d��2l�_�W�qg"���lF�ߧ3�"�������,g	D�6YGƦ��	Ux?�[��8��D��|��b�?���zS/r@[Q�%�.����QH��C�e���u�`a5&��ov<�Ǡ(�f�
o:��ۤ����Rb�̈́�V����z[���C:���?+�R�S��*U��ǽ"�*���om�� ��f7�K�x/=��đ}���ÜtN�c�a�_��v	�%g�����"'�o�oP�Z_*���P�{�q=� wt���Ba�Y��/�Ǉ�9�;g�� '��G��<����l�W�4�4��E�����x\{
"��A�c��J���Hz�xߟ�D��x�<\/pco�(�S%Dgۆ�؁�idpψ�J����2X�I{��\�<��Dm��N� gH�D���/!
_�x5�o1�֢��Rl9�h,��^�I塅���"�ٰp쯓RAb<���Z\π�J�w!s0A}�ɏH�q�,�2�0S�*���t5�W������~y0z��0��\lew|�ڣ>�
�8�l@���De�1?L0j�uLU��$@8R5��g�Jy����Ӑ�.���NR�朘4�l �2�yVTV�l|���f�
���cc���v~y���Ψ�PGZ�I�p��$�	�t*������ЩOF3&�'F̋���-�B��-�|ˑ�򢺽�w\�	T�>Kk	����0��B��tj����g����3��vZ0��4-�x�뒖~[{$RB�'�BV�Ks.E,����|2�N�ǝ9��hM�9�U]w��lq�a�8*[����������?��d�	n�H����D�n1x<��k����mP�S*���[��W��S����LuZNƩ����$W#�c؎D������BH6�KA���;ErұS���+àd��mV=H���㏗��;��	'-��yW|�I���fG�������ڡ|#ݠ����	�P�sG��� 7��
�$�Y���Ǿrڅy+�i:��sϷ�e���I>*{�/Q�[��%>����s6�1�X?�!G�#2����&�,3�]p`є������j�O���o��P񼱨^�V�NBT�˶Sh�����C |ξD��%�a�I�\�o�w��nm݇�r;�Yq5P0��:)QA�ͩ~WY�9�-`/����p�@a��#��������EA���	�wҜ�g�C���lH�	�+{�m1����?e��𺉃�
M��3��k��T��^�w$��	�����;�,�~��[�.q~�����B�j�ߢ��i�W+�1�'��c6M�ki��� ;��rX�7��K[�`��(���ʁ �>��K�����tiOGP�nJ\��ߠ<&��s��Y���_�d�����Fd����|����"GY��ݯ���l�fh^�a>��ˉb��]d}����ƈl�v�JE�[�,]8s�nx�6�|���(���4T�����dp ;�Pm<��l?���x��s6�NUxMA����-�w�r�6b*]�ȓ ��|�5��?�|���Xb;VRW�ʁ��+�`��<@�z�y��j�0������2���	a%C�+�?�3�vs�o��&[��L5��v׬��%�L?�ti���y������@r�B����k�C�Qģ��ٍw���� E��)�;����\ږ��C��\�tE���$Heҁ���D�X!:�lUE=A����*{_�$���Ԅ^���eB��
l�>�ٗ�ugt�}�c�u�wEʥ��(��QE�b��Dt9��PcEt�L%�&X�u��I���(#u�z�R�_�7�"6��[���@W���r��3T���HX�d ����:������P  ^��9�����n&��	�Xw�3-����q��!��~-�݊C�jS����/�����7�IL�XI/�ַI��Ց-n�;>�������M����+�����ߋ��:�@*Z����BTY,!�� aGQ�sB�)dʪ�b/"2��\����t5O�\� �?t��#�u�pX������#���>s�jh8(�o�f��m�aS���6�O�?�O�'����<]��x�G�b:'iv습����[*NHvN^�`����c��j	��MI��îk����RG��4�P�e��>��Gu�C��Wl5?)(c}0�WX�j��du�����um;咴w��G��<�eQ�+�Æ�a��x����wvmu�5<֓�T����
."C���Ύ�P�S�=Y�HQ�*��������ݘeO8p5$՘1��^ƫ���. �`�,����f>R�#C�,??����IW����R T0�2������ooxA�i��A~\�9d��H{`�.B�\[�5n�eV^��݁>�tFc���8�|�	{��?nwu�1М���tXX&F���Z2����W /�_����A�" ����SB���>�!��	����B�+lSŁp4�x������>��Ь�Sgr̍���zi�w�m~X��^� ��tf�?_�C�X�j�F&�95�E"��}��Ve:�
��ƀ́��;o��<������*[���M��j������	��ٱ�k���R��S���A%4�c&��l�d�?J)�v�V�>�%VN�~27�.1���iF��ʑ�`8�3��0��	��H�"�w� ���\&V��NX����{l���W��nq��~'F*����;~�E����n�����D�b���Ao��Μf��hVZ��L�H�!j���O�M�j�L�MN�z�8x�v��)j� �j���W�e��s��/��$p���l�V�k�-�^�_{���ڙҤ7Q^��u<����ב�菽����HB���d�^���ց����+>hz�IOgOG�0�n��@1����Y!��L�v-���������n�=����5��Jd�Ous7\��%|��ZXq�K��s��,�Hݪ��
�A�:�I��~�ZU�sp�[��A+J@# �|�Q��aWaLr������z���V!n��Y���
��&�G;m>�PictP�C(�&A�z�w��=���jƧ8s'�����%���Zt	t�_>��DH����jf%��������=BZθG�m��i�hs��TGxxĤhb#}�2O�5��(
�.y*̐B�,��D��p���b�4Sm���@{"`��g��߁���_�x}�Pv���Ƌ٨a�zð&��ʄ������4Z(�{�Vmބ�u��'n=|�c#l�n���0Z��3����1�y�ko;�B-q�01J}�'[ʲz�O��]�+s1���&N������p�ȯ��b.�x��;����������ap*#,!m�e>����84��];��(s�?m�u� �	�e�[�L["��r=�:�s����H��Y� ��{ o"j�|X�E	�s���j��$��}��E�^~5F�kTmWw�__�~]�K���1�A�����	�b%� ?T�*j�T�0���$^uG-�^7ȯ7��	��w/�hM6��]�v��u�.�}P�X#b<p1i��A�kϛ$�5e�uٔ�䉆 �C�V��*j���1&��s��d'YPs����s��t0�*�dNi잂�j0���(��x�QA���cF۠���ь����,�-�5��So��1,\͵���&������#��V���6~Y������UА�a���cT�'ŻU�3Z)�!4`�3���?/����@>(�$U�e�V����&�]�G�Ɲ�T���c���È[-���=�<L�p\}�� ��쨔�[w��n�D���2M#��	��:�X��U�tF�KZfJ�+���e���gÙ�R��
�`︊Xp`����I
�q��k�6�t���	������s��������?L�.��w�	|�LՋ
c��vL+9�^�k<Z>��!o�p9�����Ʌ�5�Tf���f ���\O~1i:Ӻ`�`��G,V�Ј�a��W#'\u�'C���[�/�8C�F4%/�.�U�WXHY�&�(�q�FR�o̫�[c�v�����'p}�7��s����ײ�d	��6х���;x:���3H-ө�?n#R([��R��26�kX
ʄ"n�K+2��d�,�1�랎c��H�L/�7���3�E�H�Mb�	k�ҵ���O_.di�Ì�wkSi�ST톸vh'��K��*M>"�[��`H(!��#;��t!�~��c�Gf�	T�V1@��{:6���xd��/W#�8���V��iP����� ��$��dr>=\�4ޝ��[M���E��Q�L��ۥ��N�����a<e�=���b0�HɂV^޻��bC�B���$|������O�k�����P�/���H$ &��H~�Y��i)��°z#6r��nP�7r
st����Ĩ+�2�vV-ޜ��w�kѬD��ߴLx&4���מ����8���=��"mn��譗HK��8�c����`��f�t���opDc}�-��9�\�D�h�<4hl���Z��)ݱD�^��Hf�eY82����ϤNƂ�pD�k �/+�|}Ȍ�u�g*q�%��T��0����H��S�!C�ÞZ4n
~�_���k
��A����5�[h��P�'��@�|(:�:T=���l9���d&u�$òVmW.֓���0#7|hA������K�P����q�KV 7�Q(>�(���:�"�p��Q�����u��mAC4L����>b�-T�GϏR����B3������%�3��MT��N9������/�Ǌ��*�G��.\T�����*OH<�$�����j�q��W�e ,�C_�|�Bik�
F]�L��5��dQYp�@�ƙ�Rߋ��0�YT�����/���@��w�� []-�~E	�pm-���g��]9n�`æ+�T����>�x`�ă#'LQ?�C�\!�
�&41c���:iz3U|&Y8>q�ߜ��ͱҭ�ɬ7EN��؂<���NINLY��yp���;���
���?5	�m��R��K�08!{W�������2J� .��e�p�ߏ�oP޶a|K�����'�A��ə��+Ч���7;��W�x�9%�e��H}�R���Ot6�%��bQ�4J���jW'	�wf��@�d݌��ǿܹ�9��x�O]-��~`	��;�$�0݉w5]qJ�E])��lNa�=D�6�x�,T�l����G�P�!����x�|�
�f�6�>U�qO�a7%,��ϓY�������v�O[S�+����oD���=�.n�,��W���AuL�؝�g%�Uoe�&�2�����k֤lb$Es#AŶ��쒔ƺ�q+���O ��U�@��A��;7S:���{=���W��x�/��*�1�SP�������!_}�-OB%uO#�7����k�i��4��o�ߒQ@3ɐL������>�`!v�Ye�9�1f.k�q��}E[��v%�uK�^\xm�M��^Rs�5B��lZ��������Щ�����Rq�+�/�\(.�;t��'�Q�0l	$A�]��+-��vҲ�h)Y� c:zl��a��Df��c��>Ș���H%��0:x��<4k����w��;��e�x��ˇ[
�v��zE�0I:9���bC��r���b(M.�1e^��*��Kx�8��_CgE��?.��_�T�>d�dl2�~-{gm�4GG�gz3����r(��29��G�rb?6��7� �3�<Z"vjs�Uq��r��d��X=p�������W���xP���Q��s	2�����j�,Z[[!]��m?|~��
P�}�S��Ρ�0�r���>��#sqk8�&�pfՐ4C��^��s)7PŢB�����>�hrm+j�J��Ԇy�<�Xn��O�D���KkE�rd��� +�`��h���q�x_����)C�s��Y�����6斛��h �v�j�q��	h��F��<)����
��woM?�&�l����Ra�bYGH��qS�����y�����`�s�{�P�˥{^^�v*㤞�N.��Z�.�d�2Q�$i"�1q5&�Y0D�
��R\#x}eK�Z�zv����2��;��Y�('�M�R|���A�H_��z�G���_��UI3y?�s	���_li38�d�] ��/i���E�ڥ.|L�P�0�L�����࢖���"�Ɯ���q���x��W��Z��_�HZ�*�ݏS�x��u�=wz����~�x�_�3`5Gb�7XP3��$�A�y�,�mK�4�<� 8C�q�T��8��f2|�^o�l��y����MG�I&$o A��p�2�w��_atU�v�$�#&
��JqǺ�(���F����>4��+d����h�������I8�����5H��::�Շ2�\�&�řlV���2�%�	y+���>����־LI+~�P��EY�L�/����E�}3����	<���R��&�B�Z���%���ON��3$�����RSg޼z�ggf���e�@�6�}TZ��FfC!b���Fd���1�#�;4��/��9ɶ�ﯕJ�q�q+�'�v�Bn%9B������lضT:�0}�`���k���;ŗ�np�U1E�tKϱ�T��-%6�W��Om�54��|0N�Q��Â�M~��]����*r���:)��Ǖ����N�����Kv�'b�a��-�5o��?s[!0.��#�(�}���m#44ިl�Q4���tV��J���e������:f�.�t�><^I��f?VcX$�W�~Y��ɴ����B��&:*��F��K�<
�\�'����J�;D(������h��{dv^�}�α�K�MQ�[h�4�x5�w��#�/�va6�5��ʚ���Z-�>��JA{lq?rK�^A���G�����K�$h�U��(���B�����Wa��ID�a��2j%*�3�'�-rU�!����̪����j��O$�.�Xؙ�D_�A�~M�R�z)��l�m�Ce����̰Z^W��!�Gf<,������x.�N���'�^.������a�P~O�� �8>�*���`��e�L�3`�ﶤ�����I/2��L�rEN��!M	�ȍ谴�	����z`뛛���kjM����ȁ �<�"f	�z��_> ��Z~�2����&Y@���s�X���Cϔ~�Hs�1Y�g	�^��icN*;�Ëo���<U���b^cg^�EN�v�+?�_/�ݹ�Q�;��L��b5W/O�as��<QG� ��E����&�ܙ(1��;��0��J��]��+��kr�ޒ9�F�����7�d���D/��=W��`��2��H+��SdKY{;O��0�u�Ѣ"�i��#Mۜ^سu�� �-�J�ב�T����@A�uy�(�	�m3{��&u55��7s^I��Ni��<��b�Е���h�L^���Ov��ԭ;2����b�����D�~B��^_�++HK�l�<'ٲw�K��D|���d��I��9��:�b �;h;�Y��C.�\l��sUx�J�!k~,����Ko���z�NW�['�1b?����,�"���_r{Ъi�@ ��\����_Y�����=���Oǫ�k�u��$7 ��H�Mx�<:$F͚�/�G=8ȦϑK � �.��B>���%��8z]���6I��?m9�u�ې6��5l@���%}x+(׬��؜���@Us��������=�0���I1=b�z-��� ���p?�N`F����w+{��op?��i��y�sdS_	ZS~�Cb��3��N�ŭ���%�\ā>�ȱ��'�ʌ"�,�F/j3���yz�E�H�9>�k�0�%���ڷ���ߑX�m<_��hu�?��&-�r+��[K�'�\�����@*���-l�x�Ev� A>���M��M�L��13�I���T��$��r�� (%�G�װ�Ō�gPI�`@�&ö��_������>ݬ��:���O�!6˻��n���D�c��W@m:ݥ���D��RuT�#��'tI(B�4L ���#2z�k����0�Tb��BM�6p:3s"�h�J�T����E_�g�� �Z�jc�`T�-� ^� �V�3��*���?t&�vy��p��1����٥~�0Wڰ�N�+|r�Du�}I��5�V-2t]Rjߣ��[��6-iV'�L<�~�@�ț^��P��%U��(cs-�u��>��C�K�@��Λ۾C44��Wp��Z����R�#P5V1��7fK����n[72'$�z���i��/K �~��ه�)妠K}!�8/�,�\�2˽ 0�s��H4G�m����}|\$[1fV��|����.��8p���sխ��e�F1/���'l����<��y��υ ����㳚�.xµ�j�c.�Ne�o�8���z��tY�y���e��Rw���k��,Dc�����E�d�M��c�aљ��8]��c��䯯�rز��c�5��9�H�7(�*�td��<
�f��#y"��)Lc�x|���ʦ2r˦��z+ӡ��	T��ޙ'n�5�QO�!��4z�p�����3�͟T��I��������w��q�<�k_�D��z�� �i�I�)��>K=�}[X-����M������H��4qaQ_�l/w��Z�6�K�Bg+�s� �N��z�+L��K�J����ƥ����k� :���D<H�l����2 /��Ph�w�����2�<x@�'׋���ј�V7�/�m���d�"$4_����;.��zJ��p)闐%*��������l�%Tww���H[p*��$\�����Hf��U�llΣ�ha)��+�r�nKH�1�x�*��?
2��{B��i�3-���'Q-�i)BEx�4VU�; ���Ѽ� ���徇���+OLt�}�]® ��D1�r�9�������g����bM��>Ŵ� B�n�]�sj���<	�1�q���J: �|�=�q���`�SI���z||��/��� �v~���X��3h��\f��Ѿ�1T��hg�9��r��D�� H�����
������y�Y��c�����ٗ�Z6&�}r��C���n��*A�0D���?��٣w��l��ŢF\�����)|�~x8���"E��6iW�x��vv%P35��� �Yb���~���=�۞�JJU�A-|����.����V�;�>乆�\�N��G6��}�ʇ[�u��G��:�n9��;�z��/�7�ʷ|u�C~���=zw*�o}F�Յe����"�����X�|���O�H�`#���Jc�pᗙ�ƶ~g+L�d�ۃ�5k��}��I���K��k�B���ń���V��N��*����.��6H"CѼ��X�w�=~9��]B���c|(�A@.ɪ�[�:����,�cY7�}��:�S�<X��� |�m:9�rK�ډ!��g6�
���km�C��8��
-�斬�a���t�誙��=��U�hc"��l�h��k��@ӑ�E�ˠ?��5�ОH�ױ�;g��A��nf7��������|�7Q���������uon�m�Ȯ�n�7� ���6};�ᎅ�����aG4l�sH+��w�����:t��$vQ#����� ��:1a�~dxE�6W�V�q�\?��P���Z�eg��TS��Gxn����in��J��R{�C4�
C�>��{�=����Sj�N��Ҁq�J��o(�ؖ���Lf���.sC�I���o0���j&�/�rnv�̈�s.�9 ��im��.bs>P�(@!  ���G�`
��?�����2ʦD�E�ۙ��3"�d��e����_@�����Y�4��zwh����pG��U��+�����Nn[C�X/����f�S�_�:�2�y�lG^Hm�9��0z���Z��,�~j��{^T��_��Q7tv�����le�h���ң��|�0%_urt���2J�_#7�>MhA�Ka����u�/1�+ҁﳻ)�O� k�fN�	~���M�O(A�Z�����p�W�����!�b�6P��׋P��T�Q��B��;(BxT�;�&�;�"��
�Μ|Qᶺ$���%���!��Y S��3��\o���};�4H�|����:.f/���S� �ɋ����J����-��c���|Ks��`���>�f���j��%���	�j�g����Z�o���
��R�̾X�`ΐM�]�8Z<��G��Hwj�}���ݳY����/G�9���[1�5t9�C_F陝��m}���	4*���Z�z*s71���h�ݓ/��{T]���l/���a�ŏ,H��Oꏗ�6Hjċ���菺��v���R�|�����$m����F�h+oX��ݓRBv���
��C�n��C�Ic[i���zZ�	�#�)�-��3"oIWC�YKpQ���#nmF έ}�����c�An��Bs=>�b@� M�$fVx��\HT�{U��,Z��ʲRq�!���~u�y��׼E�#�|
s�1���Y��dl짜V�\�j��A0����31/���\�b:�;�\K�����Cz�:����O��-��o<�;�:�H����������I��D=�RJ�=a�m��]�F� ZB��tɎ^�@�l`ފ
5�g���y�0���`�[��M
M����s2�õw����e?�@�K:m��ҳ��(�b�v�/F�,LO:������i���Ā�U{k8G@����;^s�x��?#$Nw�N������$	m�%m����7�yE�e�)Khddͣ���<"YhoV��]T�$P{RL��v�>v���޵{��1=����-��Rܾ����E����/^E�e볫�(�y����$��Ŋ#u�	� $���2W�´��,`�x��:���@Ǌ�s�Œ�xkǾ��2WAr�������c��^x�F��2�����)�D�v�t��av�S�'�����73�%��y�HMpi+�^�I�k�����x~��oE�g���v� �6RU+�H�DLT>�Q\(3eN��޻���� RZ����²�]P��F�w`v-�e8��<��wf��EȲ:?�/�P�1���G�SK�Ϊ4	���gٰˠC��@���%��sj��'��!�Qt����D"��];�0Ł�c�jE��%8��)�%�_�\ؐ�憱��i��>�K_�e����=;A5�o�D�����\cdWuညI?�zVCpA��5ͧ�AH�S�oR;U�+Y�	�?Q+_�	$��J-�q��~H6��/2̥fMTT�¹5�\2^��|`�8�ܩ�2����J��@Q�j��Ȳ6[,���M�MI	���s/��)l�WW��Jby���\e�ڴ�v�/i���O�٠ia^&BC��If��9�Xp��~�o�|-"�1Z,m&rS�<�r&x�Y��S��[5ҷ�B<��s�k)�\��4.?[��	w��
qr5X�YbD��O�(��ܼQ�!?)���;gc���֍���z_@u����m+s���ӧ���B�ggP(����l���x�ћ� OJ�	�v��������Y_`�3�)E��Z�Q7�3Ո|�����$9�O���OYKQ}Q`^Ua�����N*�8�o{�&����C�K����G"�2,����}�.2�.��^�{�����y�7��u��\-I��L-[ƻ��6�6��r�~T�7�O�l���aV�l�}���P��!�ʣ��$�)���(&ۊ��Y4�#��&�J�*
1��2�cetD��������q!���2�n�JKl
8��S��(�8եw�ݽ�7qٌe���j�'�}D���W*����W��p�U�8��mR{>�)T��&��v5���"�w���ܨ ��!}B�+�Z�|���3�����XI���&$ 6��h��S���9���;�x#��} ��o�ּR}[p���l�~"�f���G)A7aLW p����d��� ����g�-�jS�`;��Kڪdf<��5��y�y�E���/z cmz�J[�&�H��Ĉ�@՚��R�-GM������v���I��w撣B�&(%�v��(��UTM;]Q����U�Y6O+�<�m����U���h
�Z2��úX����TY�b#ݹ��r^�&?.{� Z�9В:$2��[PS+�m)h���+����Soz�]��b�.�2[0IaH	��A��?�?��K�׆���(�[H���G���}IM�ev�l���\�T���N�Oւ���\~�	ޖ�ϝ��6��]�g���I7���5L���w�U�S?��boH�_�(���T���/�71o�~�>�Δ�|0_5t�R��`1����h�=s�hJ�^Rף�i����6�i������]���R?��巐���o?4ЅvAǗ���?����/�{)]e����eA�zӣ.om1X�����Ã}rK�ǡj��M-�Ĥf�c�E�5G����9�w�3�Ϭ�Z�����J#pw����������%�`!74)<������� h7(�?n���Ij����&�t4�n>�lM��PT9�,R�,|+�c�۝tӥ�Zֻ�:��c�Is��%ޫ��mglSꂷ��F����d3�b �Z���lY�Į; ���� j|5��0iUq�W����}iR���؞*�
^�Vc��H*�瘟�Tp_AVo���(Z�,�D|ۭ�~�}kK[�X�2	�v����+׾H�A�֊)��`rl���/b�/�E-����� ��)���S�u�(S�j&t_��!H�����ԟ���Kz+�x�)�"��8wp����56�Q���>��m��d��a�j ����ҟ�[3/�Q&}�%��Ho�T��(��K˙Kx.r�J���It}�:�yD�	���$S�Xi_3�D�m��ӗ�
���%��Ę�i%s\������7���O��ۨ}�%(yKi���8�?��*��� >!T��~a,�k�[�S�Q�S���;�,M^p�+�Y�L�>��!>���ƹ�-!��|^pELd~���c��|�VT,�.K���?K0�f,�G1�w��ܴW/HEm���R�r�H�k՘#��s-̞`���JȤ��k�o��`�Ǔфqa�e�'�-�G̤��7��7^���	5������>D��2RW�Qkw����m4i����v@��p�f�&�:��%��
yDN:n ��ah��+���f����O��N�kk�?cP���/�#�0��yc|����/��Q� +Gs�t��'�L����O%�0������X�� Ux�h�g:y��?��34O��p�D� )L;��d��3�=}]adM��v�;��b���-Si���܋��^�9������m�f"��GOn�2��yr�4��e߉�Q�ΔgA��Eik��¯�B��0�� ��R���>�p��e��t�����˹Zr����:�+�Q�]��&�Y�9d�o�
ɒ�u�-od�1	M<,C	�P���v�W����.5+ERs�j��3������L.���5ط^ǉϾ5BJ���/�9���Z٬Dn~1�ٜr��%텢��ES2�-�E�Z��H�⺌Zy��>�M~Ix��F�GJ�5�H.��m(E1�ZZ��l�Ue�l9�S�G��	⩨
|�䚏�n��j�����t�Wħ�i��z>��@DQ�í �����TQ����?l�(�q��������u�tre�i4M�e���{�?����s�o�����M4?ƶBXAM��2�U�F�h�U2�����5�n���!
{�U4�B@@���X��^�Ӊ_��Y6j�L"�WA����| /�֐�>����x3�@�1<���0�{��.P�x$��J���(��.�P��=����Wy���Wۓ��X���j|$�;��C�N�w�=9�ڴ|�E��\�W�H}���!����xЙ���m2�xl2�U�=e�Ʃ�"��;���#0 ��%<��΍$4��'ί��+D��	�;v+���"����ˍA9�Ei�Y��w�(f�(�bi�`$V�^�1��C��K+��W;��6�W��9(^#<�k��{�s�_,H:K���fʗVV��X[�����o�L�#V_(~��rG�w�@ʿܶ��R��o�E0�~����(m�:M���2�- �X! ��Sakp����� �0,����|h\9��y|�{��#"A�~����-ԲT�I_4���~U���VQY؄OzOK�J���y�v:Q$$�v�@%f�χ9�[~D-�d�Pe����\�;����~���a�=�U�X������yUh*�sD|�DI���$P%u���9"ǭ�9��R�g�h�x (����Х�5�Ĩ/��'�3����Sf�z'm��
 �e�ͤƦ��^�E�P�$�B���*�������>���54���^=�D*��m���h[��E�����'�E�)h����U�����"��d�Ì!O�99�%섽��so�O)����p ����H���ok�т69Td�gqJi3��?�� ���|4?��/�x�=V��#�7������X�+]��u�]:r�f��DT<�0��*��Q�}sҒ��;E���g�l�-V�	?�;��Tsx�ֆ���P\i#���lxhG�(Q+ +�;&�S߇�Sl�vkJ2��,�Q9��ݪՌ���c�ST36��U{k庢�l��%3���O��j�/\�4��� ��a`��� �<�E��{��S�Rɴ�}qB�;k��)(��B"���0T���-΀�tpC���@`v���J|��&��jQ,����!�-$$�7yV7������nqK�*��PK`� ��mb"�T�V�������B�M���TS�/<N]�T}���pP��I��	!�\���ޠ�s��8g��"�:(*��GEo�������������B��n`�q��s�s5d	�Wt�ax���/I1�[K8��aa�I�EӢC�tvCߩ|܍ь$PL���VY�(����\k��ig�Ck���g�/�S�t��O�� n���f��^#���?�p	�{蚇��șֽV�i�nJG��SFguvl(}�˯¢�P��&��$Jc�t�����ļ=*�⨙���J+o~�����(�2��q��r�6���MBf2�oPiG���*������r-W+�m��v
p+�H$;�&EusC�3���R:�B��g ��b�
�f��I�ķB��ӹ��CIOr�A�W��O�q`��<��eݨ�hC��($��R���*
u�b%pJ�jZ�ZtG�M��"[�b���c�(�ڄ%�{���b����V\6��<Қ�����P��RS�U8�(c�Kц��&<�5�o�w;��<�Z��Pn�U���;K����Q�T��&���яj�$�vD�x㞥��U	��Q�);&Tw��h�g�"�`h�[k�R<��PW��H6t���j����Q0|. ��������-���a�i�|Z����z9z��Mq�@�]@���D��}�ذ�F��d�14�=a��n��D���	��"�!q8 J4�	?z��e0`�J��ͦ���0�Z�?Z�ګ#�]T���*��_�Z�ɕ�Q��l�����Y7m��9!���mpo�>��(�@`X-�yNwe��r���~��&m�"��y,��g˷/�vq/���HG�I�Hî�ICՆQp��)��n9Rߊ��׎RM1[��9��`,�2
Q�C����Ch.h.��_fl�! �#�Ѽmi�;od� 9q8��q�v��+�9������A�.]A�s�!����e�:�5�Ҟ^�Qe�
�a8�>��AԿ�ec��9�Z��!}t�3$/��Z�mKa���?jQ�"��_��|6c ސ�����]z�*�y�u)��U�؊8�W�l]�Ӓ���Խ�i�Lf��'[�T3�
���, 6X �����q��lƾ��i��,��d��qk@qUɷ�q�m��:�_P�˱�ϺV�{�5!����j������ ǽ�ꮼg�z�zb0V\[K�=�3:Y���S(,��>�
븰����Cx��%��߯]	Z'�$���fOE=���ZDxH��j�3��sM捴�����l����nJ�}�:vFO08+���`��2�C2�*�A�% ��RE%�e�ks"�մ6�\��R�����"�U#�(P_�b�$�~W��G!�tC1�Q����SЛ!ݹ|��5�Ԙ*g��E��� Leͺ�	��6�#�ň����g[���:����<.tg��p0姒����&�nFn-�f8�ӡi�"l)2�;�����,ס]-t�b�4e�u��D̕�]���o=�C� ��AVQ=Ԃ�/�%F��q�I$ #h�⿠��'莨SL�$��6ݚ���5��5���i7ޒ��G<�d��bp#�c�ɬ�~!�ѡ#���������7���I60Th������ʂ5�aE�bP ��8,�7�TE�du����ө��c͙؋w����I�܋ń_yp�Sֻ�$n�CK�g���趰y�a�%�k��u�5�r?ӌt�F����U��(	�]��$ GLa\��Jؓ2(�􃏉Y����
m{�A#�HP���)X��	1�O!��N;[!ڕ�����M�Y����t`oǺ��k�?�GQ">��FǓ�-���9�� ~�N� ?3堡��ih�S�c�w�>��տ��*T����	.���,�	����&l�3Z��lΝ�7:��q�n�?j܎j������>��nyO����7h���`�&<q$��!*�����ٺ��?�t|¹�bt�S(�ꨉ�ɥ���������@����+�����&�4�G�t����W��i�s��Xj���!w�����F��S^���*].���kw�����tAZYb�n�%��dx��`��V1N��؛����8������
s�1�+�*~P�ߪ��@�̞�7�m����U��7ڈ���)L6�e�|o��a�xa� 4i%�J/���w�c���k���_�9���A!4�پ�:�}s��*ur+����E�� ]�"�[��G��q?}�!�ȱ.�8�?�9���S� ��oc�,���k���7ֆ�\ףO�Y\���XԤ;L�e�zj�'y�S��0��D�5����g����b;F@�����팪�{�V��R+J��%~8���R �bj6Li�/����^6���`a�g%/"�/6����PV��7Fǩ�n�40�0#��gU˩�yEg�Ls�$-�Z�RZ�5,�{��p�s��:.���*��$9f���@��!����tγM��9�M��,`�a�c9���[������x��L��&�#^[>�{�z`K3��A���S+(��q�>ws����BU�}�u��Qܭ���|��
���Y��O�zW<��ph͑}5�T��	T�_:KnR�!'��m_
Jt��ڝ�D�s���Uٮm�L��U�HL8�$�!���eR����A�]g�s�G:�{�r
�S>=K̋�]��Me��;�`Oo���out��VYP��R�����I�ܩ~���!�HXgx�<Vi��ʀ��M�FQF.\�oA{����p���.�C.��t;��c�dDnJ-�J��G�6�Kt�EX��c�5��S��}�v�b
_>I�j*HD��n�ڒ_<0���������u¶J�jLεb���yrq���X�����ԴP�+2�����	�X�k�F�T3���Pb+���(�ٺ%w�C�E������J�!�K���mu��,�pu8����B��g���m	���
�>���&��8_��U��5����<�����ˆ/3�Ϥ��͈NCW�%��b��fC��h���,rv�{3������L#��(z��t�����r���S�~_"� �w��'$|%����"��뚱bԔQ�*Ǽ�ݫ��i����x5���Lt�1>.!�b*�����j�ko�Vߜ�|5��.
?:��Wu�u��[�Z�
3;	�����s{�$������+��"v��~f�����%�}9c~���s/�V_N��
v�m)!a�?y�kl�=����7��Ot=��U.����ȸ���tE/���.�.>�d�t(�̓���yh>A=� $ .�Ч�d:L��
�k� ��J�~�Q��5��n�K�I�t��d�R����S�Y�F��K�Z��*n}�C`u�l�.iAy#�l�<��@����C+ܼ
)���Ə���c�e�O|�օL�;-A�e�FST�O�Ȉ�4�Lt�'�H×�5_��qX׈�ӵ%�SJK<H&���Nd����SZ�;T�e�D��-VW{n6]ۻ*v����{wC6wL�ӯU��<D�V����J��j��l��"ȋH��Bbؕ�w���FN,�*nA#w*TŐ�]:�a���DA�kǃu�*����4�M������V�]��8��y��j`�;kW9[ڃ�9�#�.�3	p�8��{���@��(aN��)Nh���mWħ�����뎑��sUy��R��r�KI�X3��y��*Jd��c�� �ܗ�mA��S�k
�Ľ�Қ�PBz/��� �5��f v���ӱ��>#��D�����,gsr޳���N��)F�UAD+��W6�d�Ñlpe�i��+�@��o���ߥB$ɩ:ljK��A�E�S}��Y;s��o�涷k�SD.5�dK�}����=&�Ϟ}#K�:Vh dc�����wH��q�#?Cw���H76��R��g��(l$_�ir�>-~8�UҔ���7����Up��ԡ^(�µ�i�jcK���b���6%n�E��uw����j7cx��	ي�yz��jzR����)�P%����}�ç+��;�Tn>Sn�OB^N���j1�ޤ]�P�bl�Vn�]��3��w������k2�Bd�o�W�$|���A���Y����p����)�!��'L�&������f�i�c#����/X&�(m
����	{g�_�����9���%~]��2&�X}�0E�F�P��!�g��Q6o' ��h�n�+��_W����[�oȦ7���1sk�@��Y���p�rB�Ϻ�R�w�F�2h�=�t(�j~;���A�-�9���LkB9������g�ˆü�3^}}���>t����wq�����:����V��:g`x{hlFK}��1���:e�>�u�vT<.�6��C�
��J��_e������%�.޾��J��m9FLL�U.��4�����SPqPM���������v4�a9��=FY?,p�(#O����b(`(i�XvɅ#���t{��L�c!�G�c4�"2RZ:u˃j~V�T���4�W��^X��|��q�cU�9��7�6�`��G��e}+\a��q�zok����
���;�*��� (��
�z��Oҷ����Y�ߵd��֙�����(��V_!Z�Y�EMe��XJ�`��f)�ބ�n��) �a�כ��lm����h���&k�Y15z�vh�
.c^ �{}C���@чt�lu��	�$ͯ��A����s���s���쳦J�[�_u�r������8�N1�k%��&ά����{��(3;uǩ��V�,���Ԋ��Eb�b�ʄ�qTt�b0��v��"͏���A+x��X�T�grѡ�)/����X0�]GE�� �E!p�(� ��.�v%��ñ���Y]��Et�4-��!/�	f^L�(2�Dɥ���m�*F����?r�ݦ5)��ǠkѦY��0Z'A$��&~j[��3�v�?1J�|�ȗ�>���D���\�t�.�-�Z����~����Ժd���AZ	d�ҁ��P�>�N�R3�>�7�|��kY]Is �CyG����г�0��x ��B~?/�����n���H���������G�5��Bw�\E�XS9�wֈX�a�7>혝���.u�V�s��!8c�|�);��arև�:n�'	P9�i�RC�����SiI�
E��풉����O�������������x���N[Z�	]��3W�]���V)�����XI�xrq�v"�W-�����Ņ�v��0G�s3LS�/���p��~_�L��0g�2���˃�(���L>C��ykǣ��R�?*��<�MŢ�&��=��TS�E1�XV�suD��(�0}�n��Ey�6��V���P~�Y�N���O��ǈ�r]m_�譤܍�cBnr��aN����n��؇�YGZ���ɺ��O~<[��ϲ�4���u�"��s�������*%g*K���IS��
!2��<�]5p�d�"��c��F.k��&��16�c����j�����g����5�㬉�x䒝��e�|c�|�i$e#P$��L�Zd�
�5��q�ՆΈH����NAc�=�����Jol�h�|s��}�2�Q�#B��!�=���*��#w�����^[��I*����A��9O�*�<u�6a�!�<��U=AJ�_�5�)5)E��L�R���L���z�����݃�.��{?B�
���_�%k��-80<]��Asj :!�k�Kf��FA����tK7�p�&��� ����LX�ww�2�R�Gb��6Q�,v�����A�7��H%W����)��P�5�sju:��i�&��5���ަΔ�,��&�ᘗ_gP�?>3gJ�t-�+��":$���;�7."���z޿��ڥ�U���[<��%���, 
D9s�X!��ݦ_#`@���3�?V��v���̓�y�j�<l|��^��>�h�L�jU���+�6q�⏧y�*�bF)\��bĳ��FI���R�����}$_��{.�����6ג�o�k�����)S�Z�
fr`��nZ��ͅ�y	J�6�����,�e��'�Ƕ+�P�k�KE!��Z�O_3j���t6�/OUgE�c��Uy��v�D�֫Pa�0��No�q?F���a����I�:��Gf�IR�0���y�_���5\e�N{��!!����s%��n��Ї{G	1|�h��'p�7�� R��tE���#�<��LISF��Oj���Ȫ��b���qO鮤��zX�"|��LFq"}$MS�Ύ��M'k2��xuӓ�`aH����#��}q��}�|��{�2h�ce�R���9c�]�ܶ��{�3@�����-x�Kc��(�z�1 *��r�V"3�)	���U�b��ƝX�֑���m��ԡ��*_/�t/O����y4}YB+'�ؙ�h�b����G����n�쾅�$��l��"��}���@�c�N�K�䕆��_o��w7�������;}ZN�w�<I��I�#iE�(0c���L�.����9�X䰱��}H�D�z��8��S����� ��`e4�Bӑ�J`�y`R&��G�o�1��F���	�I�$�`�o	iF�?1{��~{jv�bl�I�3�������v�����_B8�Y�N�.=B(=X�WUa�&>�A2y��5�����ҝ��8%�#���� b(���k�.d�H�z�j<Q�̻	���V�����8Y�
�{y|���d�:r3|4���+E�؟���������9����h�j'��
ߨ�Y�6^�\ʿ^{7b>.mCJ O�ֈ������m��J�ho�ܹ���#Rߧu'[��d��{/��~�B}�%�+�d�d�/�-��w���}a�5%�V�=<�y��B��knJ8�,R�.G�������b �� o��!.�蓙�#���Ǚ����묌�N�
���Q���,���}����]���s�G���h�����߉$���d��Br��ea��.3.�`�𩡽��K2�$���C@T�o#6���1%!!{�^�D�4�j��~Ƶ���������w��Oo���ΐ����J�b��� �����Sn��\�=����E��e���J�~�׿?�ז�~���]W�U�4m�}r��}�E�&��M��،��\�� m�ӊ�e��xGݿ�=���b,3����,TR���C{
"ه�P�%O�mq�boe�Om�B�S��\�DѤ^ao!�~�j�f� >����֨�٥�6bE��{T��I_�����?;��Q�ݗ>/�����B0N�o� ;��$��Xr	��m�qL�?>z�Y�7|�b�ua��8j���� e�8�ʊݤe�G(^��жTz�
E�|�-bl��_�^�8R֨�ݝB���j����y���FwL�V����aiަ��QP�=���<�F��$c͋���%���bV�?Z�X�ٌ_VI�ר�gq&ob�����/���P�Q����*d��Ƀ�1l�-����5��QO���L����{n���12��@*rn�f��'}�dQ�s«L�I�F�ZYdvho�����1}���&�V���(ñN��/��_��(�Dz]
`lqs��y�������[�X�tKq_E�{Q3Re��v�P�/,`҅�R_Ѽn�MԒ����@I�+�g1���9Ub"6P�e�n���_'��1س9�C���[5�v��[��Z�2�v���T�~��ܗc��]X��&6��*)s��4L��]�>92u�J��9�h`��hD3�;�Ǖs����>&aQ�w��d��o��t��d�檊0�|�ZV�(o�)s)��I��Q(X�^��b��uϫh�� C1�v/�w����Ć�.U'{vbu��[6������Og�e>�e̒U����a	sB��@�ۙN�� U1[�(�n.}��v����*��3?.:O���ہEna���T���gA5���놬e����ё���_`�E��A�"9pBN�{��G^�;���[��v9s�]�g��aQ$m'���\ou-��Ć��N�q!��okKஙe�;���@��z�?�.J�E��v�a`���;�~@n9K�g|�Z1��(��k8����ˆ��4��K�3\�"	���?i���)��w��M����q��g��nk~���q�g�9zR��?�D�q�����t_2���L?��Hs#�R�I�[�
 ���1�`�$!/l�Ueh(1;w@�E�IGzY�P!u�-��T�����#�W��q�����R"������;��^ �(����=�H���&�K�.��ltsP��޼&��H#\ͯ��ہ�D�$�ͦ�9�8_�}������ˁ�f�|1NW}U`4�B��0��<kA�}�=!|I+ޮ�>z7�_��"��ޭ���8��u���X��eƸ�6�����kT����O�ܤtkҰ�86r�	G�.8��G�wa���Œ�)�o�����u���Z���s����L��;+����ҡ��G��L,�Y���T�\����loq��ZR�J���h�*����~�r�V���W�:�>j����x�}ԗ�X+,�1����Щ�n8d:f�l6$(��%eu�xq�utD�<���ը:߁�L`ؾ֏��Y�MǮ޴����^����M�i�*G�o�"����h	�%,��dC�F�YD�M��:N�uT��)��8x��>�8`��Sc�?h�PY�������{@��AJ��_��(�X�)�\���h��;��0��1FѾ��8%l��-��{5��r��Q��=Ǐ+aCo�Tާ!t��U�[�'.Y,����[�O8/����&
;cܨ1 8]�/a�������&@�GP��gL3ʌ�i�$5�T ��P��Ѣ%�g�T���O�O�HKG��M�_�SS � $�4�s+)�!�gGo��E���,ϩ���I����݌�x��H��\V��&�>�q�@.Tj�����`��s/>+�5����ϰMa�_(L�r���.�/����e���5�9k8NW!�y�d|.pi����s��LEL壟���ϙ��s���&�/E�.�
4�r�.1+Tב��_h>.v�h��mgM�r�v�J�~�f�HOY�F��?��P���G��'���&ꞯ��Q�b���g0!���#�LGo�^B��%�\}�|#tV��+�ւ�s&��v�W�+�0�E5,� �x���Bg>�b�i��v��K�Pb��QS�I H{�CT��nbX/���K�8)[ ��6>"H�0Q���Y"{9�XcL�I� ��������?��+Zh߄�4�o� c�3�=ſE^a��CSb�q�Y=Ir'��"�<�{A�)�G�y�.�8#_�a��P66��s���\c`<��q@���-�9D������s)FV&R8�/�6�z�
N��2��3�~��G����l�"�AD�O/dP�bR�wK<��fTW��a�Hc�F	U]�[}�!OC�0���4���EP����9��~w���^���S�۹����w@q�����kNq!&���� �]���y~EB���D��-Ƀ1e��/I�{���� _�:ַ]�60��%ha�K�d���s�����Y�6��*{�w��U^_4ɦ8�"ˤ�*H3�%����OpKm�)'>�Ե��Z���bBLzwd�v8�P��pXM^#s�?�n/v�}�R�g����U*���OY'/)���yE��(�~�-�m� ��3'���|�m���eg1W�7MX9��ԠC���Y��h���wu�X&�L���jP��n��=��2��ěn�[;D�(���T��		~�Vrz	��E��`g���v�+� [cͩ��a|C�b�N!��[)�#wD���|[T"�^	�%&���o'�!�S�GM���ȸ�.��;��� f;r�@?:�_% k��{�����7�5(�$�����(�F�6��ey���ڷ�ۊ�Һ�'<�D�|���Lo-��MY�E����(|Лh�}����:����e/9e#y���uk�;�3��Ԍ"dT�羀 {��a; ��Pl=���̥�e�s�/�X����%7�32���Iޯ*xG����b�����t����(�h��;�	�͡WD�{~Z��<��8�Q�� ��>-��?��FI�&iw�w|2�Lll�$��r�g��6��1�Cc:���������jE�����Po�J�^��u��� yD\m@��5�2�g�ρ�m�G��R�"92�:}�)ʼߔ�9?��F�u��&1���w����Q�(M�l�'���� ;�xU�Ƭ"HEB&��G]*_�鸃�^�ª��jr�2;r��&��m�|u/qL��OT���;l;���,�Y�W�
3���'���n�Z�ff�	�TZ�7�e�{�[�<zHB�	����9�\\�ށ}O��U�Yf1�z�p�v߿� O��xa�~-�CR��9Ԙ�g�(�����DR��F�==�� <͎u�H��mRj�� ���P��x02S�KW;�j��?4�!H�7(̿����8�'N� A/@�/�SmQ6S� 3_NsֽV��yg{��˭�<�~���O��F�}i�V�����:@N�1��{�gf�L�� b��,,ee� �- \xϯ�:���ת5m������A4�B;�Eƿ:A���a#v���!<1��Ϊ�H69R\�ߗ:C3��;�#�8+�̗����æ��tPe.ct�q~����F�kJ�w��^�x�(DF	4+��X�_˼T���dd��\���I���拗%޿m����aG/�{N`H�s��b��XD�%���Ż 6�M��sЄy�o��E&c����ṳ�t?2��^�����[�ʘ4w��W�s�&y ��0�������Q�Z��y��|���*yR$~��02������P�n����^E-2�S�Ye_�Ҳ���;ْa[8�b1@���4����_�4�S�t�!�����*'�q ���pW)h�Lc���/H�a�y1��fk�	��8#��)|+P��ԪW͋�"���.�$dE�����lG��C�s!R��|��� #r.!��Z��q"�����s1ݰ��M��zf��tӛY��M�C{/�!���o�h$�k���Y��S���ݎ�� Y�fE�����
��wڳ��%�^�0��eQ������[*L�D2�p��U1k����9(��&�����d+?iS�zV���s��{6's'W�~��d������|�]���I�T�����	p��j V\��;�|�6���6��ƨ�@�@FrSy��9��]A�W��|���"vi�LvokI%�
��遤�wb ������w�>��PED�B'{TQ�ʶ�$����D ���6]�e��6y)͊gmB�l�u��Dו�>cO%d��{�r ]�"V�H+X�n����N�z������'
EV��
\���?�ʡ+�>�MEw����D���i槮��Ak�.k@ϸR	R��!ÇP�L��2?��_m� ���^�5�`J�$/��_ޮ�.�N�i�VY?՘Ø!�Vt�����J\��mv]� w�ad�H씶�'b;2�#Ĩr@@>&Y�&��ԿK���6-	=�to�o��]l�ܜ����n�&��sϒv}+,^�f�q�<�sg���	��k3�c�@O��Ws"H�?TR[@�Hq����_Z�^���{ ��c'qsѕ@$L�{7�ZA�x	�P�]�y����^�y�L�CNI�m��	�R�geu��xt�.V�s�WSX5����y$���W�?G&~?DY����*ײ*�|��ۤ}������ҕx��JXm&}�$T`|�4��1Y�h��v�(�� u>!i���I���A�_<G�G��R�Kmt��¨sN����1������;��OSt���@J�¿\%Yi�<�D:�#/�G�(�jA
�'(���:�;m��'��;��s1��kE���Zf?���tKK��s���aQAY��e��
ⷳ����
rk)�C+ {�`P˷��?h֔����r������@!P��DsZy x=(Frv�������������]�n��2+��>C��A������1��3W��X�"	[)_P3a�ͩc���7>t��m�ۚ�Y�@�9����S�fM���$���r�����+
4Y
	�����J�[�,���b��.[�sB>�Zia�0����12�G��ƴp���(���Ic]��9���/�Lغ�$�|z��E��Q�춒�Q&p�4�(o[X�Im���x�v=V)E�
��u��w�v�P�C�y������	�Ԥ���x�/*�Y��s-R���Ո��ϙ������y�{O��Xz����ʼ�2K?�u3�B��L��݋�+�>���("�?i
	Mө��[q��������@7�&]���0p�����(���7�qf�^���3N�:0��4,Ji7�
J�kFq�>�'T�:��'�tK���3~X .��߃�G��W#eҷ)	�WDX�i�����i�ѕf�i\5�q�4�c�6�XG�aq�C��G��Ļc�Pc�B��,9�����0��҂*�m�}2�?�7�#[<�2<��a�A�2f�8���K3
X{���xq:X���ח�(�h\M��$���|�;>�%SL��ږXa߁��b�!��:��ޮ�;��Z��⇖)єc�{�Z�Ҡ�B����]J��+f6wX��ZY��q<��=biٛ�5dF�A9\gBsu�8oTS�3�y���~rk+ܒ��)>��[�f�x��u:2�6l�a�q�ڈY��l�'��P��?��X-��
yX�HFpq�o�V��}��a4ZV�vԒ�����J���'�x$c��)M�����0���a�u�-�.?�S5+�O.6/`�0�X]>g��]ᑤ�� �L�j�H[Y���q���3���%�O�>㦯�{�d
D7�w�;b}��pwz�ns;��� �8,��&�;��P��W%�H2?L\h�9j��Ṭ�31����a��M�]�R�絶�tlWw�bj�iZ!�� $����o�o�����^�YP��(�Δ� �%����93�D���Щ\~�Wku=��޺GG���6jϱ$9pv���	¹�N>{[^�
OV�G��NZ����|�:֢l<�Q��#�D~�?�4-̀��s��K��z)�u�B)���*R����;,ե�e����� ���m����C���n�u�z"���Q�H?¿r�~�o�K�~��Y�qeG�V|�r ��G�t�0I� ���N�Ƣ�$RM]��,+�3%q�+E���<&�}��tm���b��j�w��D���N����V�wW�j�%�č�+g�._ˀ��W���p���P�ޅ�5?��v���#Im}���Ѱ#,ctQA:n:f-2� jtU���3un����$�
�*��H7���Y�[)z��;W�؀i��:�]];�tap*��X���+��	���v��t�?�ݠ"9���0��e�4��|t<^��R_w�2���9�ᐕafU�����s�*eq;����o�QD�����ט�f$H�U���j�C�^�'xJ�kF�f�,����9wJ�M!ܓS��钿c��"d�a��Uh��4�%��lmN��F�%N��q	� C��5�w�=5b���$/�C�����UZuɵ��[���a#zFג�N\��ض,�i4j�h��Ũ��5�ゕ��V�����^NXE_��pi��'=` ��Kr����תG]ƨ �G��k=2�!L�%��l)��+vmBv����~~���� U*v8�O&�A��lZ����$�3n��H6^;���U�k.�AӘ��yN�"�G8^�3�Cwђ_�ai�6-UՍ�N�����wm㍔Ɂ������+='�eߔ�$��	8��*���'nl�g]�|�G�꼈 ��J�d�٧�:�zL����;�Ov	�.k��G��G�N6��҉�.G��`�`���3����8'r�]�ȠC�^�6<s�"9�C�pym�������.)�(��*߼��ÿo?/4ꆢSB=;�p���w�	�3 |ܦ���9��c�~['��/m�K7'w�ң�|��#����W�����݅���)*�F2ƀXx�dl�d'	�2���M�$��ғQ�૴�<���:�8�,��N���ʴ�/�+���e]*b�}���2�Q.t�1"�/>!-]��d�{�A���Dp29�jY��74$�������[��?��^�`�x���'�Q���t��Q��!(V���q�ԥe�����Ԉ4�IaT�Q����ɶ��<c�|���{�A?R֨�����% ��mƤ֛�D��w���^)�T����b�Xz�K�q�-��@p���[�����r���
�JZ�����JCӵOC�z�L�w�$:�f�����i�����ծb�Q��V�)2X����3�QN��=��[=���!�9$H��|��ڧ��5*�^���4�"�MU�c��L�{Q��tk�+t��W�~����ŀ5E:�ssY����_���a�Nj�oa4�Y:Pi2��D���������(/,��oo�J�HPe�&.�����YC=Z%׼S]�ů��M���ʖHo��,�&ǩL�.�ʂÆ�=��v�
3.ښ�C0�zյ�����$嘻���-#NB�Hs �z�ާTk�o�B���q�=��: NbxmIx�tt������xW���)jM�-�6����h�he���5�4���f'��I���2�\��4D�l���*���X��r��d��z11��=��޽�I�V�{(qA�����`�6��"~?C���P�:yc~�m��m�e�VY����#�K���V®A�P���C��rˮ�Ö����������$y�����bZ�9�$,�)�␠F��:�Z�?����b|U�6� Uq"��Ć�cF���c�i��wS����*���6k_SP��+��!ܴr��v
�!^#o�SE�0s������-3}!H舵�1�^�!o�zb����
�&��iD�9�~�ywO�����ƳF���_B��t#ڡ���SPq�(�E�{�Q��B(]�B4I�rl���3F��1��T�����Z�� �A�tK��ph�A��X��!X���5��[�|T�I�U�vZ�@��{ʡvp�}r�w���XpR���AMQM)DN%��!�F�5R�9#Gu̚�[�����/ךP�x�$�s�{��e��hk �W��Ԗ��__2R����=��yuT,�b��2E�]��/-�'ߛ9sV��j/}��S��Z���X=�qI�P�Lؗ`�5t;Q� ��R�m;������J�v�P�aƲ>M���c1 ���~y��=[�#ۆ�4��͐!"uP#�aRK3�W��6��O�
T�%�ل��t$Tm��>BVD�^a��Q�*DR ������T��IK����T�N��.^��P�Xpʴ��_�����m�p7z�u�?�H�+����f�N��+��3IVG��~]r�;��T&/5�X	<3��[�o���Ͱ'���p�.�4f�v��_^FY(+g�M�FM���6dY�O���Znڪ*�������\��PnJ6�����U��.����@���/M��a#kG4��'6��"�2[�A������-���\i�ӊR�@Іm��6����'�ݧ�3�2
T+}�-��V"?.������n�]`$���`��C�joYJ/�r���:q��#�0�9��U�Gǝ���ɡ�ko'�䧳� k0A!��B�0��uO|��<�ΠjF?�����: ��c��Z����ܚ; �)�ѵ�+��q�O�<��Y=6������QXA/���9EE�Έ�(��]X&���ҹ�)���oWm&a�o3�3%DǮ�e!�CXcm�j�����CH�?L��\�͊	�G�J>�WJ$���!�j|:�!޻���肗v/,}L�Br:�c�\
(<Qw
$ �c��
�Z���z'��|���s\���,E1�Ͷ�Y�*�(=�\��']؛�[g�K�3<��ۃ{L��?+��K�G.�X�nt����ܪ]�W;x��Ŧ��h�3@0*��K��o�1�����p��$��x�h�^�;��! ?�|k��,��LgR>������P��:T���
���/:����+���2��Zw&�Ė��x�Ny�Ռ�ԯ��%]��m(���G�)k���Ό�B8�&�:r� �U����+	�!��x=�R��TQ"��+7gJ۟��u7�Ta %��U�͍���QP���#�v@��O�?���]����zd%95��>�4�nw�G���0�.~�����Nލ2��I�uP�l8��IO� v�E�Z�����Q�Mv\���ѩ~<��#���_�6|ޣR����vK�H1a�ОyTk��953p&��|$(�����N�݅�2����^�b��*�]sQk
����	���#w��1�����2�Q� [:�~d�q�hh���ur�,��X�@�=Q��꾔ڋ�N)G�i�7A-h����i��.ʁ#'J��'�ي�����3;�.E{�-֝�@�7Ę�r��� �=:�����O�"�o�h�i��<<t���ǀ%o���W�ٌ�$+��kr�����N�����b��X�j�U'+�|��{o��r�3'�z	��qCկs*����M�9�*�>�!jw��9K[���4�V���c�����H��q|[ �zy�av�R��ȝ{�%sL�/.��hi��^����C�(�� ���x����r�sB�C���3�YhP8��j�C��޴ �sdP��h"?D]lXܵʹ���qHnBޕ����F2���D����۱q�N�Q-M8���A=;�|��Jw�Nh
j��\��t�I�Mɖ^S�}�0��0�#���t?�9k�]�n����vGޥ��!��7 �4�R����҃��*��&:�Q��w��3G�u؂�,�8p�c�L�	�y��23��F5��"���)�r-5I*�UE��(tzʪ����a������'w���lK1����a)	��q�i�
�y��:8ؽ����i�{��������MV�{xRM��g��)�)�(*�
��,Y���u�;o��F�^�B$������qΎ�I1S��v�����F���A��>�x+B�q)� �2���槪�_G�7���wi�����Ii���tPm�a}���g�N�	?/K� }/.�?��sL����#������v�EXf�w��X��1R�ѿ������$,a0+�m��͗����7�"3����=\K3F�����z'w�R�ԾQ�]�1��7�e�N!>���l�o��~���T�����r��SVx0�='r�w�Cp��#�Ϝ܈�5*�ˣ�&�_�L&����c^W
>t�%/��ɸ��;�o���T�`h��K���TĆ��x8���/"�Mq��2�a�c�
��$�_uV!z��L{gl]6{U���6��a��Yi�3�d\SZE�H��~��aMn��P��8��f�`Kae�����\�&KR�}rO�B�W�*���6}� }&�/�Ӣ%��:�@sb4�J��ɯqx:�3�W3t����B(�3r۬1����3����Ov�^�%�xR�p�A>	���+��C�DcNbkS��ߛ�O�
�����&d��|Ҁ,t".���jj�h���ۉm��i������F�N֍�_L�$��QU���j0�,xX��0��302��K�aj�7�^O*�Z:3�䆈���)E�[s�����28�-6�)�oY��4�B�1mLͿ��rĺ.?���*)�7�%���{��!�0C�ϛRh�����s�����=>���g⵴Ik�����D�຅`;�&����z�q�~M�/�z��:+Fi�R�z��q��Y��BVP�-�E��8��B�}�-�ݍzUw��/�.�l�_���Rқ��`hy����~���q"eX��1N1^�kE�G7:��b��\�)�tL~���'p�V��~q��L��~qsT�$�ɥ��1�5c�x1�F��چ
=��*J~qx{|�8b�y!�~{���yFE��ZR�Jz����]�9��~�ť#�LM�������e�$�����eDc*�ʹr��x?�[+��e�X� ��:�]N����>�`���\�������I"#����8S��!x90��Ĉ\���5}���x��Џe��u�OR/�l\�_��yCLצf�ٺx��_R`�셲��yp��-	���Ԙo��C�$X�����ܓ$y�DI�\�kbQ�R��'���*��:�5��f-�{�S �~L�E��͈a>��w�`�*�v���j��@6��~×I�j��j�(s"UI�Q�aO���jQ��!�&�Q��A�3c �t���jp�o��~1`>?.������g�2L�y�hg�F�@
��u�!Ҫ�%\��5��	��	U���'���e��O���\��;�����ntq�jg�m��h^� =�o����Yo�nD5VT��b)����:cH�d�P���e!�5��^\�P��S芏�!_O�ڹkY����	ibz-@Xr�� ^�k�t��"�O|���D'�苋�fB��?A����D6v.��`5qj#G�I6�ޫ��W�v�0��#�q�]�ޢ�&UQ��v�SE���a��&��*+����k�=���^%w�u|سg�t<+I����ee�3S� Twlx��C߃�`2�"&�.4D8p^��xAW���3m����n+k���s���D<����� /h�J�	9��V_��7�B�)�z���2*���)כ��$�ސ�ܴD���kVP���mC��ȟ��4�q����~�L�?.�ȏ跋�A�����k���Ԯ��>P"��m�m[bPc�3��tNتA���:�`������o����=1�?����!!)�p�,��XP��L�!bV�$�@����d�wkQ���̥���2��.3_53��'?3l�pc� �`8uC*�� @t�y3E�׫
Г�֊�����8pБj.v�CH�V�Ql6sv��N��p]%{+�rj�?{/a]�����!��NW�Cf�KJ%/���9KG'��㛻-2=��i�#4fQ�b���Ó�]�Tq��|���Ⓚ�[c��u��}M�;�:ɋ�~����Xk�u���*�mrY慆~�����^ytl�ݢ�!�Wc���&�R$a��[9B=|J�y �+�'w?���w��
X�i̖��U����*�G���|��hq-�K	��uN	��q_(�=�$G�E��s9��D
!魈'w��Bع�����S�Ŷ��O����MԧYtm��.*t�N#�U�H��k�v�N>���qX cnJMJ�B�X3�j�t �gVP��K����ղD�w{��1�!���^6�81*�/�xV�r������R��Zmz���a�p�JI�������oil�� �Z�J��6���!�ԝ.S�)|?TAK]"XK�:��E	.�FP��J��hN�g���,�m��+��O�Ґ�+e�9���W#d��=�'*ϴ�ݢ)6����E����昊^+�L-�ESL�O�r�*G���[j�m�((�g���MV3�A���Y��Ǯ�������짔q2�bt��e9�l�`�ȿﶏx4O���[��c$�X\ⴼs�ȭ�������ɛ�p�����.!K��l�d�*�#��n�qP.�1�J}q4�D������}v2��G�u2d�����72y�-�j�^��n���k���iB^
. �k}��a��Fܖ��`�Nzc�{%����S�ɞ�D��G/�(F�H��r����VCG����'ӈ;����X���	M�h���>�6b��8�<��&t�,���^�����$b	=C�W���}yH���2��܄bm�|Q/��K|�[-��Z=�/���ǉ!�7�E�R��နq��5
��"8HZ����1����!��6�����/ I�ٰV����O�케x����k�j!Tn�X%
�M1����H`�������y1�u�oz�`��5�͋M��h[�x�a�f�ؚ`�x�����}#� �5�l��D�2��/���T�fҔ�e�:�&���#���M���gMӃD����x��@e$���m4�e��:Zz�mP�x}�hum�������Z��&�'��v��W��#t$�7�tV�	�V������R�<U��a�pV�����U�lH�NR N�����l�k#�T
�<A����=âKOO�N�����3	G3���i�/Dbj�A]�ȵ�G�bJ��b�!��w�Ӑݿ�]��*�_�*e�1)�ܔ�Ib1�P1�/����	���<=��$��p��s�H.[�R�c�mc?���*���$��%?�I��7A���7]�)A�d`�z2���|o~8΂�����	�%X�� 9������%]\�6��޶u��(-��)��7�=H�k��-9��Bɤ)�Śp�����%�	��X��(YՔۃr�l<��|�v����_�%7�w�`�c���Ƌ7^����t�_d��	�9�p WT�"��c�����.#K����/���	�:j���Y��� ��$�^n�4��w�9XT�w�
�[��a�/<>�!� ��i�Z�E}��z4�ջ�u]�Ŀ-.�Vn�����*RMpZ��X]�v���$�^�F��n١��?����)�����A������j嵐Ŷ��9�Ȟ���ZrUeG��^�NN���҈���=,��ɸ��y�Ո �*XX��a���P��P�����؋B��F��Di��,�����,�E�8Dgri��6��|���$�Mі���,'K����e9��Tp��?>:s�P���bg:������(���6���[*���T��{%�RI��ԍ �
9�38]TH�y�S&{�"�Ê�W��ǫ;F��S�VUZ_эa5Z��Y`$�$�f�dO�)��m�'���(�=7ɪ(9Z�/}j�����g@���g�I�6��E���i��S|�l�� ��kޣϕ��?�@��8�G��ȼyD­��\mj�W�X�m�A{�Y�i��R�]��1+��S�z޺�8|�KZ�W\�e�C�`3��B��;sn�A��.�mp�<d(�{������4EB��*�S	�eF��&�(h���'C`�'��N�����O!hR_�4�5Z��w$�5�^[P�m��΄�����c�.R������+�o�����_\��iDDD��%��7{��28tdY�?�Z���C�X�������/"�	蕕���U��p�֊�Q��3�#�R��=�A���O���0��S�P>�2b��<fJ�5�Q�	�lQ��emq�C�b��پ�ꚡ��ծ���1!��{O���<Ȧ�������_ܾ�FZ>N�Ǚ�$C��j�X��m�	�lO��Y'��H!::j40�߾���"6�cυn��;8��#�cr'xb��F�"�v��/u�4��3>K���;��R���]rtKS�g��!��Z4��Z�k;$m7�nͨ������>&�t��ݶ!��\��(ȸD�1�m��Z�\����)}3�A���b}0�Qs+�E^+Vֳ����>��!��h�c�+���MZ�O/���Z����7��sV�H�6r�0��RI%�O0Ǳ_��=5=�K��b��w�IY�/��r���E���X�����y�;*C܏�4�Pl��!���t{�2Eo;�Y4��W%����$L���n�丆���[�>���L	7�s3��U)�ī0���v�����:�vϽ���u{���aσ���9��7.p�Ս5 ���=�"ٍ+�N�p�*�E�g�*;����wGa=�a4>�D�UB��e�7�.�p�x�>�d'Y��EL±�����ws�e"�٠O��X�)F"2�o����$o�?�;@��3��Yd)�t��_A���i;���R�u��S؄!�`��T�N�wl��REh_c�,�9�t3b�Ԏ���n�U��
5� w_	KaD���{A���ا��N��Н}�|���M��#�V��IӾ˓�'Л�����6/��w��K3��W����& 	��/ۗ��V���ږЛ1�M�K~J�C�C�	�g�2#5�:�ƎfJ�n}B�4	���"�k.���L�њڻ�C��W1����<�� f�C!�r��u8?��LT�����J���)�!���oUh�����@1۷˞ʦ	7�L�������:.���B�+�/�\.�zS�6m9��x@/c�]��<£jF�ϺȲs*�X,�v�rgb'�:�L��C�+|��mԸqO��4x!,y���H8�B-�)K�eX�:1b��v�Dw S<�M�qja_�æ	�K����ɑ��?Q���6
ԴK�n��@D��o�zfy'�1���hT�EuY��Y�&#���UI�]?����.����h%���ĕ��|����Ly�z
֑N����O8�",�2\�:H��ݯޫ#���&H�+����)]�U�K��6��u�k<��S���빋�h��&��}>�@�߅�l�����ýxY�h�MN��2���H��?���m���ߥכ	���ik�����T��ϋq�;����O����hG�[��
��N�3
�������Îr����ׄ����J��B8����M�ρ;xq
ܝ�jB���a�}?[PR�2.������-c���"�܎5�X:[(k���"�Z��v4?GS�ϧ;�
ۥ�pyH��'䠸tg�����[_O��摲�)I%�> �����<���:����Ͼ4�P�p�iE�F֭�,�=��w�7��D�w��͇���(C ѵ��4�L�F"���b٣뭠ͫ����u���hפC{J#�Ҏ�@j;�z�t�fx�K�	�o����Y�ɉ0E��.�ڇ"6���Dgl�gܠL�g^"i9c_�	�(�V�y�vok.��ژ�<�z˻�T�Ð]�@�fG烇'Ƭ+�+�ǈ��?���&VE&�{�Lľ�	G��n��KA'D��R���aXlAl��^ݽ�9N���'>��MȾ|_=,����$5�>-�^�p��ވ����$},�� z���)��=(8�Ď��Nyl��S&��
L�| L���伳_dZ�5Y��H�5S�o&��¾���<��|����ǐo�[�ƠE
x �q����7R�t����rU�����W��xP�%��D�8�嬥B�&Q"��Ԙ���P	��Yc�U��l6|��3�W{qbQܟ���Cz�G鮬�!�j�G����H(�[&%�VQu̪�����N	V����X6=�@�}G�E��skRb�b�pBYg/�L��a{�²�n6`���� ���?�s����(~��BuޗC�@|v�i�o "��<��j��^T<9ި�҂Ԅ>�ܜ"��d��rB}�D�<�w���ۡ��R���)rQ�dw����/[L��
֊��"it�dr��=��k������pLk]����'[�3�PK�R+B)jZ���f�obJ���ƌ��f ��B�3�U�9v$]Vw�㞞o9f���9^#���~�1JO#@ Iv����ܑ�5��Ld�R���S���E��Q�ۣ�5�"dX>�T�k���[N},ovͮ���b�~��A�su�3ڹ�ʵ>1)؏�O3�(�Y���}C� ��b�ū��u;�.	�Y���_aI�#>.b�?��v*�x�A�%�� ��x���^�x��3�� L⠓��C�A��۩��~6�;h;?e;���j~[T;+C���&�g��M+%*
�����p��_+�M�����d�H�໶G.WI�K�g�OՑf�o��(�g߉�`z�L��3�y�0����zZ�V�Gg&�º��.E��y���<�K�Yg`�� ��\�ņ\r���Ɍ9�,L�с��W�#�p>���b[�06ܽj�������2�r��8�l<4m��(�o�2����h�E:t���]�-����-�ܾ��ۡbǰT������ƍ��_��{��Ð���!ʺx�����}V_�K�H� ��\�_T�����#����9�ƪ��5(RHd�~d�r�G85j��^+�����Zq^��/R�zv׊4rqU�(���LZ��u����ڹ-5ÿ��k|���u�����w� q�o�uA~�pL�\��*'Kڵ�v�ʗ=Wз�i�"*�ڎ��ϙ���x�	 t~ܰ�t�<��� ��H|��� ��_��$�5�D�[��K��A@o!y/��̀���?+�[>��{8�ԧ�~�w�䜞��8G��`9a���$�4l��J�)��4@l�>P!�K�G�?���ҏ�ⳅ���7�XW��5���8�=z��y��)����0�2h>��V�K8ৼP��zfq�ǥ�,V����xk}([�~���N!��n����a`���剤����qI��46S}�x�j��[2'�|�7�c�}� 6�O�4<d�����1���j���ՠ1��9��߅TvB��d\���x��<;������O´�x�\����g~/��f Ek������ӖH�g̓0�"�%�� G7��tZ����_d����)�2=�[o�!M�?�h��	��R��u�~���l��p&��RT�*�h��0ڬ?���9���)�~�C&
���D�tEt�>x��Z�3�5����\��C%+K�K�j�<������"��U�s��ᅤ2�)֤��� �d��������ڿD���̗���bڤ,w6L{�;�O��a����#vB1'��	�J,�O������ѩ�6k�~ԏ�TΥ5gȴϠ�0߶�Ͻ�M2T^�u��M����[�	ê��}C�%C��t�HYאּV��)�L�J�b
�UZ�XQQf�YP}��FUvtf�b�%M�篴{��
+���ԉ�ɓ�E�i�������6t�z����ɍfz��0f��7���vROY-XX��J�1���Í���{|`��W�	�'�:d�ϝGΡ�ד�8�k�enNc��/�����(������/o�[��%��a*S�#i�S%X��a�ݹ�J�]x�7g5�/���c~��i��c c6�:��H倘R�;�gT
9.w�7d%����}/�vG��o�|g�M�b5�ƿ�^���n��n���_��;@�N:�i.��f�ɽq8������fi����5�4�W?���+�(�����?	3r~R��X����K��Mz�E�Xdrq��R�p'�Vs��e� 6]�y���oٔ�_���<�Z���]�*���3�4�5�YP�w����Osce���.;(���o9�H��K�
��SL�h�2|�Pv�3%�A�!Lq�A^�͐�(�����NT�k8(���+~���^71q�Ҁ�Ȩ���Z ?l�ɳ���H~"|B�c���K��ύ�LH�B%³���D:�@&����@�a��=i�>c�����E�����*�׏��;*嵐.{��_����#���`ä�S������i�M����נ�a��h�),�cI>�x�K�a�X��l/�#=Ň�]�	,���`�͚��1�s�}gQ����#�L��̽*A=�|;���jT��x��z�Û&7�m��9��.1́tx�T�����݂��>X�%�.��q�J_3z1�`d��F��"��֨�B�ȶ"Q�lWT�i9.�S����M᝾g�"g@4w�4��n�,�ᕱpI��/� w�^�
�K����?r�x����:ݥ�D�Bb��L��׿�����gO��~0������X��<K�	�j�Y�84��]F8ޞ��%ɩI�����t�� )�CO����f��KϦ��[K�\l��L�u�gK]%��\��<cb��M�V�.?uL��Ањ������2K)ЃV�2`Ɵ.W���Sԗ[Z���t�3� �!e���n.J_׀�G�H(�H�?�R��׊�+֘���� c�P(![����R�ԕ,ĝ<=gs�]�kP|6D2nP'������<�2m�50�G_OLM�&Q�%Id}���&�26�ݦ�3u�g�IM/<���Zrg��k�Fsf)�EkQੲ?pl��w�,��+�r-O��o�܍~sRZy�w�=�Z�"k�-�z�̃��Qdg�F�B5�YB��ju= �*���u�0OZ~�Q ��[>�i��'��ѩ+���k5xdѾ��2$���]�R��(�Ǩ��H�{e�M�v��κ�i%��˨޷����=x/U8V�`�g-�IP�j|y���)':�,�Vդ7��5���̭i<Tܰ����H������i�IGm����j���^4�uY�����	6>����BGsOɘ[|��sB��0���� y�����Aӂ@�ǐ<p�at���zK�Q-I�_��
��v�+��9��nn[��v���|qu�����c�&v�C�����\�N�g�(���i}��JT���'���P��B�ia�i5�ҧ{��J3;�2)�BF;	���g?���J[����ᠴ�v�f��Oj�;ƺ�W-���{$�T#������=���P)T>X�17�������e��
�$��EA� �LP#�R����2IU�ɶT��C��C�Q�9������.w���:e@�5N6���:��@� c_�~�}�Ě��c@��*�L��⾬Q^�Ì���r� m��H��Mm�b�����
܈���<e% �<��/�(�Wɹ(�e��ޠ�5���cOrOͦYv��u����=��O������d�
��6I�-KetP��ĝ�"��d�U�y@��Jêi� ~Lks�S�¯}�����r�12u�^X�@�[���d����I2k��,��{T�	��v/K�c�͏���R"	���r��ݳ��J�� �0� ye�=�':����g��]�m�E�?t��E����N&����|;�����4c�QΖ��Eyj��:*q����0أ<�MѺ�*�6k˰���{�@Nj�;��dq�\.2�{O�Ն滚6��T9c��$B~R0S��Zm.��"�m]����̷��	���aI��7���`>�X:C�{�Й5�B*�p��.m��z<�gWgd��d]�y:��u���4i^��}�x&CYHu����-{HJ�ty!�gHl�kgeo		Ng�A�����b�9��Uv����(���*��[�h�H�ѷ����\]��ℓpW,���IN��Cwd�m�A�A�5��o�&^ɦ���>�$���iF�`���N� L�lָr�XT�jSO�4z�aQ��`^z��ا�)���	����ӑ�����賗�$u���b/R���i�g���δ����ҳg_�]`�{�ڃ�?�r����& �p�}��^�otM�s|_�+�5Qͳ�//P�gx��L��C�h��p�eR�dŲ"&*���
���W��I���U��Dm��axOǋc3ѷ`�rJ{��[	�>z#{?C x�ᬂ	�S�>�����*5F߾�j��������j�*v��v���	x���鱕���U}�t� �a��?c�a_dU ڥ|~,���©]5&��GS�ֈqz5���s�a>s�Ns/��G:����o�Cӏdn�kPO��]����?c�\�Gh2��ܷ]��T�BgZ1��Λ���E_�p��j'y��"oK�`
v�6ԫ:s�r��+/JM����}^=���ٛ<QX_�5j<�[�����z�/8����T�8�M6��Hߡ�y��s>]�J� 3^�>�
dy��u�~�-�G��L�^���),���}�4o��t��B�Sy�A�!!�	�1�ᖔo�i ��Xt�?�y�7��f8�,�����54{��'�4 Ul䂊ƕb��W(	�8�V�y(��(b�� 2��\L���҃��������������y
lo|'е���>���_��a@�ܽ����&��j��t��x̸{I�u�EX��.pL<t}G�[����>YC`�1.融U��mTd��{�7�&P�ʊ�/���=�_]Z�~K���PE���j�UɎ1��������l��j�B!~����k4��&N��#��r����uԄ����v"VP��8/�����2<��)
�"9y/-�]��V9�����f����?�&5u�����C�(�<l����V��=�(�z�^���
��5^?��Lr�m}b���d����f�[v8ŚC{��U�Mf�׻Y@�.'حG#�^�i��?��K�Z<���3陥����ߠ��IP��*!`����6ٝ�O���=�<�S^�E�^7����=���N%���F���VyG�GC�y�0����n:(�zR��Ӂ�0f9d7*8�/�= t�K#Rƥ�:���L8I���w�/;3ɉm��s���?�6{�y�9�����c�p8�}|qV7=J��e^��w���äH���W�v���$�$ =����]�F�݂o�@{k�{��K&��ϸ�g��o;����o<E<��[�*<v^�_�Ǝ/�İ!�f]��P+x�Qfɳ�Ρ�p���C�� 64��ʾ��Y��ds��&�\)Vm&,��gUT,�kB@��y��O��c+� ��e��t}m?���QwH��6RN�A��ڮ��(A�+��i'&J���q(|������t���ɐ��  �O�KB��p���}*3�9Q�=�VOܣ�`S�����1۹���π��!Y��'D�-Sf��)@��ͭ0���7�^n3�����ZU��{.���ʁJ��������͡K�$m����V�9�+b�}���ݓ��۵1�
W�b�L�k��# �<]n��
Jld�7�� 2�^�@����eD[�Q4���(U��Cz���е���#<��H�>��r�[�V�HI.���v�R	|����M���!�2Q1��⃨�_X0�7F�BX���۹�ف�����_��(���0`�*����K����D�&;s�^���(��}v�OJhD��p���Qը�
L�U�de�G�ˇr�^^�m�O&�P!tg9d/󧡖����'��U�+�Ȑ?���!OO���DT|pz7X���2u�6!TL ��˄�?�t�ީ�p1�l�-�X�Rhe��۲L�����M�������� ��Y���[��fx�Hv>���4�-��H��I�eN��P� m~�֊ǵgyts�Jm��;���p��<�I���j��i�I~!tqh��ʹ����~�f��^��r�]���g ��隈��Ǝ��Xi�p�	9!�3b��X�ٍ�N1I�t�~͡��8^V7W��ej迈��1�O&
��mBX� ��Ȟ,�#{n K����Bo��V��޸�˷f�;��:A'�s�em�0�1k`��)������k`���<13���!�2š"GsX�����Ĝ�ht'���V�q�f_d3f�p|X� �X<رf��,F��l�H���;]�uP��?�cw���PF�E��J���gV�����s���<�Ӿ�{%�/��dH�7��5B��ʬ@X� ��%�;���_�C0Q��ބg�;�(�-5�p��a�eA�e�v�� �F!)f�a]D��E>�Y (3�5.'h,���$�v��Rzk4�h�J{����°oڠ�^���ݝ�c�H�>o]f˞~�	OL�����l�/oQ��W��U�e��f9A�X^�n�Af��QT����tJ�C�G�3�h�z��J6�ȑ�<�w#��%2P�B�B��f��C���N�Li[��N��Q�D�$��>�ߺ��0'��[5������`�X������9�e8:�Wd1���XB5�c�4�[��"w�&\r-
ÏM[SF#u�˷�\�Ӳ!�/�^8�:c�a�l�ne�o����Ʒ=�Ώ���E$<�䘻��}R�Z&6y�srו%e(S������Y~lS�~��na���%<��ŋ6 �拖�P�X��v��l�#AGc����<G�hZ 4h�b�a\�l{{'�K���J�*22�)��#��W�N��5� �Z%�ޕ3��k�͓�U-+�s=)c=�djV�Q��t}��雵���ܶZ&Q�r�̅��Q8z��h��Gb�i7#5 ��1�T��P��Y��/p���{��H�
��xz�"�?�96c5�ri`��K)�13�X9�8�!�x����Ѐ�c`7ģ������oR{q£�f���:ʍ�fXx�m��Z�	�p,#e!�9r�5�P��l���o�;g�I�t7����/�R+�>�@��~I�V�Vk©s9��"S����4Ɗ�;m�~`EK� ���<�P��UG�DE?x��j�,�����MSXo��m�B�̑��^x�*M�J�t�i3<��[	1�^{�$�hj���0]�NW	��r�fบ'��#���i�F{RJ�!�4��'�<�������
�D�;��,CC0�}M��� ��L:Q��Z�Ɖ񱞁��p$��}�8b���E_�N��"O��L�K�c����Rŭ��DXJC;3Yp��o��� ��
�v������孑��	KQS���KIX�+�lTl!����#�@ns_�����:��7��z���ʙ.��XL˯6&��-��j=6#���u1qz)q�ұ<uLi�6�vϤCT�b�e��p�= �~ň����g����vx#Q��t��;�t�
)n��I��(-�]�.\�Q��u��ѿb��/����8c9�5��5^�o�������dbɏ?�-�R�v�%2#<pĕJ�<Խ���|rJ�ԳQ|�Dr���m���5�9lG�-4u��+���ֹ��E�.�`������\1��@Li�����?�1���������rB�c "�-|���nB�"�8��״Q�{��C�BD�Aaݷ��O$~>\���θ�tn?��A�]T,�����������"����	"�j��k`g��Ł?o����J���I󻳵�a5\jH��*:,T�?�ÿDC#Rhc_2K����C=������G�C�L��J4��Vb<&{�\���{�N�_o�MV�^>�X@�E�i8)�9��HWցI��B�N�n�g�P�y�|���;��&7�)8��r��R�z�+ċ\cε��%Q�tIy搮�G��y����T4�9�Zj�4aX9�̓�Vb���=2�;E�S��$5����k�h2`�d�z21���"�	�u�<��H$�J�����)��l��(���õ0�_.8{����77��tu�J`������+O��"0�]SbJR4������1]ǰk����(��WB?yp?\�+�R䮝�u�"�Г���'�|��ۛ�? B�(ቨ��}Lš�K����R~$�^�U�Sd��}�z@
.m!c�wYT^y������9����f	8��&K�M����0���"�4���{|�ؒ�9x�R�'�z�_�(��T�V.��pf��>��4��hRS�В�i�.ߺ�-�fͲ��P�t�Q]).<����Db���&"���I�LA�yO2͟4V@����޶ۿ���'��O�����^���S����7���͠z}���*�:el \c�)r^�*��$�e�@��ŉaH6bߥ5����!�ܸ���8s�>��'�W
����ϣ�p���2`=��]@�K*G*a���xds�|��u������$t�k������r�C���
�������eOf�9���;vt������#Z��4vr~{R�[�}�F偁��a������@���k֥^��>Ш\�ma+����� �N2�W�2y(�ďhf���+�'T_�;>,�5��<�Pbk�&��fT�Jy��Ľ�Q���(﷫�T�^�aT�f���V�>,��3�g4C l��o75I��W3#{�L�X)��etu�w$璧�v�=�o߱�9�������cb� �sy�B��E6e� ��dy�p	[aT�G��qF�6���
t�nK9vS�N�V�=HN<!���$��w*'dJې쒧�]����/@��u7|I�h� )��`�G�c���W#)pC�>����?���Y����������&�4^�۩�E?ڡN��f�8�խ� H�>��e�!��6 �I\p����9�r����õ�t��֦�.��o�uS ����!'0s.N�Lu�lg�<�1ꄊ-yEeut�oP�����C7��\P���~���r'3B���7���CaaT�Cx:��޶��x�>u��Z]!�k`xH��8s��+��9�Y����֜ez��;��� *�ò�~�DK���6�M`<�e"��;P�-�ʆ�wM��s�Ld"*&SZ���ֻ���1��c�l���V0�i��Ur?U�Cr�[r�ئ�x$Oa[���Ӑs&���e�`�\9^�"�Q ��?�>w ��}�g<�/Y�
��X�n ��\<3�*M�ͥ^�4��+`�n"�B�0�i{GA=�t.9(B<:_��k��n~�Z6`�s$��`�Rt]�� a(���遍���Q�X��]��L������,s�r�μ �
l�(8��<f�TȦ�ࢿMv_Vu
�0~���=� !�A���Y*`�&y�}��*RN��a$z�zb�����Ύ�ڇr֏�������X��[8�?Sŀ�Z?���f*��Tik�+�� N{���ע;���\�_z�8h�:�p�2NR�
����>�a���j�f����i�������m8�(S8�&���C�U10��i:��`m�y9;�����zf���O��!t��࿾�>�.�YWm��D)�z����v���F�F?�% ������p��Ya	���3~�������BÀ$�z;�<��3^�|e&���#��y��0�	���z��Vd��?�wr^f6�O�2aE{}b?��"��w뫩G�92�E(Vbqa�M��u�P���Mh�@����|���"�_�f�fO�c+�M�����8�b�*�)���ZM1Ɨ�8��� �ΉE#���O���2ӯ�6��l[��K6l+r�0^��q�{ZF/���QQ�FD5�
Uκא�k��*�����	F�S���Soކ�4��/��U�K��h�#O�E3_p8�l/��hI?�0饸�)��/gE��I.P�`����qW/���H"׫��wr��)�a�>��ef���/VVCPU�ƄY�:HK�Y[�����:s�����
p��d䫒�E���|�\	�sI�� nN�0����l��X���H�0��e��	��oͺ�����S�f�m�� b�]��p%2�d\���Ӝ��6*�#�D6,�_#*5��A*�yl�<���,/��s�>I�?έ7�d �����x�g����!mLk�nsVPy,W�h\���I�N���������w�V���OT�+�@���Nj2��AB3[�;�Y�`�]2Y�1�����]g�Y����~@L��|��9~�W�����O-T�z^�m�F/|�R�\�=�P�>��V�@��w>uJS������fZ��M�`����>/d�6�p���P������ĔdM����ђ)D��������l� ��<ܩ�YNUT|�Mj�(��|�����T�c|�6y�:��S���[�D��}��5n\W�'X=YiOx}3�g��77.�i7o��3xR����[��
+S��A�h��B'y*w>�UHq3�D)H�,��%��i�s�B�~�pE�"y��
1
�Z��E�:�e�ե��<�nL�C�w.�F���>4x���!ԓ&��(��
C���OYm:A��j� ��B'�����H̹��S�����4E��N�e�i��N�#�7�y�%�?37X���^O	fE~H/w����\�,X|�|FW5:�>6��䜑py��+�+REC��"���֚:�KGD���pq�W��Y�\��$��@�[e�]�z|��Eq$��r�geX�ͩ�)6�T|�$�;>Q+gcS�6�ibJRx Ҍ0Q��p�X@��KH&N��y�T W�T;b U��mw�tG�	{Oނ'��0�W:���rR�BtL�˯��ׅP��W��:ݩ�V���W�>�޴�#f�H��G����h���C2�
�9k��c���OO�8��i��&��"�Mp9p�Hp<��ߙ~p�O�J������с
�]���K�%6���(��E��-�CL^��T��dDe�Y�$�Pr|�<E�
����"����4�����IM܇;Q��yu{���"MV2����Ra�b�"d�16��Q�6�Z�؆_u������ך�=�exu����U������dW��~�ĵ�qa� �:� �/k�dߤ$9�
q��3?�yjµ4`:C��ܑv��a��o�Y8�K��"�ې�t�>�������P��Ұn�l�=L�u(%��ϣ�w��Q�����AX������ۛV�zu��De*o���B8OD߄��S΀�uݮY��\����f���!O[��_�1���Y��r��\�*�f�r��Y��X��=N|�E����IG��Mn�:]�R�p1M1�\ZD�#�$�	]1͖���@��!\x"{n� �c� I�:V�������.K�DN�X�-��M��$2���T�s}��ļ'Ф��n�CT�hLϑ��6�ӄt�t�IP����K�����z!_�fK���Xqi���x�K@+|
���U�(k>��#�:q����n1�ei�y��o�%P��T Z��.ͱ?&�#p�p��4.��w����9��$�;9�ѱ�_r�(9�tu��Q���7fE��t�ss�cyU�n�^�{���V�$:�voC�x�:	_V��5P��6M�I�;��q�,�� �i��vý���Q�Nڄ�ғ�H)��*�f��F��=5�UO�Eh����4���D��%P�f�o���{#|tKN�V"h7!]X���2��H/#�Z�7���9FL?�ˏ��^�"�7�1��D�Ъ1-���S, ���P��Y-Y-MW*�/l2LG�`%��~���5���X�� �v>)#m�6'x�)4ߗ�FM�=)�N*<���D��)�Vj�2�J+�S���v�x=L�i��M��c�Kf񔾻���r�2�ڴ ^H����(�/,R����obaTxX5�L&Xkjŭ(��P����Et��G
��GGV�r���@i�0�*���248���i�d1~��f�~t��ݾ���ulA���/%�@k�4;��<�*�����\|7�����!B<Z�X����O���o�T�l^��s�t�5.����w��^g"��2dN�eI]��7�j���H.���1W	�o�w�Z��5�`�v�׵�yϑ�ow�gN@'8�N��/�"��(�$�K����^	����1{m�<r�!��Ģ��������j¾E�hұG[J��Ƨ8Ɨ�И�j���6�}�;Ϙ�(�V7�kA	�)Y�Tm�qi�
tgҸ��)���(���bK��q�Qu�]EpD��E:��~��H2�#A�F�6s�["����4���>Fv����͛`� ��p%��'�u��+��yE�p
9L1�ݹ�NtZL!c�t���R����0�YJ�xQ���ܪ��c�]r��I��{�o��S �k�L�8�$%b�m���>;@��=����/����`�V��G���b�f[p{�EsKGʠt�$��S��s�*#sB:�QxG�Al��C�n�@"�hwܪ|���B��&ِ���*`%Ǖ�V��p1����)JBnrh%��+p>t9)N�����1�3-��R~�w"hkUB*�ux��82�F�5�RB1���L��_!�
���J9W��B=�<]j�?��)�#��Q��D��-r�v8ƽC�R��t�/PP��^��^d:�E�������N��V��fR��l�H�����fw���Q� �k��T�&�[���FI�ݬ�K�VM,ݔ�����#�6%�H�]��D'�>�G:~��0s���"{-����!���K���V��ܑ��?C��"y�j��?�!	M��p���]6��9U�o;�k��M��?z��G;%_D��7� �e^J��y�⤈?L�6q�� 4�[��(J�<KN�����<|�A������`�I�|�ǅ����
��׃�Kw����(���77�b��y�-�v{9�ڷ)�Z��a�0���s�"M�
�
[�Ut'���l�7\;2�J#��e-�H��A1-�W�c�}�C��P�1�\�@��E�i���������,8˖��3R��@_�g���bT�N�ٺ�Iűp�M�?�i:5�H5.��!Imox�߬��؍g�� ��$�|�x����> 9��r�^�+ơ'@"o=��G3�E�e��E�k���hN=�P���d2��i\'\���a׶��WIBX�+k���Y����19�� �u6�w�<�#�
lS;/-&�����l9? ��CŦ�2[�'��"E�?k�]�b]��1D�9x6��8}�HvA'�U��Ԍfc�jˡ#�,#o�Q���MB"J*����}S5�qF���_�R<�}t{E+�BP8�x��޶��ɇ��̇5%=�i�4H�c7uŜ��MR���ʻ�s`YMȡ�� �IeP`�&3�8��~J��@��{J��-�V� �%��B9t���"
�d�s�ܺ:����طGs<A�MЩAC��S��MC\=}YT�[�E��b��V�ky�R9B�;�Y�n��&���>����ty"P�T���,�s�z�j��t'
��ưwKn00p�7��Fw-½ 9>-� 8��'�\��iϿ�2�R��C�{,by���)�U*i����-���쀇�S��f�`�_�J����_Rg�;vl��{���MIP7��9��ؼ�^b�=����cW�R$���w%�}��}١��G���KP��}Ӯ������F6�5��O���`J�㌣���S6�?΢1I�g��5U��!���Ú<}�9�&��Z?���ʸ��\#!5̤.�զ#��SK��Jw����pd��b��f�p�w���?aV����4���K�g\�1����r�'�y�k�!��w���e Ԣ%I� 7'��x�$����kP��2HW��a)���3�ʯ\	9H`�C+U���E�ΪX���KNp z��g��j=c���.xZ79���q���ݿc�0����m���w�b�IW|oSNF��
���B^/���:O&WSܣ��e�c\� �['��_`q���-�@`R��N t�V$% |�ay�m�K�R�EV��{�D 6��޿�IT�.�4b�0�'vz�1
 �~�:3 +�h-o;0[����~ǶA\D8���x�ιZ��yK�V
5+�d��؍ �Sg�P�2�I#����1:G�I���fV;s������M��q�g����n	 ���JM����yu�\i��E����'���x[�i��U��:�"�;�S�cnV�y����:��]��[|�����o�&��GKi�TP^T�dUؓX�e)�ֳ�9e���z�I2f#�C�\����d��V={.c�;2i�s��gJK��c,q��{��L~lv�쒑К���\pQ�?p�da�#Cj��e�k�T�c���I;[�wr�$�>��	�%�B2��~��3n�k����m������v�a.�߅�!5���qNh`���ж��$����r�?�R��4]����YlK�*�=
q}�)�N�Ј]`�t��1@p��q�*�Y��Z=S�<C����YDmw��j�q�V��f����;V����iP^';,!WXyGU~4ٌؔfT���6�%s�W��8L�i�W�lXD��c��,�J����F�$��ȗ_<v,a��-��_!�SК�G�|J��V��˃��%���ey�UOlW�+9���1Tǿ�[��3J]���[���T�DP^Z��7n#���p��b^���iW��Y���)H�	��V8(V%��t�H�=Q<�Ȃ��?,%�0�Ku2M]��b�l����%V�̾�R�JK���B3j���W��Ν�����y�3���E��ϊy(U�d��;��3L������a_���֘MK���7�oQ�۩���h��@�˞#�5U��5��deֱ�,�y��-��@��[z�����j������ƞ�'�u�?� i��l��4ۄ=ʹTB�dhy�|�Y�.�!TT/���ł4[c1ړ	�N����xSh�4�5b7~���\��!o��&��3!�V�7�"E�h��Ej
�|6���,�	@P-�5P�U�ue�K�$��&�ڤ�z���W8�}iQ �^ ��m]0��*f���1V��1��g����[*�3��lD0�1�@<0;0$�S!�W
�ng
Z�zӟ	'pQ�u�ٟ��:Ʒ�z5�	+���n�;�136 �,�l&9����H5��XK�	����`�����A�Y�D�蘏X��ʱ:�������n5��~��$S�*ڏT�L��� �ɭD�CUm�-agk����^l��q�,@�`�"vfE�	:M=���/���W�mcu�l���v��p]$K���#����`iB4���>V�nT��Q��l(�Cit�1�7@�v�+�0�������nT��=�1:�sO<(��Z�L�R���<���E�=n�Jg����	u��~0��C���8�1��Ӥ�&�d;�A����j��%E�k-�\t"�m��T�\��!Q
@0�'0�,�r#e��t3�)�4z����6w�-{Rg�c��\�x�ҧo=��[�IU�9ڔv��S����p�v���Պ���C?��cY��ǈ\���J�d1cdl�9zt|zQ1Ⱥak�~>l���FV�;��E�����ב�	G�J�3y!���+cU��9����JǇ�~~K���ثQWnʺ�����]n����H:�ZI�R�z^%���@W�����"pz��}��wQ;��ݷ�2��x�j��{�,�h�Q�G�δ�[Yầ����~{!7��mS^���#��.D��ZȖێ�wf�Z�G�&�_�]�%v�J4����$'���=*��B�:Eg-�H}�J04_�,�P��0�]d��y�р^��ܡ ��'�h�����X��o��?J1�ȂO�j,0��nG73=h%����L��f�8/]x�;��Pⱪ�'#%�Z������bIdڒ�3P 
+���K��M�1Vջ�vFMT?W�]�X�y�#ν^���'�u:w� �^%ߌ���\��-�-�\;�`�D9\�����ֲѮw��JaЍo�'�L	Q&`Np}��^>�w��x���{�캊�o����K�/��4��p*�ŏh�$5Of|��)Lp�F`�O@�`5S�����Ǽ[�2���L۬w�5ؔ�2��@��tuH��~~�07]Z}/�'\m�Cq���z����f8OiN��a�Ȱ�J37�C�*�{���q����k��Z ��=DCy,#�1��.6�O�������3̓�'"�ЗC�a���m�ٯ���l�n��$<�SM(b)o��3}��x
�����o����V�5�Q��G�����T������`s\�X�ڙG��'6���7V�c��L-\C���!g��;P\�"4f D����-R��:J��&Cio�"5;���� ��SMD*�NJ��͍���S@�$�%�p�~��)�#\������������G����`]�Ή�$qdc���:���к�݅�"�[ɷ���f�#�����S�DρHP�)��Y����1�'�k�<!/e&	i�g��@��;Wƶ�yD�y�Ӂ���h���W�	p�G.4�iـ|GQr�y�U��6��"�WI�3ߡ��B����Ư��_�0b�Ύ���qX&����zN=����|a��$��6M6���Xl�8���kJnV�!�N�GS�C=�fD�X���6�}�}�-���K���0��L垲)�`��R���v�z����[T�����\��E�Dt�6��Qs�EMN�P{](�0q>EIa|_�"�G��ǒ-�+�)$�}����n�g�<�W�8���kQ�5��g��AEJ� �E�	����y���o{C������Y<?`�Þ%��SVH��ã���MV�~*Vb�"�A������!d�WG>"���%���~�wq�d\�5�s�Ak1�f"X�ZŻ-�����D�|y@>���a��T��͒��6^\��S~��נP��ax�o�9�nS�f��aK�v��j��oLR^S=���|���=ل'hR�gv!@����K/8mZ3��J��9��nf�;R�D�E��e_E

6�ZJ�?��`�ۚ��{�L\��y^a���{B��+[ΉȄe']Uq�8�Hؓ̈́a�+�Da��V����*����.�͎��_O�
�i�$���&iǶ����*��Q~[��G�8�H;c�]h�H�!�5`8d�l��#��iSM��b��jeʩ@�0��$Z���ˡ�g2����wP�)o���̝�h�©�@�I>RiN�H�r�M��Qԋ}��SxN�4�nz��`b	�+m�����
Q��maw���\�pq�Ov�xNh����5�c���@�(y�/�k��G�6�<L1'>�P��}Q?�m[�#o!�r�H�D�ƀ�F�: G��&%�SdB ���B��6���OIS�X L`+��M��h�6_�=5��a5��3@T�8ý`X��)j�Pu�Pfg0��7���ZKBÇ�xF���ݪ�'�Z��%ZfNK�ꁴ�M��<�'S9�#L��ɜ�c�V�����<�����~�`@�]4r7�-x����4k�O�� ��MCGt�A�3�lK�5�T� Y��
o���.����;���T��=��ǂ�PF�`�t7[Az6��|F�)�h�,�M���]a$fv0�ޤ *�a�7����W�}����#Q���.�z��܇��ߣ!U)`L�Q��9�Hx���e���M"� ����*t���p�d+±1�o4��
W���?�y���k⏏�duo����֏�x��8xl�����{�&<��W:]�F�y_o��;�Њn�p���=��N��j��Y/�*�t�5ֿ���Or��|��'���Q��7�h��=�j����mz���S��N���Y��-��O�,
�K��ʯ.��?�W�z��|�^�z��j�"���%� Ae�5l��U��v��	z5��t�0�D�h+��X�c�XO2�I��}5��<vl�I��z
:1
��F�=ux�U��p源=�6�gl����2�Xgi���޳c���Oc�lcM�w�W�1X�_�������#�馮�����sށEĺ�%�|���O��^�h��.��m��i��7dx�H��1z:�T!4�N/vT�!�� ��oQ7K^k5GU_�_^��$V�g�K걘���/kQl4[�,T�WS�%���<>�C�i)Л��ǟ٪}�W����'�{6?���5�ڣRe���3��΍|��lc�Z;�2��¾�9y�F���Ȯ"��H�T?k/�8�#��e�.�n܁v�`q�j�ѡ��	:��2lՉS��cu=�Z��⫚Jsc�z��)&��ml5�<���.R������z")��KA� �=�g��Xqo�ۧg���D�c�����K��D@6��l�"���#��A���Q�OqA�o#\�A�Y���F��h����o�|�_P2(��/O _�@'��{ ������UYt�G;$�R�~�A/EW�%�A�b䃰4R�3w�K���_u{�"�Ƕq����=sL�������ġA�ܽ��f�#��	�%��lI]:(�%]O"��Ӆ�'B6k_��]qtڿL�z*
];߼xLb ��9���A��L��y�#����;���i������^B�-��:r���ـ;��\ശ��
����{d�g5�Q��>�[�qA��nzE|ҍV��"m�0W�XE�|�׻d<u#�zG�
`+��F�HLn�w(�~q �u��T9��Qt.>-҄�B�s�.@��Bg��g�@���#G�%���R,$�Qc���t����us"�x���k3��'�-�_0R�o6),��h�y!) "��B����

7�1�ay0.�E�5P�M%W/	�#{�.��|B�V>'{�5d(��"��uX�Qʊ4m�%KJ�xcl$���Z
%���# E@?�u�9�W=��2�L�~�M/�j�j(�:9Rd��2���9�V'&�a*>R?�ق���>�y����q?�>uC��1u1��f�p����#j_~��͎$83�~EU�F� 2�\N��h#�[d$����{:J���B��%�4+5Q���x�.������
iK#jNI�-�uz�*�i�����A��oT�.
���Ի���=A
ؿ/��w(�Zí��:^ө�A�ۙx@�5,=�^~��	���X���7Bc���y��&�]���h�S�|�{��P��}'�'3�A��)��e׃J���8���R&�hy��m��m� G��+.��4�~3�1�ʢ���K��2�=�7����c`^)�h��*���q�hK����+�ߏ|TWT]�_�·Y
=p�V��ED�"h7�a�
�z �V�4����G��U4<`��8��;��"u��E�yd��0�����+��B���c��������f��*ALM�Xv�{d�K,���̱`[0���踫�F�
�AO�:�Ǆ��Ec���4����MII�����pc���>����*��+���{�pY�3�tn�	23V7Q�d#?�S7�4�t��I��gj	�}1�g.?[i`_�l�H�}�V��= ������"�0,������������	x�Ϭp:60�KO�3_In��H�L��T�{��8q�y����2��q�R���������hD+�l���5B ��ڶ�#2�%=�ǎʁ(�q_C �`5�|N.A] Lӏ��x�X[p�E�<�u4"�V�b�M��B�VD�;X�u�y �
;����A��y5��9�d��vˣ���6s���Gg󩪪,���$[�l^���
6<��Z�3���C��`��b�;p��³\�:3J���l�ɝ�9�A��N8�$b̚+���yڌ�D�K�5oKL����P�?
�ـ��ߑ�[�O7�͜I�#9�����F�\K�mIJi��`6$�R���~��g`h��+JFޢ�=��FOHd����u�0���+ݟ���i��8�<����c���C(6�`D��k���ͱ�d�s.'~��[��#�(�Y{#�5T�I�?f=���s[N�������G�Y��8��~����`�rv���v�r�OE`����"@l�e"��`��4����΍���v�}�[-U��b�_S���Q��Ds�a淲�����_��"��A�
dc3ûH�;򥙰�(~�6��%�ao��jQT�E`�*y���uy'9H��a�:�Q-�f����Ú�41�E��[�{oç��d�r޾Q1�d~ K�^����e�t�w�1�ɑ��u�N$;���m9:��H5�m��uY�L����:!�g�������h�:wC��^����W{Kܼ;�SƼ����]�)1�#t��Z��� Y4����V�y^��Rُ��81<8�e< ��oj�;�@�t�<qY?d�s�_�s���Y�Y���#���k}��e�o���l1"����s�qG�:`�cx�b}AǢ�yB�R��>AA����X��<�{W|��x��9�Q��e⊯���j]�����)r���_ml�)hx�0��
\���Ձ.��,L��@%F2q��S����YPp��m�:�,�\��&9�<��r˅���6��@�b����T:sn�Ot9K��_��.]��_,|rF�I`W�QZO�a�r��T�83VAۚݓ9X/a���wXT��Vs�SC�����fS�i��!$��ѥ�����1���D�����u1@��}����>���������g9$�;#�˿=���?�_�ɇ1"y�ԥ!.��,R����8�:��+�UȆt�зiz1_�������Rh��z�#�#�i�)��Q�����X<Ǚ�����/�o�U�3;��?/�3G�H��G�m9v�X̤�9��$�1< $��ւ���`���T�������A]� dk,���GE��jBeJ|	�u��ہ�ȟw�&vD2���nn�<���_�>�u�����wa����k0�m�Py����1F��uC�}�`'#S�^����.)#������ZI�TQDu�;�޸h��^5��G�jq~���eD�K��2�FiLG2�EOc˼��V��j�Z�������j����[}�r����m�9O�u&y"��⁫ˌ�1���C�C{�����o�c)w�z��0l�vA{�1Ù_z(�s���6�̙��X�v|貪Zg�eJ�T�^�"�x;}��8I�v�\��młc@3E�[�`�{	���PAK�8R8�Xˮ�@}�XZ���"�:���1�:�mD'�Y{}�[�����ӣ�<�;����.�~��&j� �9hn��|���+{��۾8�=S��_�oML�7u8�q�Z=�trZ=<���8�� �gC���Jz0�z�k�[}8�*m��<�g 3�;;L{I����>�W���L���ee��L�D� (B�a7�mr�+��Rx�
�3\�l�.��*ϾRK�(�M~�%�3�66<g����_�D���C��6��)N��,H�ޤ{�R��1���Sl՟�kdE'�#N�G��D��y��\�<�'�ڂ��[l $N�?�L0C�6����<�$I8/�l�纅�2T�(`wFU��L5Q�����P���$�����	N@������a����v��a��B���	@狼��sp<N�F���]�E1~�wK�EW�U<W9#�Z���7��/�d�S(�! ��iqp4�{Z�g^.s~q�߬��ax����;$�HԪ����ך۳$����}�^��-�4p&��, �z\8{V\6 ���m��Qo�9���s������� ��}�?g��w[��ehkI�N�KeV켅��g�[���E�0���Q�L��p8i��]X�����f6�1=|&�ˌ[H_��r~�&�Iv��u�Rۭ8�SPs��+k|-���[�P����� �x(�$���k�q�_iڙM@����t�\jI#�m	x�����C?� U p8֩y���Jh�!���GB3`���襈���d���7����ی"���ɲ�=)	Zx��9A�f�,�n���G�)y|�����o�s��=�3W��S�e��df�j��9��a��h�ߖ y��Bs/��2�a�{�tM	k%�=M:"�*6�`�V~�fhUʘ�*�>���C7��1���,XqYU(m�bW���E�	�����(/����U7�Rר��]�?��zn
(v���}oIĕ��w4������te?���(o:	��ӟ��=����:�l��U�Hb�P��.��P��3J�P��Ӥ��*y��І�I+�	�3��� Aүo�D���]�E��O)cQ��������μ�	�܁g]O�lZ�6 �o}����/�N��懂,��.�K��d�?
������:vTIx,��p������{f���JȔL�)��
��0�9g��M��vϟP0��4q� �xA����?��Ӷ:v1&��-�5҂$���Y����w�0�� �<���fE�0A�ZkU�(X+�h#�UA��z�mkn�'j~�&���&�9� ��S�f��!EZA���nfى�X���r>P301�{��Q�d�)�T$xey��el3�΢6O�~��!S�V�((���5'�6�w��!@����� �ҋKZ��j�S�G'��M���Xݺ�pS��웻pæn~ى�p!�>L�1j�P;��Q^����wf�tbpLNR�0��}Fm*7���F:�RߐYU2�(�v̺T��0�`Ry-���m�*O�a�����|��-�Nx01�x�W�ip������2��X�DN���+*�V9j8���y��|�o���m��u�.�]d�?0��Ө ]���Z�W�"�DU�QFܤ�D�r\���,�Y�α�����G �o��`��^��ہ���?���R3�Okp%�ų��O�j��3�=�Ƒ��ކ�"�K��J�J�=��r�|v�s�
�n��|(��КZ�(���Yp��&�c'L�&O�WQ�T�/e��8�/ �ڰ�?�xء/+�V����[��|�G�$13	w4�v>r*�� 6��>3���=|4*+X�`��Mg�YhЬB�V���ξ� wbŧ2{terx%�[�cv��V�iU!�/�`�U�_������/2�]��.s(�B��m���vI8n��'z��&	�9*c�rX��m�;&E��m����'u����|��CJ���u���#�y�#��o�bX�K�����17f�y��Ɯ�"����ޜ|!م��Ǜ�ᒠ���z� ��Q����P�@\��l�[�:q@2�8�n� ��� ��՘ʹ��A<N�������-���s��q��#|\Φ*�
��7��R0�̭~MPO���s1��Ad����g_8M�.d��4B �����v��_'i��y��v�E\
;����}	Ma7󹱲���D*�^7y�c���$���3G�F{�
Ha��v;^:ll����l��y�]�j�ݦ:�e�O��J��	�.��s
;�7%�Ϭؒ��l:u곣Uj!��������S�>H%v�
���4���8�a����f�_&�`����hdS�9�0Q�̘�f�& )5߇��f��?���EB����� �����s衶�D�f����&���Q��SA p�(n<1K����I�Q&Ҕ���G1��f��STv������W�c�������ǃq4��T@(h.�����&}�nM���O����V9B��H��?��/�r<P0��י_��RkV ���(�Mrff�$ހ �J�9h�Y�Ud��~�B?U>����*��<I��G(cң�7�-N��g� �p�V��dD��'P�079��m0-1�ꖂ��ua���ྺ	 �A����Q��qx4��Y/�S�KG	m�R��)>K<���)�rH�6����x��7H�Zʕ�Ko�J�+X+�4R>�3�7(�9��	&4�G���� �yw��6�v_��������e����8h��w|�(���bw�3_L&Qn���[��Cd;,8.�[�u,��
A���^���2R8<Yp��F�����=1_���kk_�R��՚C�ѫ����*c��Ɏ�֠�N��*���յ�1
l�g�M�nu���6�$��$�$ �+]��.�OEo/�<E�6C�_�Lb���Kݒ!����_d�p�(��oa�����@�~�K�s�����Q���;<MH�'/W_f�@�|�Gm�@Ǽ�j����C�Rt�e���H��*����vQ��LE1�H�n�+i�"k��.q.�Y6~H<j^�x�f�#Q~MU0A�"P	0|�q����p#S�ha	��G�`&���~\�6��SE|}�eLQ��㍏�C2�ZOw�QR�Hцe��u�qC��ge�)\�Y����0�ە�����0��mʯ�h��d ��d�]�B��T��׍EvO�j����%�}�j�T�����Rڵ@��H�������-����&Go�������[���oF�9,YU�{��7��pH�\�^�^A}�"v&�N�9zl�Ò�cu3֟���^q��	���JɦR�b�����;�fH�3^���c/���B��Y72�^uE
+���f���Sm�"��k�4i�<fd	O�$�Z���P��]�EO�tM�ݫ���E��Yǀ�Mע䰖3a�Ȗ�����e�9xb�j�ΰ�ϐJ�d�N�A΋��y�پTrB��Xz��g9+k?�#PzA�__#�ha*88ZsȻd����珮��<�k�R�g���Fr=�c��U���{����i���ڢ;{[R6۠���d�Z�s��q���_��.�X�ƽF�o�8oQO�8"O��^��ZDXo�5���N8�lKG}�,Wn�.u��;��O�s@�"���%kR��J_։��nd�}@��iC�zz�R��{u�̬U��F�0:�֣Fe�#�~��<�zEy �W%��u��ט��O���{y3�����}�9��Ϧ��ϟ��'��������BFdu��2�� o�y/���[�~��� V�K���Y�Ҕ�C@�?j	-�^��:+�V�r�`��u[jŻ����7ΨfG�dw��`'��l�'�0f����;sAFG,��ȓ廵���Q�}s���e���0M�k/M�`e�o�H�m��ݗ���ƚ�Q��D���B&O�>8��뭍~��ӽp݁xn^,�
D�q4�FF�`�J�ʒ�����h��ΨO{��9�!��{R	�'�J��2�mԼ�Ή:�F6��[h��Uk\n�n�5Z@bc������0U�KԐQ	��]9;�2<z��u��_#)d$@��V��K�(���l�� �B�����,���A���_3[�,�",�z��lV��#��P�R��i��:�`dA��i[��mML�,��y�Ol�g��C8F����l@�O\�h��s e	�X�ط�%c�L%�nmu	F��C����n��ȜJz��z\2
h�%�Ey�?CA�k��Eȣ�:o�LA�5)�F z)��u��Mޢ*ν�"[�1�Z{(�;x��{*��@?`[Fb��:=`%�8� U�vh�;x?��\����8lw\L��8�" l�Wa��n��Rt�������|��� ��ɇ)�ˊ� 0E�K����g�&���*�{��4�a���O[>5>�������0/O��]'4L-���q4��N}/��޾n�{��h>9f���:��y1.�)�i��X�!�:�!eG���X�O��X�A�~&yj��E�@��#�<Y���Y���tBौ� ):�����8�ƶ�
�,���j�t	>���츿�L��zE�b�/Jy�7n�1ݫ���׍�A|_���'#8��p��4c�g�@`9p������������	�M�YE�a4�0��X�1�:�QUq߲����h78�'����\x93��m�Nh�L�����4�q��M`JwZϾ�n��]�2PCD?����׶6@ b& [;�����ƽ�^�1���G6��3��ґ�DU ��>|���Iz�O�Wk�{��z�þ����'i	�r�����83�[W!w���������SS���Qr5���nX��yX��	(���5�����l���y|q�$���Ĺo��� 㑪CӐJt�t1�Pa���Y�{ �W�X1��������NB���"��u������l	��L�d�;͠��,i%�2뗉M�w����g�`(�.��P/~e�� �Z�N�φ���K��"g���c��U�[�4�}�CF, �q��f+�'i�m�œ}����lp���sn����0�2���z���Q�[��_������6�T�o��e!�2H�� ���s�u��wt����=Է��bK��d@�:F^d㊏�Ӟ�4�j3����YDmʃ��ˡ:$��$�}]!d�ǌ5��0�s��1����IR����%oA�db��z�@L8�n�R�~�]�NJ��l�iW5��^R��M���hw,l�����ŐH��Uo1֚��8�E��p�]�"1`C���^��F
<��ʆ���M�,�Z�>�_m�!z%��&�kO�:� 8�J���%�����N�"��$Y�bo�3ќ�����������!^ep��z����HP�ʛ2yq���O�e�w�Wd����,B���FD���^袶�,��虔��͇6Rd�DsQ�f2
~�"����z�z6�l�����p���0�l��T����I���G��Kyr�����lU�0f�<6f��pC�T���Z�zT0~���{�k{�vi5����c'�Q3�kU攜���DI�R�]��&�����9yu`�A!�lu.��ë�H�%IiQ��jK1�N D��q�Ѿ��>rؒ�9b�k� ��F�B�M��d�=��+���V��P:j�����'�|���v���`^P^�\ԁ���+r
)�T�jPyޟ]Ȏ���@�ѐ�O�a��@�o�p%CG�~�khyi�GW+�vj�¯�6��-D����2�@j3��4ZA$o�jR����n�o���@&�����M��Q"�<Sx��dC��e�C���4D/�`*N�8�����Ⳇ����'k���%hԲs5��JO���ع�p��'��ߺ� ~샟�U�-��-�,2Yb�;�pF� !e��ޠ���.��o�Y�W�-���n�=��>��pZ��Q���B��už 3�M'?vb#y&�/��#e�/��W�<e{lATջG�G"P=������'�V�;ê}��}O�ހ�L���J�0�}����᭔��Dy'%��_,�!J8 ��Ml䘽L�1���龕�i-O����B�ñ����jt�M�H٢g�t�ǦڍR���Ӻ�����R�9ө/h�p΍M�Sh���9eR�-r���+�� �q���*�.���|��c���;��8Z�"��5�i��m �M���>^�%	�T̓|A�6����R�$�{]�-��(Ŗ$*��%�0b��~!{E�c���ۤ� � �q�r#�L�mY��G��I$4�9��<vBHd$-D>���%X\��\Cڼu؟Ӌąg�5����v��Aʍ�V
��v�pF�u��#>���w����q�8�G��.�� |��>�����h@ W�N�ϟ:WKz&�̶޹�B�ha^A����?��.o�Q(,;G�߫�`�\2�\���r���X_���|C_8Œ=&	�h�\ً�\
a�Ǖ��]DE�i�j��R�{L���sw���_&we�-::is@�����;�|ԻX|�6ǰ��wd��Z�0$����#d	v�+����/�<��*��3�چ�>)�NV�IŨ�ܡ��t�/AG �D��h	�{�}�:��?��xj�W]d��E�6�_=� ���|��Tvk���u2)��oË��\�`���&�^���yĀ�CJ�OK^7�ɵ�-�&?>=�D��3�*(�<��*%#�Z��EuK[�9]��4��� ��V�濄���9�����2A�k};J}�e��ׁ���ߔt�Ϲ�M`�,����Wn��O/|���P��l1�y�뤭���hH���Җz��3�|��D�Z�s�92�l~k�����-��M��J�����o���EG#��������\�aN��ϐk��֨p��Wl�����z魹un�b؆D磐�I�Y@To�8��FW��JK����Cܾg�s6_z⎜@�a֋Bi"ׄյ�IX�7��wPd�����O	2�r{�����]�8�hL��%�K����F�.l�i��ui�=���#��~��@��lN��,VeI������뙁�}r��hV�⥇O� tM� �� U���Y�e��	�� � }��KD�Tb֖-_O ?$�w���g;jS��F
����W���ˊ�2h�Ҽ��*�z	�C�J�r��p�xyv)���D�W��iP
,�6���;��@}���Ej`���J�jM��7�`������gb=aM	�Ue���e���C���u�*�����8"�[dk�HW�U½�P��Mk�Lo u~�,>��^�7~o�S���J���eg�|�]�GT��9�Y,"�G��De߃�6dXK�D�1��B���1&��yO�n�E�q�K�
��EX��5|F�W ��*W���O��W�%�'�|����*H��;��k�</�"R�_A�э(��[,zOb�1�}-����h]��X�M09�p0��]���\��GqO��=�\ �&˓�����@%fE�ZFɍl�fQ���.[�wh�|�q��K���98<�W���Oד�J&('�Cݭ3}خ+V���M���~>�B�ɑ�',6����h�d�t�i���y���1�*�ɉ�<������Qp�(�i��TGLv��eҦ=c�j���.����D��!��ӰIf�;�?�
�b���e�4�L�n���z�r�c^BW�;�, �Et��(N�?���x�IUM���+y`2b�8�A�ف�^�l���������e%W��岻��\�f}�d4m�~[
2���O�"���_���l����ϡ�=Th `+� F���>�/0�n�0�UEʹ�c��x��C�$=@��WX��
*��	zt�$`s�j15��?�<X��MX'�X�5z��z��� 0r-��]��4W�ϒ�5��J��G��|�t�)��3ʷ�Y�1�66	<���K���6Jd'���g,n�-ZT��f_�\/b|eU�lu	�C�;�.XU^oO�R�6�,��?��%���.�\��m�t�?������Z����y[��svL�`(O�-4����0aY�\s�!�XLyf�/����3VQ�ی�T�`l- �=��A,�H����\�Rq2>_p
8e���(e<�f�	:�柕�1�H��6���ղ!yIye]�\�J?�5y?����Ca��Da`e�*r[�C�ã�݆��AZ����=����ք��؝`F�lI��¡{��0���d���b80c	�z"��ir�ʰ�R[;�3��'w�ч�jp��($�^��\Kd��cto�� �6-�y�G�
Hs�c8�oC{qC����E��:�P�;�eC�o�a}��3� �ec��']`��	����6my��f���[|�mP�f)%-��� 6[���ND:]����+Q��ϸ��u|l*P.�We$q��VN���\o��������	'�{���&E�x�v�5E�3�|I&�+ɷW,�ݖ��;��~n�cTH�VC�~Y�KFϾ��Œ�}`_&R�j1t�`_�j�J�#���BxN~
���߮-���+���>� [��N@��̸�p=���~Z�ѳwSBjk�$���+�C����LPx��iI$1�u�xq��b����<*�MKP8h��1M�!O���i�r�>����� !���TƦ�cN�|��,��@r��D
���-���۔Ic'e�9�ia3�ysA���>��$1��������#��{~�|��%�S��(����?�����՞#�=�ReDX�1�Q�{�aG��ʶ�8(a�$�̰�V8S�n���b�cEY������U�+��Oeݟ[��6��(v��0.��I4,�ƶs���F����@;]��W8kˁg������Q��8!�Hc$�A�'Ea�]m&Ī+e�6��˧w��-X�����+DS1V2?�3H?��N��ǥ1-C�V"*���V�1(��t\#-&_cU52FP�V������f�Kl*�����03���j�S_$��ܿ�m��Og�T�dMa�	��YB���>�J̶I�\8�������	̀�᭱�CH��p`��>�&�kу�OX��g{��jR�y
��6>p6�x�0(?f։|�;�ڪ���L��x�M֐0�F�?,�Q,�-ۗ�y�M<j�������J�c��l�4��zZ��v�0�[��X�o�x�c��GS�P]�U7\I��k�t_�KY�,�{o��d�(� ��`RO�`�Y�. ��eJ`���f�a��q&�O���D�W�i�pG[��X�2^�����b���;�����ĩ�V��x����*��+��(9�(�&����$#��aZa�"��0)a	�{��u}*�������^�9r��x��	�`�_�z5�%��u<;eCA\"�r���;`;�P�C���g��<"�B'^�F1��Ǧj�|=p���W�~�3h��JT��e�o�;���{�%���!������~�c�E�$�Ւ�%L`�w  H�]A�k�a��x~A�D��4c������&fֹ�W���� �8�ƨ׮B��^5�K�4�Z(��"�������:VF�j��mI9�B�0�W[vQ1'1�l��o�p
ߍ,�A��Q�Z� m���J��&5axM�#��1\&�jgʃ�.��#��.;��L�����YӨ��B�"�PL�)-/J ��m�*1q{���6� �NE��E��f���}�p�|����4�gs���4ip˴�`�aeɝ�m)� ��k�R��y��J/z��C�/EH�_�P��y�<C]g`&��Q�QI���m~j�I�%�a��J±��@�_��[��+Gb@��J^����wR��}�@.��di�V�^|�x�#�f�S�aI�a� ,d�1�VGm�;p[E\���>������f�S5�.X�	⾰�����'m�Z{��h}���M�jt)y]فj�ZB��yR���k��V���%j	���u@���p��V:��I ,�Ϟ�~��Ʒ�����s��qzF�����6�x\;�����=;�"���qqj�Ru��!/r`5�L�S�/�+�����E+n��m��9��l�uu*c{	��J�)����K�z*�W:�=�����Bcs�V5#�ÖπE�'�������VY��X_}���U��ľ��U�o�L¼Kt����,���z�4���.����1���z��c+�3c���PYql^���h�:�����)9�*���p:8�N�>�d�n/�z�V���M�x ���9Z�ܶz��Ce�!��G�X\87{�3�g����et�o�NJ�Z���K�[�qI&�m,���<�<Q�뎑�ljM:�4"ф��-�'��Ң�7�mz����騿�7�3��i� �㚐��d�u���ٸ0V��[�4���8�/\��_��b���O
�=�0�"�99���7p�0,$V��o���zf��̒�W�s���O������2�R"��M��f͂C�<�ٴ���e��=�kêė��}�#�ݤA�`��n�ƊY�d����0w� F����H4���&�@zm k��0W-��`K[��ߝª/[B=d�S� k�Y�p<*'a�O��c��}:�5�s����4�[ ��'����!�Ai���*���K�bz���ڿ�[����c�&����T�$S*�TMY��F�a~)��ecXXz>�A��+�_�P�+���i�����l^2X��t��kàCi(d����mi8l�����}��e��c�aE\KHe���q[%2�����[{�5)��'���_�"Y�qyJu"+��K��"���x�~��>�mk��ᄝՑ�Lߎy� Z��3�I��95�S4D�"4=xU����(+T���ͺ�.6>��� L4S���j� ���MY �Y�ћ��ȴ���=n�9��EC���	$�&�hR�쮭�Ֆ��e�4�]��2PnN�B��R7�Nc�R��?[o���:��;���I@���]��꺖eS����*����NƏ��\��7�c��L��K�1�F�"�[�=M�N�&zP�r^	���t?�i@��4�C�� �X4����/t�D�,�t4�ޭ�K3�F�t�ϪGx��M�iʯy	�*�*����k��ՙ�7;j�k`���Ш�S�@���}s�I�W@�n� ��2( Z)b���BW�i�
��4�\e�x�t�P;�a�I�r��-浖�Q�����v[���&�ҩ�&�O��I �,�$�i�'�֍��e*Y�
�"��M�xJ���!����� �/�$ y�K9�]Qj�s���Wo���n���a��iz-�����X]2��k��"#����Yǋ^�Ȋ����<�j,�YZ0(z�z��
Qf0��1�T�t�˻?�da� �0pL(��X�@��0���L��������U?�ǆ�=�q�\ϡ,:�G�Mߣ�	�GSS@�H�;b\���q�xi;I�5�^U��I��`�ɼ�bn,e��{\�_�|]���t��%�d�0�Ϋ6��T�;�D�@�����8zŗc���qt����uN������;4U}^:���b�?��Hÿu�8%�`ޓ�?���x����G�P�;(-�۔!8k7���	$�#�c�T�!�Owf�e  �|�ﰰ
8�*���m3�)��r�T�\N^�.2��NF������FXm�-��������u����.O��z�$�A2l�}	vx�xb�����l�xK���71�+�*��Ek���Ib�UC��je7#��a�ʇt%^���^��BKmgaT:H��S?�m��(����Md�,�x�ѓ[	�`�q#���c��H��Uw��U<��.�h7�1���'�c�5W�u6�S��3Y�x��"`�H$�?�k|a��A����k�k(�<}(�W@[;[э�+S"�r����9���i�̐#eNmY]�)��N2ω7���T��:!0��(SF؟��Er��T�J%j�}:�}�fh�ƅB���ׁ0-���e�ȟ:��������J8�1��Ž��$�I������`�ff,sy7��\p�I!�h|Z��!/�,�0@�h�hQ�E�rk'�����!�~�Ŵ��d+~��f:,�� �v����y�a,{|�>�R�5U�����O
�a�P�]�\�dܕ��L�͏y^Q����������*}�7��k���}ɴ
*O �b@��C��w����7�Ұ�y�-�,�s���כN;���o�Uֽ�|	��Ja��xh���Z��K&L�e�O골LB��D�bk���$J4���F?Cf�W #%���T��#���8og�)E��\�X�ű=���g��p_!���V6
a0J|����Q�&7nWe,��G�r���w�-@�H�c�<:�t"���齙g����D�.h�j�SMqJ5�E���R���C��q���qo:5�K�!��HqK~j��pgY�9V�w�4*a���;��4ʮ�^5_h:��`+�}
���,m1��&��T�ػY?A30l_�uiÔ�$܋;�[��Cή��D�7�󐥣�
?c<���GP�f)�"���{�����9��5'�wb���"�,c���2���A����T/_�F�����l_g*�8J%�������BȮiCD�cm^ڴ~�Q��_|�ihR���,�2��̬s��.n�L����2�����n|�֥j���xdKL���hL0}_,V�ꢣ���7��Wr������:�ÜC	�%��,�^w��-�gi!.�xq��������4�f�����-���e^���8cp/� v:0\'�󆿤��0e�!#j�} ��T���w�̮Ј�?r�ҁ��%��_�������֞�ZB,��,^6S�/<�U���m�7Nc%0I�M5��`	6���#���)Od�a�
uab�;`i�H�E߽o��'�u4<���HR�/�W6Ӽ�F����ň'����<,JΔ�p����g�"�קB�u�����x �Ĺ�����P`��u0ﮣ�^L��� �t}�i��v��x娶��	k�fs�90�&�R��(
W{ʌ��=�(�%c�e�|�,�>_�/��j�_5�r�a���|�*�Y�M���/��a� ������2�����)�����I�N�G��' �VഒnR�fPun�c9[��u�XX����P~�(�7$ ���K��B�e�
ܣϐ��ݽ��5���[��M`�_�,=�9Ƙ�JV���t*�F��U�Hz�R4}
\14�����$�;���<P������& �f"RI��'*L���c4)Lhݏ�Ô�	!t�K���)C��,P\@�rj,�/��UQ��b�_6^]A�D����>#�Ϡ��M�n���yD�Q�? S���s�(�1��׮����+���&�D��'�0��:1tpi_��.߸eGL���b�M��('E�^e��r0O:]�GXE�ױ�8~�B[=���YE(�a�bs',����ދ%`bp�)bөϖ�I;g���o�@	٠a\��./~�Sr�-'��y½��R��hAȣ� �������� ,z���ԙ��;ʄ��y;�v	,���d�s���j���O^L���i�"?�� 9!W���p��$(�LY��d�������%S~�Z}~Zc�F�/]��]E騣�0�q����ϑM5�ĳ��h��w;�1�eD3���>� R˱�D�o":@{#�G����j��~���	ٯ�0�Ȃ�k]C��h�z����:|�M��o̞f�����j��Fun����Àu���]�w5G����Y�t0��Z��<�*C���'�(��g�ƍɁdR��� ���Ap��_B77W����_X����O�����,>B��!��V�h!z}J��=
�P���;@�zz��ܢ�2�(1/�t8���Mȝ�~�p
ފV��a�-��@�/���ҝ��#�@dy��rJ�E��b���	�*�� ��NF����Z�l%�ծ_lԇ��r	���24�T$���gC��&q�h��[8a�f��#�s3��0d_��jw�g9�Q1?���[Ł������Q�g�aOA3���	E]ow+٥�?N����֒�%
7w��/����$���9^��,��k���@|K�_�{�#��0n��L���unC�0�;De��b>����!�p�+|�]Wý����f���'�'P�ڽt�_9�o��1~�Y#�#�d�S�E6�E� `	R�R�Sm�!m��2� h��uY���9P�%�鸚J��ᦛ~�'1��RY�Ə�U��<��k�脝�@c(1lK��S'���&F�D��(����R�P��I}~2�-����=F���J�*�Ȼt��1	���:��>�)��'�$q�1��-��{kɖ"���=�̍�vKB�,�]����=���$7�f����a�����sRt�м[���0��W���Io���Ţ_	�d_8�q��Ot�� �P	@�h<=W0u�#������AG�H�10�] ��mz�!|�2��/?%�r���}1
�qP�J���P�j�5�Qj�U�D��rpl��nٝ���ӣg:����S{�Zu9�JH\���c?dy ���ΌXt]
�os���s��<FOqD8Ւ������Mrj����7O�C��ǔ[Q���4*����LXn�V}Y\���� ��å���7�U&c}���	[�;H�YƬg`�R���x�&JOZ/�� c�Cb�	Ki�^��בK�"����߲I���Wɽo�NÄ�;yp��e��D@u"�b;�@��v[x?�f&�P|Nv�,)�RD��S�d���P-�]�Ce(�9>`��ʢ��)'���|w9l$+���[��4���*�we��Tޯq4��)c���/��0lNklgs�������KXw1���d��5n���&�xG�1��#�kw�f�����̶���H�VY	M�sgਐ�]��cOU���d;:B�!nuJ3�C"�*���S�ď�,U����=N��xLhi���� �lLw"F�]]��W[�8J�]��Y������캡:�W�9k':=�i�F��E��H�Is�=�<�\|�s��*w���[����{]���0�?B��.8��B�(�:�}��dIЙ7��u�dY�z�lL�'�x�Ĺ��H��LuI,��M7�P����@zN����C�'V�n�^l��y3$ʲϋ-5FD��� D~��p��f���m �7g�ė��B4�9�ˮ��,CM@a��TL��hN)�I�����r��+����V K*��U���k)Ȍ7�?z�ֈC���{@Y����n5'<�4�1�PfP��J�#/x��s���N1�t_R�Ńv�v�1��6=��Mb��-����� �� �����x�E4l��[�G�G٩�2����":�;��0�Ǿ���fG�A�l@I�y�;�桐Vh5�t^�x���$�]�q��.?ȍ�/�8��Z�	Q����~��~�5�+'��`�&@fR�N�	�M�$|���41�q�{z[�*:�y���Y��ڪ`a|/��d�^���h��G:=�=��qJ�9"c3Y�mO��](�qX�0��M���*U|;�����[�<�f:T��P�؂㩨�6=R��g��i�i��~�iFL��	򋍄�@�<�5Um�XgH%��۝�!����[����9D9���]�������W��s�PyK;�����6h�@�Óڙf����N���k��L^�hf���g��|ͭB�傼7�]��~6����A���Lo�~VU 5C����ZxY��m�������3�*'����[�7I�Ju�H�u�B_�w�Ń[bw ����_b�E����aasA�|���.m�eɸD�cF��{֌Go���~6>��O��"��<#򴂲������81��I�ҭ�ǣ���=�2�
��\��0-��y?���N�H&%RYp��a�ww�O\�����@�t@j`���^MO�'�Ľ���ޔ��j ɱFa�TG?� ���ҜDb{O����l��j���J�34S��%ң��(~<�6��j�V�����B��k�:�j	u�x��!a=���J1[�s�����V�4J{�s�L'��ۄ"Jl�[����ݣ$ �\�H׼z�;����,#S��!;���Y��R�s���]v��n�Ǚ����؇�׀{5�Ə�s�yW�A ��yV���b�ғ�-y��^DO<�pn��v���}�K��S,tk��ovD�!"�z�>�����C[��w3R�q��G�e4q��u�T�3��^��[<Uc/r= �4���?8U
T��įe��l�HRx��t5�R��'hO�y������#k�#c�:}z6	�f�� @C�?��KT"�B�����N0e�	��3��{� �Kh�U�&��<�Da�x���&jSמPi���](����C���C�۷��(O���į�3�E%���b�E�o�sV*�$2�g�?�G�f4n�9U�ss�Ț��WhL�������'_`a.�$� A�	S."&�k+�v���(�+��p��@A�HW@c���w�C��s�(�{+�[~�&�d}�L%]���GY�fåZ����W��DHk*C�`�ל��R�(ڼ�I�(�x)����+�$ /���٦).4�/���&ea��Hy��?��F]O�����;�g�3^�5�7F$�D���@� ;%Y�	<�׿��GUF8m��4��Vti�v�)��%|���&�p����.�i�_��!E�&}��؜%��8�	�������oaOz�����fQBOQw!ş���E9kLY�_ʐ��:��N!lK���5� �49M�_س��~�E�Iq^<��y���ӕe�j�ܙ�r�B%�y��:��/�i4-)߿|cp2d�2���4���Z���g�Cqf#n%�s]�j��ɄĂA�Ⱥj�����ߥ�������wNxR��J�kJ�˫<XN�RF��劸-!��67[��;��q��r�i���=g�%��pӺb�k�M���K&.r?!~<�z����U��ڋ���m.���g	[{��H>��eC���|z��Ϟ	�SZ��#І���_"�� ��T�X���t�N{�@�A!�e�dnQI�����~���M^�m����XE`n�����	@��m��&L�V���:k�]���
hi�P�������x1�z�ؙ���[!ۣ���coS��T<D~s'�-�hN
��,�&�s�x��Q��x\���4�9Fcc����\i�w�p��Jv����T�����E���{ՉFe�\b�J��`�n�����n~R�Y���$��v��J�K;@�@���z3���8)ƞ���ꪼ�*b�9���|���HC��! ���?�IUK�Q�.j=�
���v�Õ�4 � ��W�3�Q��"�`��O!g	�����[d���Y�����M�>tk��l���kM���C߿7Ò��m������gg���I��o����ƶ>I*زB�X��T�ڿ^�v�Ʀ-d�?#!�����������hl���YT��	d�ha_.�M�,�դ�-�\d�F������=.�%��2%�+*��l}�BR��Ɣ@O����R���aT��EG���:*�_>� l�m�^�	�z1@��/k|�r����)z�l@U�Z��Vb�=d�b|�J��%loXp� �q�����0�\����!�,̌��W�7J@ȃ�i7�,��,xA���ŝ�w0G���Pr�T��)�=YK��{<��5R䅢>�����ʷx��d�/	����X��-:wj�78h���.o��af���)���O�J��P�5��ƾ@�+��/�U���Z��'��N��y�6}����X�p�v1?W�}Џ@�����Y�(��Σ��x��IH�C�؛\:�r��g2�6�3p͍���w�W��!�6)�r)����}����vGKǸ3�M�)�O�Dx��Ūjy���EU��5��cq���ytXǱ[۾/��`X0��g��6�~;m'���-�Wߪ#��/��"���q����V|�~.�d�9]3e�(�?p��9H����G;��:xŧB��t��/"�{���\��\@������D����v0����إ�U�p�w���=��7�)�_��3ؼB���%�������g_�ǖ])�N]��'jΙ�i�r(�]��� �ޤ���R��X��I���o��78B����l���.C@��HK`8��s�=_�gƓ)!�R(�4Uߚ�4�hçR5\ ->���@/D%���f�7̕�����H�pv�� ďau帶M����td_�adF�~��E�[�Vex:
T L���$gX��K��l�X���C����\-α��狰�·
�V_���;Ձ�i��K0��]s���]%Tqrȝ$[ǢkKט���pG���]+��ߜuB��*�ӫQ�����S$�7t��oI	mN?nV���� L���?���@��K���]p��>(�������Ԣ��by#�P~�Dg����Bwq~�>�����b�Ň&�|��Vp2�&	U&Lr)�_��302��|�n�%�	�����������fj8�F��ğ]#��OQ5�Zr��p�8��L���#p��%�%�\V�yDOL��
�Z�S��C5k��2��B�[SW�s�����$k��YNՊ�+�dNo�wj�/ {�����R5����9}�����#O�$f�6�{�7��sU����T_1a^�s�ԛ%wH�ы�K��h�Z���\Aha%^Y����|�1k����9���&O��F_0Êub܋~���atدP�8�������M���<�h'�	U�o���rb�V��[؋�4/I��ާ7����s�9鏱^^� љ��*R�,&�W�S�C"֠�8��a�݁G�������yH���2���,�.q��he�:��t����m����{�pD��cq~�����%����q�m#߆D�>v'��	��-��k�c��Y-���ar��L��6&��%L�A�?�Z���ΔR���o2�*��~�1�%��W�����_Q��M�3�~+.��Q��A���ٚ:;���	vٛ?�vqo͈��C3�85*�ڲ��p�Qp�ھ��e�w5j�E���c/ `ٴ��!fu՟�'a�*mԒm���}�;dѺk:�S�
�-�TH��G����SZf:c(�ګ)2�IwDQ'6�����qwn���{�+�l�ZU& ��62��(�'>ma��#*�K����FˎthT�s����"�k8c�su\9�6� ��F*_�����w��Ɣ��u, )W�{����Ǝ�w5Q�ćj��ڋG�ꆭU<1�r�����S	M��Ao�{�����GZ��g�)JX|��nU=�p���Ѥ��,mԒ�/B����p���J/��/�g�� p�(E?��_�]��0��U�ܔ'���6\�A�������2���~'ms�o:�KLJ��Q�N�9v�:�zD�@/��/��Y�Hݴ\�rU6��5���8ܧ1�ZC1��U8ٶ�'�"ק9��ڸĒ�)����@�	�+�LQ��AuM"�V¦��n_.l���?�A�z�+�-Ο�L��<ſ��cm���F�G���y@#"r�~J�s��r��i&�}��,K ��|#��#SE�j�P�"�x��]�u;����؅��m�B6#���)�S��yQ�l�C�� on�N`��+���R��DU�`j{��ߖCn�4M��8�0$9�V�T�.�
�U�E"��摨e�*�̗*і̟�`�Ll���9��5�u)x��;��mo�1���J��3��y~z :�g�`���i�oq� ��n4yw���L�_EelHD���Mh��7���U�¨��)�V���I`|�U�~� �v}ֈ�����ۊ0�>�K �\��`�z�SQ��c�~����˫��$��B����CfD��"����	�K+�f5W������E�Uh�)p�{:9��'Z��� f&/��߳�V��Uѹ�}���ټ��Şcf��)�!4����ff�"�ݠ|��� U�ޡ���,"%����ʺf0YU|��HvJ�*'�b:�I;^���W�%��!.�IB���J�&G�ɟ��.@~e���A%Ǖ�2��s��	��&�i_]�)q�����rZPb
֮de'�##	܋_sjE5O`xjXR����i6eI�)M��"�k��I���w����<����� /�=��gR�Ap�U��6�x�c�*�&�^�]ևTm% g��KC5��A؆�P���rHl�`�6��+��@.;����	nV�,�S�D�d��[��ך���XQ��U�±�+����HD�f�h}c�:��Ǯҧ��T	(RD(�h�P{9�ʴS�6�5LHt$e�$��ܨ��$�Y���k�f����b�4`��h�M��v�K�U��K<r����;Gb{ [��%�Q���ӽZz���yd��s�x���]��x�A�i���M��H"��8?n3�yֆW%W��H|�Bo:Z{-��CɅ��nS+[�]uOl�w���vF�֪zK8h��T\d�
�}��0_�����KN��&����آs��6�q�w
�v����NM}@kƑ�^I��?n\�[л"���s�S�o��xt}�#��Z	��A�P�'�%8l��;B���5�"��x���w��>���ogg� ұY���rd���܈;��m������5Ȋ	מ.�h�xⓄ�	V������vh�����>ʹ��4��;�!En���T16g�l�S@�5�c� �Ɗ�+g����L�69�S�����¼"U��0�I����k�=\a��Ln/�������Ϗ`2h2;�u����^���gY^����	'`v�6����l�'�]͝����f�ݨ�4���½�ѥI@m}�B��'�������ɳ�����yW�� �3%���Ҵ�4�Sݫ�:9��P	]̋��`&v	2�0C���
6f0��9v���P�cE���o��܉Y`~��g��[t�,��S��iA 
=��d�����v��E���$Z
�i���Q9J�AYl�����Ιf8��D��:G��QJD�x�1j���h��>���YV@P)�]{��d�jk�.�L���7���|��q-��8�e+脙���.ו}p/3@b��.�I�Al�hX�̔G ��h0\2�� ��3�m+k�b����.,SDªL��#2��P��'��pI�B��A�k�����:�1�b� �z�W�h�'�d�68�)�v�R�%�h�����iUkǠ�}�a��&CĺT&��s&7�������[�]�fæ<JXD=�ruC��A�s�R�6�M�: kT2�c�Ղ����{M�s(R�e�%NvҮ=~H������b�@aGK���,�RTY�����1S��t���޿;��'F\�����E2���-!�."A�̌�D̻��0��� ��d.6&Q��F���%�j�g�����k^�(��쾳Ce�wxo�-�!0������bJ��H<kTWfsc{9�5�c��~�~���������H�<��4'��=V�q�'�24�FV@%�����qUc���w� ��>Z�q{�o�ѥ�{]x*�K޶͹�p�3�.�$@�P�I6u��=Īm�Y���&�qH����i_+�,�vP6K�sʯ����'��
�^�>e]��)p[�ˇ�>�'�,��dx[��$���n���I@FV��~(�g�Δ*g=�#T<;���	��PɌ?�7B�i����`妴HF�	��D���>��]�����mX��Xw�y��~)�e�m��k'y��䧉�X�\"��Ǐ�	�>tj(�Hϙ�:�mp�8��.��l�b�8�t�r>����r\Q��9;�CDeS�>������ĩ7�pK*��mR+v�4{���;����]�K�=n�T�,0�RS�����fܵA��"2�B�����EâC�%�Z�U�5�ˊ8�;�:vc�����
�S10��zNL̶9T-&��]٠#a��|��,�p�z�A�^���c�C��C�5��@�&������;T�7Ͻ��ȡ�&�7���{s.\�ϰ����+���D���?�I�=B=�c������J)!$j)���|�~�@��\�����i�ʂ*��eu:��g��++
	�0+�����o���"����H4z�L�c͐�r��L��C�Y�s���+g>B��7�㗜����t�L��z��kп����G������@Ν��ཥ������-y�ҝ��E��_D�G���PᏯ�<~}�љ%r��B6�H{�/I�W�L�cQ'���ב@��w�����q�i���x�?�і��o�_xB=�vH`��$�����i �n�rF���$��-1���T2���=�&WS�ML5��10���,z�en��c(�t��o*� :���$���H��ځ��/�h��[t���Q�kiQ��:dʘa�0�`����1�����(���a#�g�S^ۘCv�ְ�J6�X��{p�h�z�{��t�)��=cL�GOM$�$����I�o[k�-K])F �+��;�d��Җ�A&U�pO�l��*��E$��j���mZc 3����u����HC�doM(I(;�m�c4`�Z��j�?9x0`,����q�l9w#4��a�ʹ�2c\(�N$�5�5v����.��)�@�d��C}е͟����>��m��YPi��Q�2t,f��c6HI�h�昰�J���ź���E��mä=ҝ��Y��"*���~#���X
[T�e�r(i�P@��!� hq��9'���6���%t���M����i���:��#T�Ƨ)��x��zyJz��9�~�;6�t��;F��s��y�z:����{�5.��%��X�t,����p�̄$�W&�at��9@O��%9������|���+(I�}�!ǴL�#J�����H!��	�"���2>��{p�ʬ�ʛ�)v�Yy�9Z�5џ���-K�!yA��T�XC$\V���%f�Ⱦ���Qu��͡��u�X=�o����N�a�$�����E�a�ʟD7���y]������Z�	�?WG��]Ju�m��CJ4e��~ތq/1�,�H�W=׵Y�r�ȍ�y=�?p4�S���� ��D~��wْ��>P_�#AU�C�)�ԭk�ذ���A�����	^y���|� S=�D�)��G;2?P�f�#��>���5�<R���H�%}
"q����S���٨��>3��.J��̼H�gX�7�P(���EbGKc՞�ʴrD��z׃�wpՂ���1e�c@0&�U�����)�"�h{�u�d��b�j~�f�f'4�q�;e�N�x���
�ol������d��IY�؆9�>V��Q*�6�-�X�����@r ����&����v��S�H���� �Y��C(�K���q����.�a�~� �1�^>�A����1�Y��|+&1ײi��D�܆o`��V�uI���1���;�C�}Uؒ{Պˍ��b�Aa���Qaj�s)%�R�����7�81ߊ��=FK��7�m��L=!�u��{t ��a�2�gVɯ�`�繄B�"��ʷ9�T��>9o��h𩦝ǫ�v�HT����o�,���i=�_��+K~%N��ES�������X�bE�����<bd��4Gr%�
�r�S��!cP��Dƒ%�VF�%�?�p�8/�<@��F.ivCQ>�2�>T%��I�Vx���pަ��:\1\P��6lA�^�i�@S����PG��X#)3|�fe��!E;e>�K�O�]ˣ���y���ٵ�+'��{ j�эH�b��fE�K<V�,�>���Z��;�����^{h�˾�1���ǯ��p'�%XY;F .�=䫊��1,��)�X�7cr�Q7�{�L����V��>#�u������
ɻK}W���M�䒾_,��a�3�.4�_�%.aK&$u�`z��LMg��4���0�O����p9���G����K�ۧy��!o6�R'm�{2aViZ���y,!+O-��/�Ŕ�i�	ƕ��Xu]�*��;T��BU�4m�TTM-=:�@<駚�/��re��!��M���5d3�xE]�;~aoΨ��bE4�!)�nUN]]�U�CQ�Ԍ��Q�l7� WNa�sɝ6��%>|��Fx?���S%J��.����{��x����E�;,M�[YN������%$eT
3�<q���ȩXӅ/ud̥c����ENT)�6Ѐ�d	D(!�����\�	�Hʜ8H��F���s����V���N�H���(J9 b�^�B�h6��W~�k���Ф�0=R�R�Hzg��lk>�b� ��n�Fv�;!~���d���NR�sɦ7 "e�t��>{@w�-d���)���NE�;H7���\:+�/�ve�z���0%�����M^P��KD���P��MP�e-�L�:������`IΛ�TB���C�x�I�W����(åB���p"k��V�#+�����eSgitx�)üc�$�J
��Z$��0r0��
���G�����'�ќً�1�h)E_�����⡺�o��K�bM"Ỏ	fT�����=�&-V8��6����,x��S���Ot��ޯ�0���� U��^"�>�'�;<�S���U���m��DĆ���0�R`���U�-��t�X*�)�t���c|̼Mɷ���+�����̱�� ڸ���L�XC����� ��9��-���ޞ0�xc�¹@q�}�����YM��ᎯN��"\�J�Ӌ��n��%`���j�:�'x��cx'Ҏ͟���)AW�#��X��>p������S���oݦ��y3�綁��^wG=�h#���;��}=>�-����jgv�p��g��l���Ķ�Rh��W�5��<>�uMQ"��1ڊX���,����%0)�*8ƭ�(����J�������u��1K�n�4 ᧭e�}�f��0�8�&�l����7��Ҧ�Ƴ@0of?����*T�ܒ?rs{����$ٕ鎩A�ܴ��5��h��]�rꓷ_�W;�McJ�ߔ?� ?~��i��9p�4���X��$'�A������ ���2�Q �� ��a;������6A8L�cG�봿w����c� }(M;�in�$Z�O�Q�������A��IZ�UP��C���$��"�F�>ՊU�l�'�C��/
�z�@M�I���طY?>�	��y?}���.֐����|%�
 K��sĨ�,ar\읷D	g��I]��v�ق�oK8$L���Zݐ��;�R3��1)}
�%�G�x|@�jQ�w��n
����l&"Ҁ��I���/J/��,;v*_L��Yy�R��)��+V����B���9)K����M��1���3;-��>J����+�z:(=k۳Wgd�3m��YI�;C�;0����tm�K&D�S0#�I�`�H
���c����z̀hޏ_F���қ�e���i߭wU�Z��l��n����	�I�Rf��U;hF�Ii���}�<���'�y�f�d#�.��^�9�J�
�	Ώ� N	��������Z�A�����G3�����6��|�|�G��.�ߑ�JZD2�e��8���H�@�Y������o���+Y�/d�Ӯ��,��sܟ),���u���emP��Vv������]�`�*-]~�9ž��
�p��긺����(�'̶H˯Jaw�r�-��dj5j�B��1�U�(�'�Ti?[@���	�P{�s�ĄhB���wW�"����|�I0WU\�����QA����ސf�G�#�'�A��{ڪZvњ�Ș����8����v�0�i?dK@�&��!��^ΊO��a�G�jNϒ'@��p�]��/rN����o�U�W�M� �SK���F�����o��_�V qJ�>*pG��츦����ɱ�����-��vƝ1ҟbM�ZE��}���($`�o�O�ᬺ���xW<n�p�^_bE݃�,`��Vr�tpy_��E����ެ���
Ve9u
�;��R�'ѯ��� �[{V�����L{�A�>�p������:��TT*���v
����*5>U��y���/BtV��ah�h�ґ#���Ǖv�m��E<oR����|�����p�D�8��x�0�:v�`�JPљ
�b�TX�9�j`���SIe/^T�Tjf��EM�j鱕֒r�2��mD-��o����#�g���v�D��Y�.T)Ld4x�I0sxb*��h���"[����*d2�舁ApW(WK�6�~%�/.*���HK���2�4('� *w��ŭȒ�4)H��bxx�d[E�-����=x����sܨ(f��X��%����L���F��ր�����#V Ñ�W�����$cᘱ9�`�\�����8�o�7�ۗ,��牵{�G��t_�{Q��3s7�g�H��Fˬ#�K�K���4�_�H��Tu"�1���Wk���~7�9�Q|$��\3D$\TS�h�"3¤[*�	�͖x���sB��j^�X@��@����d��������:���>��������cB�D$ž���l�Fd�S��� 0ѧgn��������r#��	�}SÝ�}}����x��j�o�{ť;�=��xn����G�����zS��~�V;�EJD�`>N�$�/0�d^&���F�{�
�Q�?�9 h�n��C�2���-�;ޮ��-l���l��T�F�8���Xk�ZN�	�~|ؿ�}q���ř�rL��m����d)�"k����;�Ǒ��.a�ُ�!�#{������sp��:}�TE�2%Q���ĹZ��E������ H�;��T���'b�;q�z��M{R�*w"X�O�o�
vG�o�!l�h�cy����^:H���Β%�Y�1G�ؾ�Í���8YD�����~G�i`�b�r=��@tuAh������^n�G
8C��ٚPN���h��;#J�]f�aO�g���%z����J���h�Z�\Ϸ�������9p?������֮� ���Sv7po���
U0M����[=�o�j���k醽���{Lo#��i��8���`!����kبOj(��d�sS���2m�xHk�T�d�j*�����J@m��ЯD>�#�����R���FU�G�Qk!���Z,������E��6%Z���μ^�f��x���(�yxr����N���I�)2�,�+�h�P�N�@j}�X^B�q�R�8���C�e����a��3�C��<R��
����Rԑ�AKJ�(�T�
v�O)5��^�3��MY��4���R���ݸ�C��⣷D{�a�|�f�e9{�/�X-�οC�+Ș�G����b��!�y�D������❥ UZ>�����s-��2���:�ԅ�F2��vL�bcnQ/ظ��L1N�X���򱦬�6U��Xq���ny���/Bx,��$�����ݮک���(�Re{6� �hoð�9����#\#\��b��^l���u�#{}���x�UR�7�s���H��s.�zΕ�j��u�VZ��z�e��e�����9�������s�sG����z�C"&�T�����z�8��H�۬���`h���K�S���!������6qstx3���ٔ{��f�:��uq�	�-6R,Q���K�2�����r�$��Y�Q+�9d�ܺ͂a\��i�d�d]�;���CI9-��&Av� Kc�4Z���|��I׿#��d�Q�m�2�\�b����OՄ$����E�Zȯ������]�[����������߅Wx�^v�i2���M��9#/�%�����S>Uj��4�'����?y6�3��l�%��\����a(<Ӯ΂��\��:m�Lag��gs����U1V����8i��݆�����]��5��<fX���K9i��u�X<vy'�(x�� Ƕ�<M7��9	���&��:�2f��Q���'<\C�0��]��D:ef���Ht���gD���@��xzBiT�������*����[p�R��'*\�{@f��N&ko����EC���y����h}kX�ׯ�3�x����	
�p����(�������Z؆�};1D�|�^WM�v\��'� i�w9��Kߵ��/B�^b��z��0���i
{8*_`�J��ql�����>�$��R�Q}Yp~r��)Ha3\W��'�o�+/-�]c��[D�#�u=�XN�Q���e�߷�Fl�&,]�8�̖j �y����i��i-����*.ܝ��k����4�!ek6��n͜U����m|���<Ɖ
2.�d�e8�ݜ�A�<9��q@�Ss���k!Z|�0+t<�����k�DqZ*�Gq��ʕ�����3�[yL*�lR��b˟������������JpX�?�U%�xH�!j
c��Ƚ��ϐM�}SK@�� ڹ7�~��!��^AMW	L�k�=���������9��޽T໬0������sX�r��G)�b� ��D@�	+Z�6�_dʸ�����<�#�2�%Thc��񕲤Tͳ�����g\�4��ƙ�s΄ J�n�o���Md��&�A��R�sbs�B��[
�P�����[8FJ����B���'��������/p2e���~�ڰ���9h�ٌe���S�]V��SHD|�_T9$��t*��7���l�74��ǢR����I��`�xC`r1�������#�_B+C�����my�6�/�_}WY���D�#̧)�l�HA���}�n6A��sE%P��L'��oP�V)��y�x�S�s&����\��wO��8[.���{�V4�GM��E�!#��j���GP:�~��s�մ���@7g����Mv�aW�W�^�/��<�e>d��̇�H
<zT�D
M�z�a<����;��Gn@���� v��~�t$��<���t���*�6�a��{���o'��O��>7C�*l�e(Ky���Z�Xm[�G�Bn/;�BY'Ʊ[�N�+ux��BV��"(.ٛf�^Eͦ�B��k��0֥�xO=<�5��EV ���%]�׾	�d�^�?�Ze4��yL?W#�}5
L(��MQ��D�N�Ǫ$5V�e�=�:���ƴ�h��H1*U�0�@I���]1*-Lc���e;;I�к���F �-kJ$6�S�SQ��^���_�ꕟ����Q�4�3.�x�CǤVg�ͱ�|�"����c��ØrK�>_p�kp0��D�;]/�4uH��h?j�6m>����8��kK�O3�������hd�b����6C�y�J��<��\�oAr��\Gۺ+ɮK�Z�t,�Ү��U�AA�N��4]`��m~��"��8+����Ě_�Vˆ�@M�Qfd��lcqD����uz��?��E��s�/�8�`�g��e�-��Nս����9�6��E�����iM�H���3�t�&���Ub�lg3�ˎ��5B�<��!��]Ex�x\�ڤXw�����&��զy����K��n��⍙��9i.�O�%��H�����9�Q��%�b7ᆶJ7��y�|���n�'!m]~�b�m���ʌ�e��f�}���_a�oԒ�;l�_���
��ɻA#!�џ���gH��:-1���o�eb���&H�g�R�*�Pz��z�6|��[���N��]I����8��T����i`�-�x��U,�Z��_� д�%`��e����?�����`�j%�cԶ��+oتʟٍ4(.���6>�i�"]�,��)���BT`\���zG�Ĝ�I�oA�!�C������n�t|:�34���v߬RTc��N���[�c4�E�RBt2�$�p��m�F���?�)��ϼOd�A�"�I7�׎s�4&m���A^T?!����u�H��
������y����qH>����E�r��Nm�HÄ�Z;��x!�2�R ���o��Fv��@�A�w)�%!�2���',�����^fI-g`��?[-!Fp�#7&B�aL��AF��jخ9B��;��q�������6�}�u+T4����E�{Yj�ȭ9�A�e���f�B�u���t�����ۿ�E�ԮG�ڡ��������.�^�S0{�Lη���S�{���L�!�Ǘ�<�/|`	�2U�ڢbڛ�����*H�,#bN�%uYa����\�nUg8Z��AR��� *^�����"7ϷB��T}��̮��۬e����(�L�,�;C� u�EJ ڊ�qCaY��,�n�*�Ps.z%�V�G�����+���&[�%�K���Q��-���׷���Ӗ�P�	��T��`�8��?w�B��a��7})��n��,���V"�	۲�,��f�xH�}͌���u|�k�[X`��

&�E��qvlV��'I������[`L{<5�V�R�e�����@��eN�$��~������4,����,,P)R�|;z�T�^=gpMߐI�~Pھ�pUFdq+���3���a�:^��>%i*� �O��kW��:�S���S0�R9x;L��]�>ϚW�a���߳�P����k�x���W�N]��l�;׏�l��d����DhC��}��eo*���8vmO�Mi�y+��[�x]���o����||R�z�M5ã�������~����
q��1E�5�0qw��f��S����7�b�+��}0�Ո�~��&��[�e�</��O��C�Q3� �Dn �m��5���]�O$ƅ�ȡ��
ɫD�N���� �'K�0%DH�������P0��)z;X����^%���ɬ~5�db�[��#�@�������R��Xϫ;�Zt�S8���|\R�+q��p,~�鱩�hAAwVsrPCl�7>.�`y�y��`4>�ȳ���b�퍼��{s�N�cz�I��t�B�NQ{�\���[���c� �)!��@�\�_�+pk9(�4���j�I���"#�Nqꁄ�|-إ	�n0����CB`'�t�tz�l�'��`"�AW�-�����K�mb��@;���E�:�D���%��)lEC��ޯ��ằW�	�\>��KcY���{lǖ=��m��͈8i�G�Z�bGs7��(vh��D�F��@Q\5�fZ�5ZN�h{z
կ~'�N��L%�ٯF[W�
�-ҿ���"�7��J;��J�Ki^�ޟl�t��Uע�6|������?z�顡*�=ɬ%�g9Ӹk�;��*�b0X9g]�PzaV<���/�o���ݍ��@x����D�jv�+�&\C��+@�ΰ���S�^Y�����^b	.Z�'��0A�����XQo��a��l�˟�å����x:%$.�����mY�6T
p�V~���t�>����0��	[Ceֱ������ΤN�2��5q�v�}��fQ�_�{m��d��=�[WLr�yTmtw%5�]�y�!��c�u���~[A>��vE�p��3��	T���f#��MP�扈����&Ch�&]�8�R1 ����l�j��|�]�r�J�L�\�5ƍ�(���sK�v@a��D}\bu#�[2i�͹�Ұ�%����tna���h�IY=�<Xkl}�/�	L�G]V��g�V�)�;��	�==�$i:{�b>8G��9�Mf/�2n���9]%�:�I�*I@�}%�h�R��@̦U���� �#[g��$�K�]L���W-�Z�����pq�LS	���?y���a�t���D�g��n���4����b�4b�t7�Ei��=��4%7Z	�����E�m�����'D����:�UT��%�$���~���$���������J��ʲ�7,���r�' C���{0>��ld	b��L�@�>����޳���w{�m;yO�$�_/ �!(q*S#.o+p�I7�vt	����>���sd%��-/Hi��(3��e'NG��t��m?8n�I���I���,�����ռY�����2���j����Ҷo0ѩ���8�#:$�,S�uۮ�v�X��ъ��7�Au>�:��C��QS�,s��2Eg�K�j6��f�ӡ�q��H��a&~�Iid�}� 8׵&��Wsn���6epĵZBGW��>C��v�*���g���w|������쎛�t���I�X&w�À{�T
(�`h�|�uD��Τm���|O�/`���s~R*Ƞ7��M�UΘ�lwJ������r�0�7����TT��g#u<@/K::k�Zz\���d�gHP��:��\rc �?L�k�Q��Sz�dv�S����"S�u,���;%������A��K3�GD,)�.ǎ"+�m[)�oeX�#��[���8���t`�~0,S�Q^��§��$w��U����3c���5�c���MJ'���=�JA���#��W]`��#��n'�}j�Ώ^n'�'�MO`��:��Ċ�7Y�p[�J��L���Op���nM	�|H���-�.[A�<�b�{�7��ܟA_tf���=&��	(�.� u� z��E���&ߟ�gޱk��슸,��v��\_mr9a��'�>;��e=�։#��D�y��V?�n�`\�~�m���X��7>e�l�ˣ�"8�����؃��i��~���K����(���D ���'�	kP���3L��mI	�ps���ƝA&�(KQ�~g<��*$�telڂit�<���l�<-�V�z������������^V��u3s��;cj�V��f{
O:i(��-'1Gu�=��٣���=9���nh�b!���]9��vE[���`eg��	��躮[�;��\O}�3En2j�|,~�w�*���78�ڑ��~�� X�cr役����U ^y��G��'%a�1�)I�����n��Z��B�-��B	9q���x�7��S��`"ױ�o�˓T��X��,w����5��dZ�:�h���X�)�A������T�D�b*��TZ�խ&��@F������o_�7����E"��M��q��H	�{﫡�p��S�$�'�g-�W��_�N�� ��r�͏���~�!"���#�y0*L�M�93)Ͱ�k��?�M�ߢ���O�j�Fw���A5�,�t�o�!�
�)L;43�A&)/�nb-y���"��2�V�s��w����3�v�H]2p�L,N�U�r��6Fn������"{�e{-�ª���jU�`� �65[�0�$�N�~" ����꿡�r4���-��ꢅ�<T@8N���d��c*2T�aԪ+��U
~`��'ѡ�g�K���<�u{s\�;)l���E �ΰ7�I��h"ȼ�L�'-ߣ��Dw1������Y��`;� �'<*�@�I_���Aa��a�����hM�� w!�A�=�ԁ�\�Q�7���*e( bűm�K;]V���/�Z�?f�K�Po�cXȉ,Ї�u!\��� ���Uץ4"u��7���y_/��<��孈	�<�VgR�!��"�]���}�Dj'�ϖW���b�:�#V�?y6�>�$GÿlKq�8y�_i5:���Esغ@���`L���9R�h�%�)�}c
���;h�8ou����*د�\̩3�ifx:��7�vڹf�03ԛ>]D����0<x�Zm�ؚ]��dZ3����C���f��1t諮��zP��}v��O�p[jC�k��G��E8+M <��A�ZO#ڳ�b&��.�~N 2&v��;�]�v�˺�4Db���<���lg�N�9��}����4x�`�2$[����b�^��pJE����:�q��g4�P�Zǥd��&s�^wa'�K;��i��3x�*O+rcqf|�ة������~�����dOU��B�7[+zm��W?QU��]P�Z�����o��v�`�M�ce&�×������@`��)c)�Gtؒ/����ݖ8[,	���}z2�P`���[��)\��I�~Ⱦ�яH�5�I'�́7�d2�r�[�~��&���=Dº���4��m��F��-/��E��~�{X�,&Q6MiW��Ʊ٫�Nk�����C��rz�Wn�#`����mW(�4�?�x�<��l��������G�=���M#6����-�J�S-�2��'�Q������:H��N'�_��I��7�^�M�m�F+uVT����=Z��,�|�b�ϰ#�D���?�=�p-�ص�*Vh�5XQ�S��E�V�`��i՗��ނaIՔÄSo��e:D�L�!OD�W.k��"����UQ˿��YB@���jFyƠ���$�{�7����!�O�JFv������l��"�G���N��gTO]@E�tv�7[ܖ���l�m��E-yҶX��7�b
OS%
��Ue�i��h���(�UJ�O9nW�A�F�E.�؛�ĵYh6:�03ꢯ圗O��~aP�O`Rw�+a^+t�3"�|ٮ3ޤC�4Z�2��A--����"�Y���5���S���a��J�;�KM`|LF��$�����px{C#[�C��n'���%0�̖9��	(VX�v�p��ו�>%�{6
�7�C���7*�|�[������%j��d  �Z��g�,
������%��"&BP
�y�4���`�d�O���֊�Q�����-;6���dge �K3]��8��@�-�/v[�J�wF�6����Qa0��gh�����A�M�i.bgeSH�$��1v �=��]?��"�'��u�*�5��0����������靔���n�����-�p#L��^Z�}	;Tf��,תּҶ�����`t�c���=��� �3(�H��Z����32��D������F��6�.*��������k�ы�*�i4�m�?H�>F��6N+��.~�ߺ����e=��&k���꛹!�c�N�� Ż�[�:n.w��l��g��Zʬ��G2��#CT��s=��<s��W�"/L�8o5�")���Φ=4���
MqWb��(6�]Wa3��[`{�~��3���ZL��uj2�w;�@��{��X����7F���I���BL�5�j�8C�I�%z�<u��NUS�::ReHn��mcY�<&�2�(~��I�!kq��E֎�������;AU���C��q�QW�_F�m�tu&�����Kڕ�BG]G��J[��$�;i|Ƿ>�z&y<H�֟Qv*G�'�J�Gy� ����oܐ#u!�Ӳw!�G&Q�0[�x4���پ4Qq�ʵ�'Z�m�����|R�Q��]��Ϝ�g��s�T���;E���Dؒ������e��/�IİEuE��Cv� ��@�YN��҅,�0j_�Ϊ��^s�mk�\�� �� ���ڨ�&��X�*=뽼rN����=Jzq��+�/�S��<٪ɰ�I*/ި�zA�u������z��{�D�9��2���̠���6w���J?6�*� 0�D$��߿!����^BfCfpf"Qf�ͺ6���mEr��ؠ�1|yV�p�N���Y�Sk���v �D*&����:Ą�QǴyK͎�%��"rX�>zWV�����������7���צ��_�{�!c��Ѫ�T�u�VT��F"��C�P�<#�#�����fsoq.���`T`�'Ǽ#���V�]�=k%�"s�^s��K��6��>�<M��@#���:�ԏ$��M�����:�<^���6����U��i�(f�d�'�W�pvS'o?��c�n�}6��i6��Js���:�ϐ����h�|����f��x�~VҙM���^�$o��q�'(�O���z_<���M*@��v�-���a2�Aw�yKq�6J�P+4��P2ꅸղ{�	]���֒n�yy4��8�=�2��i�(��x��`� nԳ޷��j���-�!)L��V��@5 Z�i�C:�Q�n��
7=�G��&ݢ^g�*^ZD��Q�T���¸(� ��U��OUS����&R�a�]�Toh�A�)��h�\P���}S2=���-�{��䇌1��]�LF)�����l,b�IU�$�XT�(u�9Ĵ7SK8�/m�UR����堡Y��p��UA�������Z����jh)����yF��k��~�@�0.X%���Bp���l�*�	{t��.�Mּ������b�KM9N���9z��i�';�;t1�{Ah���{�rt�XD���h�_*A������C��8����NDK�K<�D��7��UG_A�����l�O�=�|�<W�p!mS�?.�P?�'��^��`#��o�^^�'�O��&�n��>��OMJ5j:|�t��W:*����Y���ލ����A��BR��V̇�`G�띩UE�q�u�,�z��KV`�y�{\$��	U���G��m�\��J���'g
h닻i�e����>vg";cD���KǙD�|�놑OMކ̉Lo6�)�k��^(�^��u[檊B�]�E��1a�:��kj�x��q�"~v�~��Җ�+�W�;��n$7�}��.i������aq��"�M�X[I~S�g5�{���� ��Z�d"ـi{�.��#8h: ��#�e�3z�L����������'I�pU���ڇ٠�Q���O>��XG�9�$a=r$� YIO��Y
��Z�'�= ͩ��;w��!v��u�$.[���=.�]A�H7�������D��>���?�������x�C="
���Hs�q	�:[SS����k/���@��/����]5��)@t�O��ڦ�aXZ����'@"��i4Mf�,����(�󛧦���	=^Qk	w�K�?g�����S��u�+|XC1^PQއw�i��/��bc�X���O���O?(��%�5�2S?A��A=��2�V���ж��(�<[f�M��$`v�4������|�6���^V���W�F0�w������Z<�d�F m����Ψ�[*O����zn�x�@���\4����!��:ⶠ@�� �]��3I�8�a��pGU�S&E}������ �ṣ}y�V'�k.�7��� �	��#��2���M6iP8���'�X����_�]Qv�⃟j��B����jWª���R-hn�,4������pY�ُT�h��*S��ׅ�A[ĥ�豬qF��U��w�����ͩz̚�������9������	vؘL�&&�3�6�.V�^)T��w�Oj��E�=���5s��vx����yW�|��kY���PF"Ƣ��<La��7el9@u��.��-v��C���S[aZ���a��!6@�9�q��=:�g�=���������O��f�dr�
$b�"�/8<Ղ�RK�	�-���m�w�i'��*wš�L��[�y���Lr��m[ܸ͛~�(T�1���@�InL�P��9 ��j*�����:k9���FS��MJ�"����R��T)��n�컇��b��o W�r� P>�<�eq��ח��7Xs�+���E����Mz�fpX\��<bt�SՏ5b�O��iQ��mI���9�]����ñ\j�����֎ĉ\��v_U�|���G�-�	K��� �o�v��b��A�����a
�_��4��X���E�[J%"�4��BC���n���ɢ�;+,��\k&�\1ހ1�F7��6v��+���UWhN�/���2�>h��\����XG�&�ѫ�P��i��=�O˵�K������h$Ӫ����Q�~�@)� p')�(�4�����{<��q`�Փ�х��2�����7n�q0�����q�ʵA_q�⎰�+~k$��p��hiI�����Y~�b���#nJ{o�[^qܒ��+����7�%r
!�:���{^�#�W�w-e#���^F<��r�E�9��v���s �#������M�d��NY6�~򇊊c�R��"Z~�_s|�/w�?��G��8b��݊�����x����~v�Q��x�B3ٍ���j'�+h��n`�K#���M1rv�*�b�ͼ�ϴ���殫�d��X����C�A$i��$�+�ߖ����+Q�㔎��b$U��d�{��ϋ%mxqൡ���g<�C�7{�%i�f�OP�{�wvXm��;��I��Q�6=���0��hLZI��(� t�RpT?���JE��E�:�����u����(�8�F�������x�u�oq��&N^}6�7�SV4���8��������w�k��sl]9�����5� 9��������UbZnMB�E`���c�d����h\O��`��)|��{d�'�!��Ʃ!-b�n�G��ti��l7��T�1;mE��U)��dA���``3f�=)�q<��n�G����R��k¥�ǐa��������HU�az)X���Å�)Qynqw��Z�M/�!XXv��R�$��{8��I�ٷ�� ��	�*��`�}�O�V2���|��q���W��9]X�ʤ�+f�lqZ��Ã,��U<�ոI���e����I]���P(�mL��	���߸�o��1���˞�?ʎ�S��ʐo� �tn�
��o�fA~��?�Шnb3���ͿvI���fB:���A�ƂN�<S�KQf�z�z�,�gg�������d�	q��:?�����x�j����&vrJ�&�������_Νv&���]�^Ԋ�/��
�@��#�����(Ȼ@?�!��
��?����i�hҒ��=� ���x�Z�״9z7BE���GrC��7�  H��!�d�B�:����p�y��6�̨��o�x�x}`ţwP̸�>	��M`̬+�s��6c{ V�^���;�*k}�A�2/W�� W�K�`M�a������]:�I���7�'���0� e+�]:夥�������Bo[�0�0�!JEj"�L������!یr��t�r���o��>��r��G��Ιq:�Ks��.����;��ۻ7�g��0�g.��F��9�C`N:g)�5>>#G��R t;�g0�9�%��}~�Z݇�����ٹÖ�a���Ff:�~�L�e]F�8��o���mx �IԂR7`N���ԕ:b��T�}���Ws�A$K�N��)Xv�_��>.v+Y�����QL�R-ҁ
��q�T��|DBK��u�k�1{_#�y����>ƹ'̉�Y%]y�i�Ѽ�rH�G��>���!�b����O�y�����3���>{:���
�ۂu��^wJ���	? ґ*"��Z�(\*��x��:\�|vRO�b�w�ti�rU��fIĉ��t"U�?��4	� 4pϢ��*�O��1{�߷�48:�B�a���awK��|hq��a��1���)J���k��ָ�y���G*3�A������l��_)�#�α��H[D�{���%�Ԭا�i&I����Dc"����k�O/����W�َ�������@�A�2�*�"��$�6������ĝ�^k�	
���r]�w<�?�׏�4,�[F`��O6��΃f,�&E>;���Q���a	(�
\����y�򩥼�{�4�ɀ�D	��u��\ǶA"-\F>Q�L02��	Ks��ݷ�'�F���c��^��IL�	��L>��D��ǥ�+���3c*�?�ED�$-?ݦ�~.,��K +�?sr�˱,1k����H/�K�"��"m�k���0��E�L�����B���+�)�he+�I�.�;�p��'��+�����+}�ȷM�3�(����5�I���uջ���-�(J�%����b3�N��������=�;������z�e.�����	�Ȑw8��6Ҁ݄�9���6GB����7f&�-u�׹S
���|_�Z��X-�~��AJ���"���a�U;��l�-""�ƺ)��>2�X	�MY��J�����L�)�:�8��ae����շ�GGA�����kF	�0�R��8V�8�fP=GH\⽄w8,v�\�����!*D��E� ��Za�>ED�!���k����/Y 1a�)�8Lk��S�����&�Nb�mG�/Jp�z+x9v���wel��5e��De�s��]U�~q�v<�S�|��S�X��Q|_��L���>p9ի�F�O�z��B�"ײ b�~=���iϜ��KʤXg��<�ДS���U�:����00�Z��)��DU�^A�6j�Q�ń/Ǐ��\�i�7}I~�H`����O�k�7�~�v�Ǩ���o�z9Ob1M�̸��������F�ǔ5.���T5�Qd�Em�֎jG*�T�/D���SW��$8�`�3���9�}G/XL@��:�L;F�-����,�/��|<�*�*s
'��"���J)n�o�^���$�Y��;�3'Bn���ႋ���TPYM�x�D
>�4� �y6��/K
�T����R�������@$i��1��q�)OS�S����?�Q��؇�8V�e`9}��7�>�	s.��p�,��N�.��V;i}�#wzL�m�vl$�����̳%�F��n�����p�J �i@Ɗ��3��Ef�M����ZwN+���+��Ž5 ����/h#?��Aa�8.E^<Y����	إ:�:�fW�.D�i��դ��>As�`y���D!E�\��p���h��TFޏ�U�1J҂�ao���4�vr[���-�=���}'J�48,��yx���8�&�L�=gbb�/xa�;�i!^̷'�T��j��ҕį�D��3�+��a���m����h��V��V8��1Iw�G�$�W;�
�Y o<�߇�.8X�z)l|
���4 �Τ��6	�`y^�~w�C�=����G&�u�]�+r�ƿ�m�k���;;��m��ʢ|i�� ���;X�?D���:��)A@"/6ݷ�=Z	��l�4�H���a�*�E��0�������j�� ��	z�z�Flj��r<vAx²�"X؉��aQ/%�Aϟ!UwO������qU�U�8��D��#_>�Į
?e���(���Z����4�#I���QIL�s����$Pe���u���j��z�a��Q�S �2���c�&��B�j9��+�Fҹ�Y������l���1q�ӕ�(���0md���E�KC8�{B�=��/�imO�ryJ�b!�gct�q�S�
� ��ٚ/q#u.*z��l�;��*A�1��2���Yց%���l��L��An �Bqj�A� >�Á�g�>��m�-��υ����NT���*�����W����q�g5/>��lP�ݿs�'�٩���2��_�ƪ�(nՄ�����W�YUs���-yW�MD&4�o_L�V*��r�[�����^��P6��5r�x1P��}*�=#o�G�5SMy%T��>s��8�+�x���$���21���$sd�3L�Y8���?,*���eb��&�s�
@	q��}��byz�E��V����Q�<�����-� v����I|�6�|���<O�<�P
k`�Yh�-<��Xv��-	+�*�/��3��U�tB�b.���5!���g��i'T846��-���XB���X4��b�f��F#枮kmup�B?C�tx�t�
�C��q�;�'����Q/F�'r��A_����Psأg\ƹ�5��'W��VJ��F���*��B)���"��]7������Ť��X4Z�ǫ�×��*2������|%�`�K�$�Td&�m@�gC�G����s(�L�b�4��Vz��h*�O�	��n���(f	�T�Q�t6ȁJc"��5��7VwA	I���Y�	2����5����1��E�~_�e�p{��b�ROj2�)�y�L�-Y/Q���YθOͲ��ztq�3
-��"��ݾ_�@Dl̿5-��~�:�0bbo����&Pd
G�Xvi��r��o�ru����R>o"�^��0t���wU��D
}�1�����eo�2���=��Fh���@���_m�1q�J�]�2�;�Ǳ�����%`�4�dZ[Ӯ���{@)`׳�RWJ�i}}���I���?�@ɣ��ŗX�)@�c�⪨��mMAH�P*p��1>��#��B���2x�q�����~�����=�g��]?����8�?���e1.N�,�H{��g�ڛ��
>�ߔ��rO)��z��4*��l��m�$y�u%㪒~��!�9!9���5Z/���2t��M,�B7ә`�黌@�GϺ;@��j|*�������J��)_�S�ģ��(�:g`r��B��A����{STR�c�!�C��pg�Z旸?Q��Zٸ�W[���$��8�|�l�[�6+	�`��hJIn�'����C��|U�<�~��(����������IJ&�����S�|	��k���O�d����Ǔ���v3e�t�>#�ު|�5��3�V���S�HB]S��%q���L笽�>�^/DŞb�?q���R<����E��0V���6�p�o�e"����Z��3җ����
���U^�flG��C�؆��������v���&�/�o���ZM�7���/��d�9K���c�`��d�D;i��$��H2�����HJ��׮��M�M2t����5A��|�H��k�|{��z㭤�ܴ�u@����묃I;'��g���LiE�K��N��!e8�%N-'&̝��)k�d�Xjǲ���n�$��g��4��ꉥ�rk��Rf�f�M5��;ŝ�6�/����5?9IY%ˤ�uHQ.}���)����I�Nw���Nc�L��B�U,��0�r`���0]�A#B�I~F��\1)2��XA@��zm4�7����hbta*ډ �Y(Jtg�����50�c|�m>�/'�_�dy0U��5\�jh6-Be&�� [`����>�N�)��3���I1�@6� �O���.�[L��r��}�R�/�(�}�| ̨���nb���a|���������xh[���l�O�b$�Ӎ<�E�P̾��Y��:�
 wRtI���mD�_B/�i��8��::��H7cf��w�:y�y�����si�W{2;�R (�����^����Z.9|��Q7kvІ8E���g&H�*�c��A�OOu����[>ʊ�G��bh�T*ҕ��E��%����Y���ev0	�qZ�Έ$C:�)`��g>�&$�q踣z|�hzD�S(g+�Ob�c�}�3���Y�	��XΫ�V�֩[¯2��2>���`��up�o�28�
LgF����}���TZ]�])?����$ё<���f����tobG8�~{��UK8��B1�ou��9zD3�ԡ��Ɇ�Igv�����ӯ�]�|˫�k|Z�"D���,��.�QV@��������w6��#�W��<�k�L��!�ʉoo�jiօi�����hU���<�D)���HG�_iHZ۾�q�IG�ƚ�a�Z���ϒ��g
�>9PC�K�y	nq��S/ɈYv���5�����Y��M��^�l�<�:+H8�A�����d�;�����5��Գ��x�`����Z�LD���.�f%M!��̽I֜��e�&!o�Os�at���]4r�o5��X��xZ>�T1��wk�Z��B��B	�>������^Z����a�y�,�s:+�N	��i��(�w�)��y�>u$	�RA�T8s����U����͕K�ds~��PSr,�z'Q�aH ��֓�F��h�Q6��lB�d-ҏp"d\M��툭��5 Jռ,���N:i���Nǜ§�6b���֝@Wkc9��k`*����6��D{�9 ����gm��k���M�k��p��"'s\̌f`k�L_�2>�P��X�b�#[dfU�ާI�"����S�%��F��Ø�f�0�R��� ��x���FW|H �l�(��HLx�9/�~.'SC���
��'��{�N
esCP�z+��Lĵ�Zl�e�A����1�Mh���G[9b�j�M��z�i��~�_�:��S��tWY���`��͛�_�	��Us�C�@*�6�bg&;c@?)�'�t5�7ȓ�����.����q���&Q�]���^�Bh+3���i9������ ���ӻ�\|� U���Zѡ���{^(�x����/�z)���}4��%�]c��h~����"�6{6���W��D{��$�N �iYA���'6�Fqi��L������gt�}�6���Ќ�S]#��*�ռ{q��KFo�t�yyQ�-1O��hc�#g�HӇ���r��S��|W��Xf�&Mq�,���F��lvՓ��f/�1O�6����2�AmP(�&���ޢ[�¥�q��>g����GM� �vK��g*� �Ui���Kw��e�Rl��ܡy+c�ߧ%�6Ǻ^ctm���y�Wض�w����h�A .�0�l�N��>� xk�B���ƅ�\�
J3�6���ߚ*�,��E�y�JߠZ�e�$0ϙBw�4�FZ;�fBH��ۅF��;#��n�4��^�6ؖ��	'�&rV+�vJ��i��v��dg�L��8��Y�	��]�(f��D�,�����&{ܼ$��]Z�p5O����o�Zu���L_]	��{D^��F��mՕC%��,����h���k=�Ϭ�!�2��6����!�+�/m�uG�����1L����25՚K��d"|6!'��=7B�|��E[�����l�F��=�h��q�,������G5�������{D�:��hGg������*G�4�B�b�-#rA�h�B��<��ȿ��ΘzPl�	��,��{����Q�}Y�.�%ἷ����՗;)b��&˺ ��p	?�N�$�����;�}x{F�B�Y������Ik���QC� ��ƺZ}��W^���EOC$`���m#P�n[��������i�"�5:bU�����h������Z��Ke��ȯ'Jg��9	2���=w�k�r�5$�7�^�#��R��
-�A/�=dYW�|����+P!NB�@�u�Y���h�ݵ�A�� ۵�\���Q*���h�`�_��`êv�8��� po�t7:o�f�1�5Cz�%K\]}�e�1�z�(��M~�µ�
`�[��>n��\<�f�I��+�Iڑq��+���y���;0|�9���a���J�q|��G���xl9��9�y������lĻ�w� Z/��J���mu�Mb��]wGL~����2ݽ@H�J�=�Jeʽ���,Ӆ�	��ɓ�97�H��yU�Z㐌�^U���p�2��������wTd�1b޿�,o0��toXu�lak\����E�:�,޳�
�#�i:t��*�oH-�I�ɔ��P��a����wr�l�Ǧ7
�cM�S��H OM؏S)ceU�I����x�+!%���%j�'ʃU��; ^*�'з�����j&����2U�(�Bf)���\9E��7�>,2���ЭcUA3�ST�¼5~g��%\�#D�Q��5�S	�=J�o^ԁ8J~�Y�h` �;���r�������d�����Qr�؆Wځ�W����*�iP�!�p=��� ��%Dg�A��'z���4�=��C4R�7�\;���Ts	����h3�{�� ���pi%��%�G�	��J6ƛ�}=Tj���g��8F5���"���V�k��D0o墝+-[� �Yl�����H,[��ȝ��w��t��L=�e�xt�5q݃���s��D\��FQ���(C	B"���`:m]x�����T�����������c�|�^k�)������G�v㖀.)bw��\+8����3��"Q��Pj�(��-�m���%�
��#�r𥷍�[�x�s�>�f�x��q�[\��iS+G
�7� P>U�+�*��xElMY��
:=�\���t�C�K�f�Ң�7�^\�֤�Ob�}����3�h��>ִ�x�x05q�!h-���������s�* ��0]V�9s���S�XX	�YrK���4y�\�Q}�=��W0d�����o�_��ҁ���UuA��>�_DoTEN��:����V]�R�M	r+.���s%�$�sm�B@ٕ]b�zp�P_��0�O8����#V<���O<]s���˩�)f��%N�?��q��N��/�q|J��g�ڃ�󊆓}f�w0�0&Yl��'XL*�E5�	kz����Yk[4m��g;�L��SI=��s��i�`������:�Ns�J�V��^䫁�V�B<Q}F�" I�]8�w�ڍV����~hQb.����d���S���X��.��2a�u�7��룯Aa����V��RVy�3�҅����R,����tE�\dzA5�҉�n�!�:��G����Oy>R-�j�A������сuLgZ�T����ݓ"l�� ��g�o�{������$��Ξ�_�n\�/ � ��>�Es6�%ZN<N���J�&�k�+[#�m@���]����[[��a�"�j�m�Ժ�D�E�~�H��ٶ���<��_HP�'�!\���:?8�����a �p��m�wRs����l�h�¦��alh�r7=M�7ғ�93�B������Ƒ?��!�.J�I'.��!��6$E�Aăf<��!�2}f�����Xh[T.��0�m�G��K���,f�ė�����ax�¶ܡ�β�c3��)5�	�1����ji]:���}çٸ*��sB��3b1���O��&�:�A��*��7N�6(��j��r尹�l\�׆Y^�q�I�\�H���J�d"{��&n_��'D�$��+.�e"����rCZF�{�"p˞�������-\���BI����m_�1
Q�� y^�5���_C���
�w�#X]#!߽5:��丏Dˬ�/��yaPd'�z��	�pjKu���]G��Ӓ�ٴLM�0[֔�~���oڵ<�ʗ,���XN�u��$��\S�SE֍6(���m�Dw%�5@)+��%���/W��Z�Nm�A#OT���!�o�.���E�����Nŭo1��v"�o�[�jwC��|'��Q�����09�y��k��z���m?�P�X
u�'3w�~D�>2�>6�)��វ���!V��T���X�Q,�҂GK�����+Z�?��k�������d���{�'��6*�Z��X��L@�j}��t���W>8��I�v� ��|A�fj��CM�ZW��e�FJU��E�_�B`ܫ_ �#ܴ�(����OT����m�q>���O�� �5�`��ɏ$��;�-x+p�'T��>X,����׿��@G�i�Ԭ�ol�<FM����h��rKmL)tƜ����C�ex3�vyi�����d��o^"����WJÏT�̹��T��T�鿍M͝���!�]���l���
��6j����;�Y��w\R(��w�ZFj��C:q�ǐï��)�/S�sA�,�;�`9�U�Z�p���;�i,���ٟ�/γ�1�u/X�Y��;Wh��IF>�� j�?�𩊈Bi1-F귕mn'Y��f�^�h�
ka:�������Fw�-�]�q���r�}h!���v�{'.�v��2xhK�����u�>h��ژo���T�ˋ�+�g�ش�Ωi�z*<�J���*%�ʺB��ߛ��%`�9�[�,|Z@�<a�� ��yJ��`i�\�0hA�Z�b��/�L?�;�\+Ɨޱ�(7U�%h�5D��E����l9eX
*K�T��c!���^Z�O��z����r���m��B�v�=�>�G!1���I�H
� �c���#���ڹ������:��R��8��)��?�a]����Z�2��6���i�4d<�8F����h��a�b9A_�׆XZd��DA|�p#������Er�n*z�U4	*��yeI@��t�����(~�������*���R����7���k�H�}@�][��Q���k���-z���n��
��}z
�e��鶱�!�+�l�C�� ��3�/6�8嚭{r�^`��5���C��x����`�
8\00tӎ���d@�ןK��Q/�A����m":�!��Qz"��)�n3HqV�d��Y67��I����{��Q(��7���ʥ��(��u<u�B��2���i]����O�XŹQXе�C��0��Xӳ[�)<]#�M�%��i�8{NS	94f� ���e�9���]��L?Ҏ
2��)oH�| �D�,�����4�D�y}�m�!8��?�n�9�v6%醋0�C�{�����d�^䆊�����[�y �a�V���)!l4��`@-�^�¢9�v!
o V�Y���(�+.�8�ޗ�2����k���=Y�Z�  m���ĸ�h���G+T�gEݗ���w��'sߌ�F,�П'��X����P�� �3$��vmU�@8%�`�J?)V���nST�SVWT�;R�)��C�_��R֊�!������<��|�̼O[߮���j�56��^_ʞ3ŏu��k-����;�o?�KI&�@�>m..�=0����[�ht�9?yE%�4�l�UV��F�yŪ*H��^;n&�qp�"'b���"�W�@������'��ofN�|��N�g��r�P#E���4�y�����d�	)@�dv��h&5Z��IF��Fr�ŧ���gY�J�x��6OL�t�Kު�	z���:�U�����G���y��Bd<�.�����  Zn��������]�)�x�'.ن�.�$Cs�4�g���]Z�_�.X_� � ��7cm��h�>ք(�3�21CCf�����
nG0/�_B�>�g���Lk��'������ׂ�|p�gJb�Z���y|Cu���jy��j�k��$��L�_G��)rzf��Cq���,B��u��[av�q����3L��0��3%a��r@�]g��{�� v���#���"��ETX�L~ť�d��]����f�i(S%Ağ��F7E��n��p�2OcZ�Y⸑z�$����}#Rr��D��Ti�X��j���&ʔ�����	(cӔ��"z x�i�]���&���r�]!���?jcb�."�"Q@��⢴N3��_�&3��K]nFA�ߊ+}#D�\4(���Gpy�^�u�B��>#ބ�y,�n�g?���~Mj���ןWue}��N��/o�Fo�(��鐿܄:���(TZ�1�N�L۾A����tZ}�t���=��j˭�Nە�?������m��dZ�2�x�!�w|'%���'u��.�þ1ǅA�y���ǲ�2]n�J�yT?�W�דD�ӭ^Ѽ�-�
�l��d��6�h�,$=8���Su�,1�ظ�~����+�~cvf���$.2��Xi�����sx������4dn4 !Vj�VT���qJl�|�"�L���2��	��C��ű7HP�uT�K%瑓�W�)���c���J��XL�N�p���H$�醀�Y��\��X��XX�9�ސXJq(';�"�����`!�Tu,�4r��*J�� ~��C� ���ao>�a��Q'fr�bv�O�Ǯ��(}������[bbeH}��DƵ��b�yQ���|'����]��"���A�{W���ʴB�z��;�Kӱ#��*x��Bۺi����Էl�ֶ��>�53I��@�J�M��;�P��߈O����J<_Qb���#�����M8���pG@�K_E'�|z+q� �������p�-�s~�TK�0�A�,B��l�A���_�gq���OY�u�atW����Ό��m�0�
���I=��s6�� #��~��a�(�4�ޏ!�~�Fl+㜯�n�	�˽���j��Y��Av"p�+�QG(~C��C�����f�F�}��z��C�;3h�򽦫4��Ο���3H�@򂮶I��:g���������(�N�D>Ԍ#��욣~-��h��ʆ��iH����=?{��l4�Z�W���'O<(aZ��3�W����{p�D����|�����I3pS�6]K��
=r�I?�RJ7�0uTj�Ȉ�}3{n#rb�p��Mеb�e�������=2�䐾�&SKB= �K��8i6�|
|��&��dI8
�@�5�v`an�T9�>a,v��?�K��㪲:1�[��
��\��%�����K7@���Ȑ�+}�FΎ�u~P�W�12	%I���v�h�Q�����eHѫ`�M3<QG�v�QU�=G����\3�#;o������R�lmƯ���5�F�E�)����2MCk�U�-X�8��
zxfS�C��H<�G�	`C��P�K�(@˙��kW3�A���@5���W��s�-��o�'܃��P�-��Z�Hq(����0Z��Cߎ��G/�������q�ҙ��Ͱ�fg�Wȓ%f&4%�#@�Xf�}�!���V�&�e��V޽Z/��m��ַH'I2��l�tE��L�<� �B�%�%&˭f��  ����m���T���� �jj����^�b�@pI6q/w�E9�� (R���4�||4�ҿ�r5�a�ű�}T�|F/��|ѩE�;�r[���Ǖ��Y�_QɁ�^D�;��k��G�ƫq�k8�[����V�U�/Ӹ�/�$DZ�B�vZ����sC��bj��Hh.$�i�D��/�bW&SH����7kV	�B���=��3���T�JA�ǺK��H�|d�|u�Ǘe�h�? ��X��g+Ԩ�\B������g�#�'��PC03u��<v?��J'��D�WS�W ��� �������g��$�+�	�5�/
<X}_�x}�Ri^���6�@hk$�k����c^���V�ڏ��d����4�Y$���;�~��CWaS��qXqO_L�ub��g���p��ɼ�Ȅf~JP� �w8�{A�������x����d����T&��������h�^P�%��605�an�036�α>�J�@���36�l�0U8��*�x�:>"���ŷ_m��[ߊ?!9���C��Fb|�>���8׎���<����V������u�>�%7;��Zׅ��;4�ZrU�M�it���Y,�4U9{����:9G��� �L�W�_W©�+�,S���AP�Ios1���P��M�~����*�cS���𺐰�j͂] ��9��i�L����!�u>��@��6Ե�/�pۃW�3��Z�޿�������-p+�4�C���~�+�����殉S�+o�b�<��v��Ұ�Io����ۊY��;p�G{a���^ɧ�a�HH��+��b���p��^�!�{h�����y"�(����6��nT�.�?�k�׹��{�՗ғ�1E;�j~��|�b�y>���ﻃ���̓����*�g.Uy�,n�-ƌ@�^�́xI���õ��a[�y�M���&�N�w^'-*<���[�h�;Zyܱ��]�0 -��%��E���{��w�2c�B�:��F�=}�Y�K_�d�#B���n?b��WcINFu�L�j�i�Y<�퓉�i�*E��Е3�+m��&��-]�����L*!�Z��s�[��~��~~s�9�� �ʁD�+��e���Z�z��&ǯ��T'���9�1��X��o�3ؓ��Z[��=�l���Ήt0����9��ૂ�	�o	=�l�݋jr��/��*s)���oV%���f�~��/�
2V�~�3�y�BY�L�P�kx/Rf��/-T_5��x���!�
�qM�!�py��Di�Q��W9�w�lv��I�K�h��Ow#*�K�eId�nPxbT�����	btn���u� 4[�6x;��jWڵEa�եhh�7_z:9/d�I��Ȯ�u16d�@d�ۆ��G�]�.[��Ԫ��h/YI�Y���B�u���M�]<	9V&����?����!Lº�C,9w�l���ņ`��1<dߗ�.`�#�n����`4i1>J�5| K湈 cњ�!��cnu嬕��X���W�8"?��G�z����(6�1�V��� W�<��xo�*����e�����-�m���`1u���g87�2,��T�-)���F�,�?�<�W2����T��A�.�-&��XtYQl�3'Ow���r�X�1P�p�>�P.�R��Lf>�_�� ��Ҏ��h1b���[�̺p��0tz���q}�(D��8������|V��ZI�]����?f"�m�vN}��F�c@��wE��%(�d̨��f��a�V����JR8�� ��㙀�%��3�ݰ�ӄ�����7�x��GN��mX�y&M�l}���g�=1=���O�/��t5�T���_
�B�v�K�a���]�UɬA�3b�#�p���+�t�QmN���8's�e�[��ԅd�R �"�)�G��w�?Pne9�_@ƘL�A|�8���;J,7U"[o:c_���Ȇl&K�$t�7�k ��L���K>�������F�%�CC$��������DC�>+��a'���,�aO5�Ǉ���bď�T�ᥝ�aޠ��p/3V9�_*�=/�!��]��Çzg�G��6b5�W�%7���{`��_T�]rM�S"+k�[�C�>��M��p�lzkP,;2����2��LG�`�ţ)A�+�4�̇-���}E��������#��!�Hs�܅� ���x��8�K�C��g�#���(��.�<6�$�_R"3�e!����i��y�i�M��3���28�I �7Xi�0��dd��\�M�!$Sg9d��o�v���:�ٻ�-�=R<��e��5^�g;�K�w�3|�-!%��__��|��˳����j	Z��_��A�XR��>�E��BI����<���$��Tqn�w7�c����A1�'�?(:f��BH�*؊���j��.�3o�0tzA�:56�9:���=����T�.@�����6#N&l�1�JF3��=}SR4���@�P��0�qY��j�ϙG���mC�l�����.�KA��N�V��G������#�Uޢ&Ơ�g3��ShvG@d��C����bN���E�hK��IAփ��Gq�L�������]N��|�`��HY���Ћg�y�d<"�Zw����׎��4#c�ԣ���/����p;����Eb�qV��Vv��������ʠL`B��C�X��s�/���#� �5��x)p�~4�Q�(pZ >AVN'��ã�9��&\��ML�}��!��{���-�)�ً*g.Aj<a8�eL�)a�������U��*�<���G�9���s��R������)x��f��k�����U��P�h���/p#-��L��\�"�9�w��h�[O�P���+���+�T�� <���x�@�R\Y�g�r)iGe���~ً�(��T����X���e$����J��4r���縠�<x���
��Ԝ�a�I��翅����^�"Z)��^L�"�4��%�q,��ҾH.v�ȼ�����?j��&WGK�A�%-��"�����?���{v���TqpE5� �~*�1�`��N�=X:����Ǽ�҇_�3�����ɲD$f���Rm�؄�����i���=}� r��������*������ΐ��@̏��f�<���N:{�Gv�L��N�����u��]/ja)���?���h�$��)��Ꙟǵ�5��A7y�z��0R�#�����2��z����Ք�i6��3ͤ�;��r݋�K6/�!��US#�k���.��yK{H��	���Q��;�5Aud��]
���-��ix���V�[�8�t{b�=��:蔯KE'܄���{�8d����=����S�b�QDNa���s;n��RB�¤���H�"#�⯡����v�d�����L��m�4y����S,�S��,X���#C�M]$67uT)P��Zc��P!���IT��F���T ��.ݜ����u^�O���F�ٓ ��:w2!0�����R��>i[(s������t�u�tM�@ε�����h�a,�Ac(��8Oq��P `��1S���g��L����ob������41K>�wQCt�)
����%�1UB�O䬧�t�1M��ݩ�P>���˾E����J����E���ޖ�КO�ۈ���0��n.u��lw|��YC�}]��N���A's��V��w���{0�-@}q*�������=����Ӽ�j���/�L�L�����n�9u=����"��M(V,t!W{��{��:��n�-y�C�lP����U�]]Un��D#�^�tb����xgpM,��,�ط�)2�n���@��:�K���hh����7��{�Z�A�i�^�0Egp�
�nLr���1㭙1��8\Ưm�r���GS�����)�׃�`���@��N�I�R���W���*���4Ӻ�>���������Gi�r\���@���D�P>�c���=S&V���qi��@�꒖Ǹ��A�Х���X°����o�)�lt���=���Y�r���������R���.���j�,���*�p'$R���x��9�"���(w�9�%���]jLˎ�s>��T��n&$�7���ᯝ�cZ���-�8��6n�,��4�b ch�-,�<46v��nr>�&՟�-�;�	H>��\�7�Z# }A�e	y*vl�d�V*y&88Uڤ��ְ�Þ14;�/��@3�����Ü������]��WZ��������XQ���x+t-ȋ�el&7!M+߼��p��.��O���$�^�$�=U?�����>?40l_R�c)4�>�2mg�'�C����1��}�<�07�F[����<,1����'�gq�1\ͯ���4������WSk�����,P���{I�h�Ks,�	�l��7ks�?�eE�]#ͥ�nBd�L)���[CB�TshF���i�@[��85"�m=��c:�h�hpЧT½�`?u�5NA:�}�� ,��^��I�������=���%m��)�O�iOC��M�и���1f�:���|S<���.q{1fNR���ɉa�ЭT>��ܳ(<n��*Y�f� ��M.ԧ�|2_���U����,T�����i|ц�$�	a䖕	�C{��@�iϖn
���4e��}��\�:5)9��B�[rP�;ħ�R^�8a��]�2��Z�c��?7���;ƣF_k�L�QasծЌ^���¹%���e�5���h����"�TK���~҅cruʜt?N�i8����Q�Zd��A�40�滇Ԉ�#4x���Š)�d&{a�@Z��5m�����AW�Բ��5yO! �s����q�*k���LS�R�	��"�O��:��b����
h�uF�ZUH��76G�*�?,��;�����cj �����r ^اr������<�捇z��g�z�0J灑C�	��X�I��ڎ�|��?J��j�\γ��]}q<	%��`���22��2�M��ݎই�@�$��I�Q�n�x����NwUjg�D5�b��5_N�JBԁe��uv7�M}Z�[���*V�t91b
>}��ql	�$����NJf�b/���ʇIlȀ�0���{�?�"�і��(�Ϡ�՝�Ǵ�ì�ͷn;���V��_~q��wGHx|�M�NB�ِ>k�+z��c F�US��K����'�̣�����܁L�����\�Ak�Ⱦ6��U���̃M��N; �9q��Y�xW��y`��(��6�C]�֔ϑ��� ���'F�	^>��Ġ�A��Ƨ��쾷�[�]��j���sb3�
�\y4�%4���-k���B�ߘ���@D6V��ʥ0���I���k���xd�0�F+�v�!1(�_�2ɲ%���<#9�P������曄1e��, 1�vs�o:v�,1��	GX}(��M2�/vb5�柄AV*���M�nl�`�&��,�����;����s�t1r�ֳB�71a$u^��Ԓ�.c:���}��u���4hS#n�rk������y��n�h+y�^�<��;)�@M�`� ���Ɲ庐����ذ���x��1�N��ki�_E��Rn�V�w�Y<�����\J�~�����q� s�\6��(bu%�oF�W����>�M�p,X(P�erP��-�"��tc3���z��I"�D^0��
�HǈÅ�пj��\_�ۨ�,h�^�YtΎ%��ʊt�R&��
��A���P���Byحy���m��vFȾ��Z�=��E�T����O�a�͂:w�Jq�7i��Bt�B�@�^�hF/��/��)9��l��n�1�܇*T���ͨ�ZA�����$��0d��(�$|mP��x㿛�d�B��;W/pB�%�b�n@9 Wr���׃���@���:tY�Q��Xq�&�,�>ۉN%��>W(�����yx��=��#ȜL}����b'0�ʭe]���,ᥧx�e�+��[�H��Ǻ1�˨�$�B�_'�?�!.c��Ͷ,�|��՚�(*��A���aW�+� �"$D���r:���f$�gk�m����W&������bV	�~�~ ��h���P���`�\�b�?e*��0�\����޸�˹}4�P0D{(�׆����8>��̘�g�W0�j�%࡙a?܁�E~^!v�����\���CT.~{�es�a�9'��)�+����D���X}߽�\!D�A�^YJ|D��:A8�5(�֖E����Pճ�Lݐ<Nٶ�;����I$Z�=]d�'\!���
�����Si{���#*�Խ֡:-ۏ��j?�=�c�t:��]�	*g�ZJns���WY ��k���`]
���!V{�S[��@��@궗��XV#@�p�x�{�X���,SQ�*\��Yk���AS���>��>+KpĸI�x|��o�]�J����x���;�b�º��k��`vc����W�w��M.r�V	��"$=�+���M3���viY����.x��g�Z�qؑ���.ދ̵�:��ۺ����؋ϼ������ ��ȪR��v��g��=3����J�c#A����`m�����-�4��:}���Q�5]uN�H���M����=�X�w53���iɲeW$Z2�sz��bW���4��=U�^��X�쩌-�� �n�������9Ga�D`D� 鎫��n�̷H�F��x����B�����F��z<�m��́i��'��	X����_�m���������n#���/P@��[��I�J��晤8􁣉C��/�֞�3���H�tX��/��T+�rxu*�+��� ؝X��7�-߹��.�l�����'�no3�%{�43Xꢉ�0����a-�B��f��m��;♓WQacn��B'K3A���1ߋ|D�Hڇdo�
��M9�GFN^�Q��ė<
c���ƛt��8�ז�Ewt�b��z������dTRkWt�K�>���+�;}�|��S��"���}WF����|�;����Ҥ%3��1�`�+�+��s�@�����{u��hʡ'*�]}+X,���bde�oJDc:�ͥ��u��vC�̈́	�IGZ�����]����w�����B�0�@ɑ�"W���݁C�	�A_){��qߖ�]j�M���292uS���	��c��׀�2'�N?�9w鬒d�5���b�H�`���t�� M;9f�+s��m4�M�]S@��%R�����f�J�v
~VH�ST���f�.���7����d%�
��T�PPZuWޡ��oX�MaMp%���wQ����u�s�]&�q�E3��JN�,�[�;-V3�aW��
���Y�[�B�����rY� �_�a߃�_㗎謹<�3g� �k���s��oPǾ5��s�!ޘ)�@B�����64�g�8�0��(y�%d�!Y�$�G~˙r�Y��pg���4�}��Im
�ݻ�F�vQ���s�qR���JFܕ{�+�n���'~�`�=m�#e��yUB"M��E�����$C���#i�C֤�;Q�'us��B�e���O�)��,	+O!Ԉc�1MR�g�[$!�6�DHl�
7�Q��|�Ӛ(P�=�������?&����wD�\����@r��) VIAG$��qI���s�Ӫ��=�ֳ��;������U� B���1\����7�t|�f�أ��:����մ���p�uB�Bp�SB��o|�?��j�K�`��eƔ=��ן�qb>/�&�Tc)��=ˤ�%�u������CaЎ�/��`2^�����ͨ/oZ�gH%�_�]'�Gxݮ��� 4�/;:_qZ~i�b�+�q2��X���Ԙ�!++���A@�:������J���F���I�����eܫ��G)��<=����3?y�ӷڗ�NԯI
z��C|�Q^͡��oRnC,<ʔ�N�"*�M���Q�.@�����rΉ`��[/��Qy;@Қ��T�W� ��7	X�|���/�B�W�m�M!`j�h�ȝ��� _�4ZdFW����v�m���G�,7�|���!V�Nf��:�mBr,�3�"0}��
��`�wf=�D�TiՑƖ����Yf� �,�
^�AS�	�0�u�9E�,@��|�&���i�$�N�	��HT#�&&F�H�n��6?�g:��X�$&#qg��@nBL�5�[��߹W9�k�Ř-ʅ�%�fN<�Z��!e�StNPbE�:3DU���[���E�ao�e�M�;t�����=������h$�D���!��R�����ͳݛjjB�-xv�!H0��ehE����/�u	�m��Hj�ܐgs���l�r�lWS�vM\L}��p���Q�������ל�'[lR����V.�g���'�;>vo0��9��J�!�H/�0�Xn�4%h�����RQÔ[�� ��jf"t���5�γ��,�#��ݗ���H�vF����^#�$��M0*9��Bv�.ԍ8�h�s�����S�j�lT�P�ǽ�"]=�kh�	3,�~�ᢞ�2��k��Kn�#g���8H^��'��<��3#�\�7+�y�]9GPܷJ���'*��m����a�vb�;"Ur��,�B߷w�΋�eyE O�N�{#x��MkAy����,��H���V���
V���KA�]M+eo$[Z�D��t���UixL��v�?	�Խ�<U��ĊI��Q���!#������,�%�����"��މZg������-s��c�uˡ��za��p��ud���?I��0��H2'�z�E��$�����SJڟ�Eg��Z���\�#���bR�}��_�yϧ����<��Iu�*rg����z��3��N�߇�rq�E'vv}H���׹,���8��Y�u���|P3t��0���-�n���)4�Dm:�Q�I6�f	�s�̦��w
���#�"�|
?�Z.�:��/�dK����9:��Ѷ��y�!:�F10J$٢��&�,�~�L~�p�8g֐(���h��a?qp�\w��~q�&���4��Y�K&-Ҏa�59w��L���)��C�M��B9|�7������X�.��L��<�@���A�g�d(����d�WF\ķt�����f�������F�¦3�b��'�͜�3I/0�k�e�����hG�{ނ}5F�s�@��ﶤ���.w#�N�?#Կ����A91��ɛ��;گ&C+ka!Q_�H-� Je]�c�l�ph��z���ʯQ.=���u�>P�kulP>[�u�ߪ����;�I(�n�n���p*�.���.Fk�4vCks�k�sk���?�
5���Ӟ�7�u��VےC�巓��!pc��F���e����;h\�9���أ�f=�Sa���Y�?���_B�M�0����0���
��	�zU~<���0S{ɵqö��K�a\K�K*�^���!��]>A�)l1�pw�6��������	˲ɈuH�K2�,���C��c�t�u�t��hX��p���lLc���I�1�9<����`+ڋ�9��P����t8]�S�j�}V�-���j�e`�?0���׋2x�n��.kv��H\)�j�0��;�"9�@��*_f� �Xҗ�f,y�O��E���ե�%�R�^�1K���� |���z|} #r�:��Tn�n�a2c�Q���n�J�!0N�eB�z�����4e������$�K("oś]�,�\��� �4�o #��uw�q��Y3���]����Ԑ)��O1w{�wUYxغ�cO~t��8�U�j�Xlm��wD��b���R��N� Q�LLl�3��Ic!����R���g%?�/z�$p�垛3�纉�ݻ�^���#���l�X�F'�=����t�D􍒃7���`��K���|�־�zWe	����"���g �%%��~����K&[?2������@�-���y��I3�2�0P�Y������.
��M���h�5��b2�΍89��mTߡW6�UN
�,%�IZ�^�4��;�Đ��\�EiW���qM�	.�3�Ka�S�i�4�����7���&����)�r �� �;�N,�
#u\S'�m�2b����i�{k�-1tt�U~T����ЏJn��ʥ��|ũ��}����J���<CP�]<�wV�����U!h���˘�G�H�{33�ڼ>�OY�o��߇��k�)�hjl>��T%�m���j8腧�I�fu�.R�Hk��d0I���#� �B�3us��N
%�Qǁ�ًě���W��%\41(��\��~m}�RV�](�6����x��Bѽ�ʆ�'����l��-�%�����h����9:���>�{���Ä�/�%�������;冿�-�'����W�ڠ�}cƈ��vv��ęX�w(H�Auκ�/WH�ۮ�$�&�(9�Qa��hI�m~�����2��P�%(
d�a�u~VN��:fK�J/ԡ�&�|���H.;�m��˳I'�E�j���H#���/w%x��I�mM��/�_-S)�$�A&︺W.'��ch)lO�rT/�F �Y�D|�;���4��B��ӡq �]N�F�(�Y�&�5<KD����<u8u��]��V�z���i
��6;�5d��tP�V�FC!��	�h�h�qFv%i��V;�y��$L���*z���Ę	�|WS�Yj���͈��3۞�r2#(}Q���_m4��H���//��:���'8V�!�%��G��R�!M�����}36Bs���zR������l�^�6���زKH2.�j<[�H�w��1잰���	�s�P�Md�O����Ad&���SO �R�?m@��@��Du�A���������pvR�7l�{s�N}s�<���-���Hsݺ
�����傽a� �=F.ˮ�XϦ����qi��P��~>쫶�m�Z�p<���c��B߬Kp��ys�u���)�B���FnX�rۡO�b�5�_���J�ɹ�rA�ܥY��`A;�,�s��2�bKa��L�(Nea!��<��-e��kA��q����'Ps�d�£./g{I� %����|�~(��)�0Eը�c��8[5;gB��G�����u唡�>&4��)L'�Fb�fC�%X71+�=Yցa��za�'})A�w�̰>:�Af]�H���3�˾���L������;azI�v��o�������N��4���Iy�z�z�@� �F��<Q?�c��¬͖�iU�}!���Į2�n��������	qiI��§:��b�y�}�-��h
ʙ����et����ex�o�
��)Ou�P�}�}�4U�SSs ���)p��K.N�WM$�����u�s뙉�z:�r��2XԞ��6�P��Y/��5y��B����U�iC��`!��ץ%�C�ؕY(�v�7v��v���{C�;����V�(��P+�'t�>e�^�_.���K�ۙE7BǢ-՘�A�(Df�o�hzz�"�/���V�G���B�[���!�4)�t�K�zv��xG{�N�O�&��}ʍX���}�}�(����%�FER�Q��5]k\�
� ��B[�fB������5N�=�=�Ev_�x	��4��tiG6����������b��]�@�Mn+�y��b�(H���S�t���6)w�R	)���,��7����9�:�Vَ�t��}��$eNX�Z;�ܽ|�Lpǘ��۞�wXʃ
����/$���F�"~J+hXtq�xoyc#�6n�ϩnК]��������6�g'�@q:�ѷ��V- �@N�%Vc���zެ���7u3X���+��WQ��qk9c{(Z�Ѣ8pA߈�#����aӭEѫ6E]4D?����;q�	~�;s�j�$15y[f�H���GS�LG�Q`N7lehR4@�/UaD.V	����B��k�G��S�����.���;*㛸�y`�u������]$\��7�O0�a3�����ח�d���1%�8��������yK(���t$G�y�թ���I�!�
�$�B�b!<H|�x�$n���u��f��BV�GnQ�s@�a���ć��`%T(�"��G��vA�7[����ry-/x��q��Q՞��$��ӏՆ2v�8|�o���>�Ni38�B��.��6a�E��b���ء7K҅��'��7uO�]���n�����_�R��B�?���C��?�'p�=6���]؇��R��*��7�5��3�HRG�i����:J�i � ��=%��WW�"^�'��	�ﵺ �4I"�����������;C�	$�� ��eeJ����4mWGFHj���N����0ąR�kä>�k�;M_�5��F�5�O�J2�Qa|�rwlɕ�����1��)�a���ނ�ˣ^y8�r�`2 J�?M�5أ���)�gy��>(���x�;�z�	|@��}HX��@β�S�3�G�����WXn۔kP���ȜGQ��%n�L�5ti7I��݁:�ʇ����F�3Z>-��5ұ���G 4��en4�U�h�e�W�c�?O���h��+��x^i�ڃ�3_"��r����u:�屢�V�;晼2�غBR�j&l�<G���YI,�5=^�(C��ۆc�N��H��<3ZÝ�ŷF�^�br�0I�tr��l��q��A������ἁ�154��L޵��w[��l��b��Q���G�a�C��a׊��&)5gl�������#�s��S�������v�x�����8�ť��?v�^�����G�Np�����(.T�~z��G}p�6���G���N|_����L�~i�e�^?��п60�x�)���և��3c��fb��e���J �a��m]��̘?���ﺓ��ƿ�.\R�{ٝs�{�{�a�T�2���!T����hV����m������K�ʦ���{��>�<z���D�	�W�e��qr7!����D��ļ��J�>�]�9Z=�u�=�����KL'P�h�� ���13�;�]ho�>h��yG�J�m��p]��hެ@soHu�~|;ʻ��RJ��uTq��em�O��f{W�C]��O��%�ꉶ�Qiq�r�Nz�O���++�?3iǤ8��ia�=t�H-��u!�TU/t���d���C����nmfH��:�_g���תe��z��ѷ.
�?�Y�C���$ܭt�U}��ߋʑ������o�P���l�icx\1��������;� �-�S�崊��ϋ���W��K[ǘ�\5au2%����+p>������9��j���� U�E��c����{��D�ؘ�ු� ��(
�YO6o5k܈����c��Fv��"���,��\�E��l�Iw0c�V�N�!�7�~	�����h�����䳰�g�[�B1p���e���VQ�z�K���^��ύ[oR�M@ũ�n��4���`\���H��/?��_B4a-��-,^4i`�#w-4y���Q�r�<�[;K�����Kg��gB.O
���.��!�G;��C]Ĺ@�z�/IK\9\�Ϋ�Cz���T;%>*�2,��$"�Fg��.ј݃��ΤS�l���-^�2���ھ���"�>:ó���Mb�Oz���`+��U��ĕ�j�L7T��.��7�Z�\����Ȗ���]t�4l�MZl�3�e�9>9��l<�o�Z�p�9q�EG���$Rۯx�^�bz(����H�����#T�?p�?��(C1�/<�[��r�b�Wi]
|���ϣ�JRA��[(�E��ϣ��%l���p��(�����-)j��������S7�#���}BXL�U��b��|��T�b��!�0{��k�g3 �êȮli�98��M}����zD��A�kI�DB��0
4Kf'�?0��~&�]'���ئ��*_��y���0���n)]H�y����*�!���lZ&��yN�:P��d���Gл�(T��U�q ��FI	x�"<T2_<�n��0 	~�^�;I���"�
�ht��\>=҂/'��j0Y�i1��b7��������z��uؿ��1P���.I��������̒5G+P�A�/h�A�����+����+�y^}	�� ])Ɇ��[V��>�٭2?UH7y?+e\=c���C����7�/$�Or?�T��3���Z@&!����)�5to��CC��߽��م�o�0�H���黹*1���
Z��_Y����j@b�`Ȼ�Q+4�C�س��s�*�g,\UT�>���\V������b~/"ؗJ/AWa깫� _�����d��OC_V;<�ZWU�1+މ�@��`X#y���J�qn1O?O��$sJԟv�5�IAU~�!|RO
7L'���A�x���l������^�-�j�~)N��&��~Ν�M�:D~i݇Y��VKp��b�d4c��p������/�ڀY��l�4�W�T�*e��?��l���>DӓW�AL��OpHhe�1�GY{#`V����j��Hh8����o �y��$mʹTr��IK~���8�Z{fA?�U\�m�AH���sWf8b�rϑ+�"a�-��;�D�!�*�͚i�3��X�ĸ9AE%�o��t��g��m��ܛ�D_���G��ۥ(1� ��J�4i<K�e���(M�`��4�Eb|!�>_�,bLkq�y���h�_̿gT�C�Ű���=�����h]�����7���#�֚^�(��}t#V)/�CpsЩ}�Wj�i�ʄ�Ώ�ո�����o�φ @1K̜+/�[�RUD��&�Z��d6��䶵������⧡�[�\��7P�*�������h�>D�m����g�}&���ި��X4�^���n9e���C<���\Q�P�qE����S�l�.j����0�$�j@G����
���\��P�\C��Ͻ��)����H.���2@M���m^���Zʭ���4>��\�$�ysEsDdj���m�"��}`/���]�i#D�7�IJ��K��⡊THݑ����b���%�f�\)hGY2v�f}.�r��aĽ���"p��x��u�ë�R�9]B`-�RF�?�� v�Ν_/����3���k�[5ND�oO�y�Z�����zL�O��b8H?_7�*zQb���8����wR5�*����g|2����Y]B�Ǡ���,8�M���K��0g��T��K	a�JDd�hS�&A �3|�)ҹdź�����Պ���J�9�@
l�+TxP���q��4F"���Rͳm�H^�B��p�I��b aw�"���ԍ�"O�3�>�ھ,��1��խ�y}C���.#��0Zט0��&m��,	���,`}�P�5�~R�Y�s����ڸ ��;Q=}!h&�;_�x�`W���^�Y�A���'�BI�H3��8��(�ÂS
w~}{�-�^j�'YQB(��RG�F��"��=��+����?h <����NIll�i�_ P�s�ʣm`���0�:bq� >&���z~��9�=�>
u�F�B�:��W��������~�� ��R\R��{On"'Ō�����#�OO��[@����&%�B>���FC+.�Y�v��+zx�U�{{}�3�<��v�*�&P�&J��7fL����<}E/�wqL%+�S�7B�k܍�d�.�e'Ұ�"���0������tZ��j2�ς�,W�=���Y��)+{�KM5�c��R+��!Y�f螅g�N}?֎3�̓	���4p��u�2eY����X6�xG�rԳ���X�&{����C��fo���z�a�m�/]'���-���.Sb�`�=��9ώ�C�H.�;��'��Y��\s%��\R����Z(���@.ڨ���F���&�Y��.� ^�xqAK��"�ܣ��;��ȝ��p}�k~K���-�<e.��F�O��~c�˖�fh�	�E��8͎���R����k}p��=�Dv�%Mƈ�D����乵nS�O�j�%�7DM�!&��إ
����k�۲z�z��_E(�I�(�j��k�"��,�S�̟)Ь=%�vh�s�Z�?[���B��U3w?[4���w$��@�qC��Ns��V}�����VC��v�����7_�h��H���D�h��Ǐ�c�R#��q7G����zBn�f+���u��DB����(�oi��P��7Eb��lƀru{ƌ�A5h$�d�����J����#�zo��1�n�2(�_��(�!���+E�^w�;��s0�%��? 4�
ė�p��8��=h�#7L��%@��g��S1�I���ڐ9��+���=�[���W+cT����zO�I�6���|Z�%�����n���d'Z�C�LTa��%��	�v�OZI4@�H6@�C_k���;#�mt�6[x�V���BW��_�>�Y�.�v���-���Imhn��[���`eHAՃh�2ƨ;����9��a�2��tV���ư<HL3��-Q�l���:JqM���~X���x�����������<'<)����EyLE'#V�/�I1D��rkv�'ɽ(C�8��@9du���r�#0��rY]��7o��x޺Ӌ}��\�k��㓣�aQ�\��/OQ�9����>}�P��d'�9�ޓ�y�a�Oe]��	α�ؚ��og�f�J����(�c���gf�vm��m��;~�'�ެ?9�^�A*X:.���8:�"�J��Z��MN�A��^+��j��f!�(�%��,��o9!��&�8��(�p���"_�_�3���{�Tǧ0?��AE�L�HiOQ���Q$��/w�gC�xJ5�� �Y 	*>���"�_5ÈS�1�(�4̘`'���m��%.���2��B�)u�^�����)l��m"2	#*�B�r� �?��