��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~��OMa��@��{[��(k��cm!��.+>��U?&x;5�2�,S�+uW��	��T�Feq	��h���ؤo��?&���D�P5t��/5�Z"3�m���D���ͩ��B�&�~�Ѫm��^o�a�� �󶱗��k@�Nk/����������Vӭ���r�.�
�8��x��t �]!�{X[iJmLD�hN磊�H�_e
�tV��3Q�����y�j��ש��x��ӝ12����KÃ'�1�&�8}NIw����>TK#ؼ���G%�C���u�5X���b�r	"�\�G�%b]`��b#�ݼ�v�FL!�Sܸ�<ʋ$�i��Dŝ#�y�	&n@�y���u�,��E�jYk��NQȚ'�3[u�?ˇ�У�+��1; ��J\\��ٛ���{�̄eܘ�+k�#p�ͭ���.�3��m��`�[:Ha��y#�t_�0���]��ܚ���V�nN�{���L0�G"���]����&%|�)τ(����|�]�$$H������$�h6
�#��Ô�M��SPʶDuTw��,�sJ��z#P�W3�����B��$���	/���=`G��2L�;p�-��ര�A�xtG��ޫ�0� ��M�?w��8��xoi2CVP|�s��R��E>?0_��L�^c�f߫˦�p����~s�lw5	'T�ԝ�Wu�u�]��M�O���fg߽
�M��v\�d)]T&�x|#�,�1�g�j̅y4z��f�X�z�����Ô�/���¨��a/��3 ܄\�5q��g�wC]���Ç�l9w�����v�����L��?�H�>��R�;�P���*��ͬn���ckFU��⿿�wX�o�@y\f[�J?�إ|�������Jq5Ͷ���s)�z�z$x�z/:�Ef����c}r!lo����*�#ְ{^��&sJ�fB�^6��6T�Zl�w�;��~��◘�x���
"���;#쬣�)�Dݔ�U�t)����O𝗔��a��맾Ͼ��������:�7P!���Z�꩛��������-//U��������q�]��lE�cV2(h�%�/b*8f3�g���I�	�BZƬ��י�w�eF.0���S݃�:�P���솿$ʇ�(��$@�����S����f��,8�|�A�����O��.�����|����n��P-�m/
k,H��z��g���[�u:�Yo����Cx�O�
B',|R�vS����5l[���G����X�e���|����!����k*��K�q�ZG�G�*Ǵ8&���6��,6kFͶ��k��3,CPS˒.�:���ޭ
͜�o6��ld`��Q�,�ήQ��@���s�ͥ��dt�ݱ��J(dZE;̎�~���Ps�&�*\q\���Q�T{8��<�z�j��O./:�щ����;�ټ�ٟSI���+�]c�N٢���6��ꒊ����ׂ��Qݏ��0��7�ES�+��vF�=}O�����A#^ڑ�-#�F�/�|�7ڡ̀����5�8�L�_��s���m�H
ƭ��z��C>����<�-���Ȭ�vH��݀ۅR�l`��Q�8IB/�%�k�KZ	B�1����Z�_l�dv]h%��{
�99��b+$g�\�T�k�t+�;��]�Ԫ
<D�����Q��ս��)Ԛ����g0��e�<�L�r��k@{-� �Z��� �O�@3��$�hiR����# ���I�	l�+��1?��O|û��t1�X���
�5��G@�ڠ����򷍧lw�d1�у�O&�t�`LI�la�/��u�]׍3�P*;P��ϯ��#ֱ(㘘�.�Y0fy}I�*��ĵz3��&��L�v��K�$7���Nj:�8�%�����Q0�����e�o��$ѹ�]A4��T�e�h��^�[��N�[W��1�q�q�8y~.AՋ#�I�WzfX�����V^��|ߗ��O-ޗ��>��S�@z�D�:�V.�- -��R�&�8��Q���fP�4�4f>Td'Eq����h���",/�����݊��;=3���IFTF��{�����?�!5���?�[�ь��xo�z����P�1�o���k���ܬ�H�a�"w����	?u��3��������e>�pe0�s�kZ	
������'H�Mr*ˡ\�H�[�R����v��1r�U�6��J^ȁ|/<�^;Ss/����P~�G�/*n�����GxD_��ϰUG㢧��T4g#?)��2�}֏�-���sTR��tt����ks���/5�S��Z�SI7����#v,+�&6X�R`b�EZ�>�:X��ϒ�x哋T�<��U�V�c�{/eb,k1�4�G{�Ƀ[�x�+�^��}�ȣza��"�Ql&�-P�oK��L-�
��V�����&����տ�s��}�=A:O��{�d{�t����(��P4���!t��!<;7�@gİqd��܇��ح;g|�j���XS��g�N�ޜ�鱁�o1N�Ho�`��	㱍�Q���������t0�9e�^������K��d��NcEܴ��Ubs�S\�6m[*e#g����C �.�X�C���}D
�ו$ND֕��ql�b�1�x�ySS�,o�lK%>&��wb��yx�@��v)T,Zғw�s�lև:��x���fܠ��,���&^-w`#�fq�𰧼D@��Z�-�^W`��G~�F^6Y�]�&�]-J�#���alW-��E���6��e�rZ�d��z ���"���^s�R�e���b�;���O�n�����O5���h��J��Ч��3X����o�P9��{��{��u��%����H?	�Y#���<F�>Rs���
bm�qb�,/;��w�I7F�$��N&�4o�,��Ɏ�޹F|Z��d�<��L�P���o�cŨS�ޥ�^[�''�����Ed��v#�fjǶ��1���JB�d��?l�"�Z"5~��۳�t+�bg'�\Իe�]hҩ0��zR�A�W��_���ՍI�#e@�7�KJZ�vG�/�+�N7�\LK>�o:�%�|���)D 7��7�@��:Љ(S�o��S����+�`��O��|�k��N��7�!;��m�斃FXL; ݪ�����%��V�i�.\�0��w�nP��܉
|��s p�1�r)2��	喂K6��1+6X�Rʌ>M������Bh�"�E�Ȣ'6����PE�?+�����A��[.���g�>������g�R���	��n����J�H/ 1�UM��4���-"�Ϩ�x�p>��D<�cf��\S�9��{S�ˋ����]�{��i���K ���Y���z����Qk�>)��7�?Rg�sb:�.�u��E��Q0��/������ �0n����J=�͜�^�]��,�K���\�G��j_SG�-�b�<�\YJA��O�ن*�gH�fh6���@�X���'�vz���������:rϰ8➍��z��"J�(�>�|�&|�w� 8��?5i�\f"�"�Bx6c	a�n�w4���/�eYƉ��t��B�ϪQ�ۂ�*H�$��(�iy����S�wS��>a�&�N�v�I�v'?�M)��={Ҡb91M|����
Q�	������(��d��Omټ)9v%��e��h�S�L��&����c;
�K�_T�VÌ�E����|u`�������
_`���>���kN|7s_��܄�@�HT	���'��Zfw�ڐ����=n�����������.u[�rx����_j�n�;s�NB%�(ܸ�|ӌ��:�;J���W8�		Q�k����ӡJ��0���CC<.\ذ�ݺ^�0��{gtW����������FV���q���-[��F�I&&����I�a�����Xj|��R?�S�j�����qc*^�<97\�+ͼU���_�㟉V�W�w�vN��[��:�4~/WOp���B�����}^^��8d{1��	k���������_5[ӓ�~�4z>l���E�%h�a�����K¼�U���aM^�"��6"��� �~䷘,w��8T��_ZR9C�$���X�)v�wڀ�[��+�\� [�y�;m�\��aJ�΁�'�+_�!S���p�C۾���ס
7���T��MD(᭐f]T���7����{+ۦSj���w�#<،&���5��1�F#5�U7�D�M�0���x�'��UҎm��Hv�+Y��R��=w�
;���O�-I�YP��l
 X��kh��v�& ��c]��"-��i����?be��t�Pf"���F��!E{�20�Y�M)&�e�rTS��{��0	�c��x�Rш7^�jM��BH�ߚw^���[�z>
q?~F�iD�¸޺Q��I�dPd��)$�P;��-��E���
�2���`�"�KI��X�4Ʒ`�_|���W�X$en$��]�֏ZRz��o��7!J�S@��; z\b./_��eՊ�\�2�b������T&�Ӝܡ�����UжC8X�.����m7zQ���ֻ�F`��)O��ۍ������������J�{�aY�ۻR�o8�!���;�������I�OY�)��6�^�4+34�u@3���3���Afcd�%E7#F�`id�S�74�:�oo�ٳP�����,�4�h�e[�x��IЁ�����Xu��Ձ��Kq!�������i��r�+_�`�CH8M+*��Z)0u�1�s��aw�Cߞ�FJa���sY�Ű�]�j0hAԃ���I��<�Z�1��r�Q+*����4gi�'�r�So?��i�^>��>�,;������QR��N��bQ4��m��
�DJ����*.D�S{8�^-�������UjÌ�i�}3xlAE� Jk��*��}e�& +�&ah@f��FR���v�0��:0�d����w�����[:>C_�:rbv�k����'��A����*$@����A������lD�� ����ER���bX���T�E:����M��&�,��́��$��P�Waݓa�qA"�e4mq8��]:�Ҳ������`��,�����JVR>���������O}��5����ԭ)Ⱥ��eA�A�-u��{�T��ן�6�ˤB��!�q��ݠ��z���43?P<��9l;���d�-�>4���1�t���SKP9�D�w��9G'��Ň��	z)Y���ZLxJ���W�-��������fY� ��`B�Q�����in#S�#���i\�S�@A5����y��q�N���k�$��rI�Vy_�).�$�2�Do1ݔpժ�(��s�u>��;)��]�*n�[($�r3�4D��x� C=������yX�^<�1f��\g\�M^fDZ9m쨶&0 ܘ5O�}ּ�BV\QÈTJg6�vZƌ<)M�'P/9�u��'9Ϣ<��h�����ÆE�IlQZt
Q�P�/%TGF<^i� I�)Ӹ���-�ly����l���g�6�YG�n�׺<gd#piYf3�ꞐjH��/���֛���r�H<L�Ud�ϱ�Ե̷��ExPS`�.Gb'/��yx�	����[����L�e�9��Mɛ�Y"P^P:�	*� ��+	��MMYԙ}�)�e�z�·�F�Of�AW�;M��QK&I:�>r^��F�)�2�`_�Ж	�(KUC7�.]Rɪ=4�k���h��&A:l'��o�f�1qz���Q/U�٦�©!�S�F`k�crI�	o�c�d��G�S�k��(_��n�¾�W��D�d���C����S�-�x���@k�3��|Im(QxK�5o
�y_p4��t9�7���x��p��.�g��7ɱ�5%Q��:������eU�;'� m���.�~&��d�.���?�����u7W{�{*M/�!{�C�s���Iُ*AB5l�cf�,��-?�Q�~eG�����Ц��0���[K��Tސ(�1�jiҝ��u3���#<���@!}:dlTږ��ǚ�\�������Ozg�JŖ���K�aī������%K�,�DHl�v��[Jvp��J����#�ܖ]����	�Ju���+/M��� �e���W���ѷ-��	ĩt~ ��c���� �k��e��RcQu}ŧ,��5�{ܘ>��0���<>\|A�4���M�>!�o/W�=��ĺ}���a�c��Զ���nit��':�����>z�u���i�Ot�4��to\U������ƭ
�7��lT�{O��(��!Æo�H��O�|�36�4���!*�(2������R�1��_��e@E�s��&��%D5�/�x�Gb�'SztrQ��W��9W�]�)2�[K�/��#��[=�5SG�d�0O�`�Œ
	��L{��$��Ѷ�g{�&��eC��#��a#�q¹�B)�C"~D�Em����7�f�E�� �a����Q�Sc[�PmS�O{6�j%E����+c���5��a��
�[E��1!n,�y����o�Ӝ\VɎԗ5$���גrJ��ɶ�bF
��R���[�[%��M i��t��x3L8#�N�57�������4a��.���1�v�y�Qj�Ydҧ�^�5�x�x��w�do׺������T��|92z���0ͻ߱E�[4U��5�7�z���VɈ�|�z������*��~�r"��?�6�]"l����_��z��d���g�R��9�f��e�Zz���B��%��w�^-��9:vϋw�(^���fO �e����}�@Gp�R��fF�;��ω�vz���z�Z	"�qEI����(������ܷ�yۙ�Q��a}�Ս�y����[c�TlT%1	{�/jD�\�X $J��	hQ�@V���0��L��]`�_G���ǻMP~4����2�I.��(��O�Ԥ��-!|׷��j�Z�}G�!A�!��q�v�$��N�@̘�X$p�F�4z���=��=���U�-��Lsl[�U�沂4BT�j�-8'��6��:~��f/�3@e\���3;Xf��xM�x%�g�m:p���Ȋ��C�ŚC��P�j�)L����_8o�4���6|P�bHgF[dh�p5g%}sȂ�����V�K��'ch ==� �|�S_S0��32 �OY�Y�T�M��o'�.��1v��K��p��-��gG�d@��GnY����K���ݪz���,��oR��Ծ'��#{o��g��)��l`��h���ֈ�O �8�uOM#D�
�F������eq��D����!>��ྉq6�o�a��� �ߒ�'T�\^͟����o�% ���D�K�UܵbƮ��"�fml� $�h긗n���We�%�>��i����^1����(�����Ǡ�T<o��7%UrPde��N_�le���2�~ 9���4Ĳ�0DK�2�*s���2��&N%6���X}��IY�܎��eR���$k.ChӣD(�S��%���d*�V����䌭+챁�v=�(L��
�Ae� ��I�"����}՟bOz�����ӭ����`��%
�q�E����Y"���9�%��[<La�n����(F}��>-�]�{������d�r�r�c�ڊ�����h�&}�O�8�YN}ԓ���Ѫ��a()z=~�C���b�.Y�����W
	J���\��B�A����=9
B'���+�0p����RF���a���u���'�~�Ҩ�ǒ�?����ۑ��%RV�-���h3e&�õK&���Kr�}��VNb�Р��#�V��-i�l�I�l8�	k��r�-���v�z)��Å��:O|����)Y�w�'I�O�����P-��y-����
�����Wl����g�d��T �k��� �μN�`�M%�Ȩ<S��L~�1�^i�ݔeq|z�_�=2�k�	��ͱ���gˆ�,��MM{�}����|h���&�E��J�eе��cM��茶�ه������dP���m��ݦ]��fĠ�{t��3��y��Q�~C'M1���!"��Q�s����xf뚨@eYd��x( �+|����H�b�~TN��&��} �ٔ�W�4����@�?��k��T�e���h*���μ�19�!���K���l״�����~�� �����.�d1X_o��ځ���
�V��5c/������
�s�kE|ʅb�����ߥyӫ�A��@�K� ���2�B�l�8qKe'��+`�Rc������j���^p��u�_�A;v��i�u8�7F�օs����/œ�P�x�ʾ�}U��!��6h�	�3�}#��\_~D��n����D8����bK��h�X��4ŗ�e���ֲ���j�M�_��i}8i��РR�7���w����[�r3�gҮkuh'{�����\i�˄��oysA%�N���LJާe�S��)_�K��'��(�
��=^�OyLy�%�3VT�F����W,�d@�K�^����!"�q�ꆒ�����$�ϐ藀YG!=ɷ����-�O:'�U�4\��+���H���:
s��7�G� `o=��]/����<`�=�QWth�YԶɜ��E�1�͜��Q��xǮ\�(
�J*�a{��ަ�� �Q����t�>V$�EG�߀Ab�1�z#�X����3����Ŭ��i:�;wv���d�ڞ(���!d�/�| �/0���j�km�_R�&���JBM�D�sI�)�0�!y2 ��Ss���B*�Bҩ��ꉭE*��= )��"���	-�nP�/fG�R�����+f��F��{����:���쪜;f�ٜ��ƟCժ"�\\�L�s�����t3(�2sb�n����J�X׎@�:�|?��k Q-����/��i@h�}Z��h�*�o��P]�BJ������|=S����CKd��ޠ��T��N��S%|�J�#Ս���a)N���B�i���e�p_��ݢ~�)��^{��bB�'�6x_%�c!����>0$'1+0��#_{�9��/�¤mBF
�{����M#���0}̡�
�|�~�X*�b�>��C$���ߌ�!�B�>��gb�(Ɉ��h{ί�s��Ցa?�� Vm3P�K�JoJKY�XJ{D��!|�����x��&����(oyI�N��'����D�v&$
�}EP<��e�v�Lvo( ]"�B����D�e�|6�(����v\�[�t"L<�Z�gP4�+�<�:��C.��R�ı����6$z���:k��U���c��: -�\���v1��S=�(���� �����p��İɞ,~o�N�EMw�j8���߳��Y
�8���\�ᰞ��2��=Aa�c%�>��}��[���U��2ϧz��$�l��nG�T��� ��_�p�*�H�H����/�q���A�mu]I�� Ϭ��;���&�)�6LL����Q#�b
5���≮������c�MDe�2���E���2�?� �Ot�
�>s|��uG2�߮醿y�D�4��Ʒ�K�0 +V�x�j���Y�>E����z�SÌ0�G�g͝�\t��@�$cj�����.��rܠ	���}��Pt��ݨ�������j��S�^��d����4�����|�%�"sYU��c��ty�m��_���ԦB�.?��I��X0�M2k���M ����a/w �ҿ5w�ϢH_\3�q�ZܜI�5z1ۺ.������j�kª޼tHD�q	>"��P�oK�K��F�6w���bہ�г
�:BweљtI��|��#��`yz^VgF��n���ɩ�{�,+��q����`��~a6O*7�8�{�=""��F͈���^g�%�y����C�~�����F�L8;��[�v�R�"���O��"�<g�>��卛Ԏ���6��X�%0�4����k��:o$s�^Q%N}�{)nG��׫.���0�-����b�#ax��NZ2u0~�޾
�|	Wrm~�Ϳ/>j}�rT�߀}�d��#^�2l`��	q{�yK����7�Q7�R�7�[��Tgѹ���T*?bq�y���j���Y�|��V�����4BL���Z[�Yq-��<q�����I�n"����}?jd.�D��"<R~Z�h�y��ſu	�>�6�7-3s u�����gy
��u7��0��8c#I��Ԡ����辔yu�s�_�"��	�}0C�HVJbRȌn�45��oQ����G	s'Ƭ��$x��a�7���9ܺM�l�F~cQ�T��0����n{o�п=$�s\�8k��k����nH��x
�N1��L�+�+k�� ;���c5�kx�3h8��z�uf�+L�9[ǘ:*N��N�g�]�o�՗4��{�<>�݉������ Nl iݟl��(�'�d�C#��}�[�%��]�}��D�G��ñS~���,�@=�+�u��Ttq���dz��� H��%X� {�3��Ӱ6N#Ǘ��[�x���rxq�S�H(ƀ�c�����4�Ǹ�F�[��1�����O+�Fr�v�蒶��4,�%���دo�q����z�o]�M������a��M�����e��]Y?>b͕b�)�P03�}��zua�<6�M�ʅ�a��G��N^*NsQ�V/��8�7�jܫ�
:��4ǰv�5y�ha=�I#�s� =j��9�a���s���ǭ��|��|���"o�����y���Ŭ/B/�RC����f��1�>��v�s�ڍ��o��}SZ�҃�%\ɨ��5�;-���@��3O��~i��`h|c�t9>�ɢ���Aܓ�������]�'�V�M>��|y~R�[���ޕ�&e�Vս�d�筢��}�����~�1~$N��I�w�����֛_0:J�)z�����GS4�6�/�3�>z�I�┨��������r�D��R�Ǽ#)��':"�7�_p�;H#�������R����K��}�gh&?����]���F'���������#Q�=�R�D�ਗ਼�i�m��m�J���������R�9�1C1**3<���H���ľ#�Rj8�;�$ޖ�����D�~TH�f��=���HQ�!�`�yF������w5�l	��;�>;��^�7�P�8����\]����pAax�|��K�eӷNJ�ļ�4��M
6bѧ�Bh"|�c��[#l�@#{�^�hFA�,�$v�����%����8�O�h�eN�(Y�*FR L��:���c�$W����� ��!�\(�F�]ھ$�;�ǐe.�'͐r�8����xV��؅�O37��h|d���\@�z*����l7-C��Nk%���nmtcO��+��S��xR���n��4��9���1N=A�u��;���cx�~ʘ�(T}�ױ��e.�gL��&ժnQT����Ԛ1#T����MɣJ�K�v�(�G��ao�r�㚠p݀�xKr�7�v��݁�X>��{����?��ۥ��%�y�`Ƨ6Τ��I���9vB�@y��@��Yބ�<4s]�ًB�o�:����˒�'@M'�A'e����ۍ�2W���p˦�ح���2Hr}�j;��IcA��*�rA�X��WI��P[���~�\"�є�Gkh�y��*u���E4����u� Q�^#�j�F�i���6ۊb�3���Ck�F^V�����O&��t�K��z��U���m|��,D���q|!��c��@Ā�Eڣܪ����@Cix]�־�R�{v�2w,�0��8��歯�%�P!4�yr���|-4����Z�(8�n_�B��� �TIU��Qsӥ���slq�����=��ϛ�A��~��J�U�D�C��ޮ�l���	�C�!5^ٽH#�rk���	Lm����x������k\5z�D���,��8v�����oR�T����k�1 �ӏ��KC�r֞B=��h�S?�+\�Y��RM�e��Y���s�_�8&ͧ��؍�[��7г��vy �K���!�X�t�v����wl���5�ʭ��w����B�M��*
g������-��?�� �N��6@��&��i�䞧�L�v��X��g�n��Ju�&�E]�J6���+@ʪ�È}�׭Oi�"�@kA��Ge놱yIn�£������~҈b�ч�"�fW`���^�3���)&�i�9.����O��.��2xJ<gR�&�l�Ӷ��#�|����x���i�n ŷ_٩!�O�~_ �����6!����E�]M�>�Oy:�h%�P����^�l�nιWv>���_��%s���"����8�-_	Tp�����	�U%~a+-�Q��sԐ�BP�W6��3���=��H�k|�&����L\$��|rXP��D��
0��fH	�9���(�E�j x����Ԕ4]�"�1����Eʃ�;N{��Ô&҆�ؿ�q,)�_�u��kv�W@D�H�1�r喫�o�}0 ��\������tZ�ǂNP~2�"Ùv��y0G�0�5P��m�#��(���<[<8.|�O�K�������`���X��Z�&�nWz=�CzO!�^X��٫H��bFaȸ�4C� ��
�_{S.�{��f����d�x����_� ��D�QH?W��7[Ϳ����b#�����g�P�_�J�4������$x�	�j�"'����.�x�]���O�uU��ڃ�񔄨���TW5pi8g~!�� ��NMa=���Z.��q��.��<.�V��*q�7�C���|k}�x�$�W0ٚ�1�]ܧ#�(^���h^T%��DC�
��a>\NW��4�~1������=�πB�;�HӾ�xT\�c���:����&����"�,,� ��֐i��.0�����5|F�B&�J�ؖ��em�܃H3]�V���>y�@"�-$��9B�#$�j�!ta�~��>S�M$�9�S�� �ޑ�W��|�j)/PZ�� o�!�dOc�b2�m���Q?�5�Ƹ��X^��f&�Q9���(u�B��Z	��M�g4K%�M�Ν *��6[�&[�CFq`�n�Ȏ�ٕ�M�4��.��Lw4Z�H����Hm!uXsL�H�ְΟ9�i2�7��8�iw���	����r]s���D���5)�s����윜���?U'ᐃH>�^W�I�'Yu�4�8ؐ.!��&������gT��;:����'Ks�_�G"7�i��ibeqhz]�Ԋխ(�S����g��I�M�<̔J$ �?�Ǿ���5� �Rz9��%�@��Ux�4��V��_�ə�g@��G���n�8�n�#t��ӑ`�eU'��ų�3gx{�wL\Vo��B�I���.#X�}�~﬷ݩ*��;���<]d�f'Qء���~oR

P���pgc��$&Z�^EH��I�M�U�J�߮k?$gu���v<f�U7�_�����|��`������vM&�@��Ѫl�2���h2"s��̞����9{�Y�пwp�lm��%��>t}��g�̀�2`*A3����-�}s�3�H��w���<�?-W�?ωY�*�J�������ui>����of�"Ҍ4�Ta]�������ݺ�,��j�a6?��1f�V���ܾ�����E2;:���G�^����a��o�� ���&��6���Bś.�����K{�-V��F��޼��H�j�(�T��e�Y�wڡ�u,������i��
���\f�#4#v�%�fS����j�'�p�E�b�xNWe[ Z��6w?������Ɋ�C�29O������h1�≱�Z ��^&�t����N�3���އ'ڞ;�_��� Y�O6I��"�P���)�0\�|>���ȔI�,�N��P�cO��>L�gQ̸���X~Y�j��A�*�W���9��j��׿a����&���n���
����;���1���K�u��������F�3��l��q�"�Ax+w�)����g}�	e���#����]M�V�
{�C�^;��v��{@�m����ěO?W�<I�H����po�Y&g�E�G�qpâ6��a>x��g��W�|�����1���*^3qG�9j�LaCD_8�0#�>vm�oF�b{1�����
��/�:`>(fJ�j�O�GD�?�}�$��˟~�dW6��0ъsЏ4��0�M<%�O��$f�wf6���xnW��y�F� -l?��'p�q�d����`��9Tb0�y�ZYH!��uБ�S���B-n�h�W�|�[���蓐wz#�2�ZKcR�$ػ�ҏ{hݭ���_ؗ���I�]3�og:&_�KQbD���/;=�<����I
h���|\�C�W�����Q� ^��1�O�k;Ә9]�2w�y��2p��b2�d���~�l���@�@˦���p餉�5�	i)�M4��2T�_��		���Hm�էo��N �='A��D� S:_Yq�Jn��?�WW8�,)h�:�}�����L[�8�"!n���a�"ښ���� vrY�����2�x�Ѕ1A�8��}�s��f&��H�&z���.1��Fz���H2��e��-)|~�z����FZ`��?�4��)���Q���7��w�#I{p�H����"D��EYbiB���Q�B��F�n Tp�a���I/���&[
r\�Y���5L]�J��oɒ�`�:����7E��+˞j3rk�U��3�L�-��C�FH�$-�|vT�,�dk�%p��i@�/�[����|��t�e��[g�&�=�f-������z�e�`k�!��ŀ�e�M,�*���O�`AB�a��p���O��7�ل��1h�\-|����L�Ԗ.g(���<J�q�>B��[�~�3�85�Oo'��3���T�@�͙|�ˉ-ܝ�y���ʑ_���8�(9U(�.ҭ丠?}�#E�����#4=i����V_��BFC��-Ή/�>� �����>+���q*�� ����@U��^@�f�ˌk��b�I�Og\s�إ 꾃�TJ5�'U15�#F���k�Y?�@��߄C\�l�,��#Ϝ�����WtT�?�t��6��0 P���B|��m�� �"D�lBg���zi��>�������R���E��`�b�ws]������8�';~`������yU�3Ƅ<�v���S'��H�s���>�ȅ�v�i��,�.���P=��O�
_�;����+@?��Q�Dr�:g�kiUٳ�kD�;���v�'� )����w]S���v��8�^��a>�Qg�'UƊJy�d^O��2�$Z->S�"V���r{�2}�s�j�L �XB��.K�?��+
{�>ꥍ7џ�%^ 8ph-���=�$�����Σ����o<�w=��V2��C�f��Q3�F%�Il�d#;�q*<N�0�+��{l�3��P/�V���L�n�P�i1W�P�)��������ެ~��x!_�ц'�c�f�K]Q�a]�~��)i�����	��͕��[S�M-U�V��].�߻?'ɇf&��2)ȸ�G��^�y�x ��ݶ�HF5P/���w0�5�rj���IR�_k���]�'e�9n�!���D��>Y+�h7�[c:'h�~�3�W�Z��AϠZ@͝^E+&X	mC��S�.��w�Yw�W�<D�v^��	Q.t��5?0���R���[��["�'	[��̜{��gM&�V�6�u��k�:_
j�	D�Uj�sR� �+t0d*i�
+5��b>f+#�٬*��Y��:=�|���C�o	�\�\���G�L��)�FK��Mt�AM� �d��5l�*�%d;��V���>'�'�����%�g�\%�{+D��M��v���$��|���p� �%���"lI- ������D�3�"�' 1��/���Gu�����-�=�Ƽ4x�K�"T�m���u��a�6Bb��bC�uc(H�b�b	�.�ސ���o�)�k�$qf�m�k3��w��R�(x���Tb���8��"�q�C�OC�&�n���<~�"d<����B�t�-?x_fW
��H���g��e�mQ��*2O�����Ї"ʾl��}�����f�IQ�&:�V�&�t�v/��0Y�,a��.�!x�H�A�����[�$�@+,�T�U��C;aVmZ�vg�Ro����&ގ���"���X���Ȉc��@�Ŧ<�v�n�wm��b�L3�!�2S��o�H���.�q��[�o��:~
�(bbY/Kwx�6M�-AM��K�8u؆+p_�cp�ƃs�Xre����o�E.���?t嗸8�290�F\��� �(%n�z�� .	Y�Bu��&�ǛipHٜ �X�A�����A:r���X�p\�!_�5^G�d�G9�wh���$j�{�e���4��N�¾i�ʆ�@w)�"}#ZJ��+�@j�a���1#�
˒�Qa2�q�ٕܮZ��Ӛ~|�w�^��ۢ/$@t�&9)���T2.���5i�;��9���������܅���7?5�����L�ٓ�/��@;�p�"��U��R��׍"U�F��G��ro �#<�ȳ~5�@�S��(�.�(�C9ɨ0g�:��N��
�UP �v���G?R�go-�@�s��c��YRSV:��f_ČR���H�uF��:@�J.�6͸E�趯=��C��M�aH��/�q�"r�-�᣻��"�Ԩ���9e_�+:�$�������r���~ӥ�댃�`��Nx�yX;E�k�!̰�=f��f,�;/�k�=�OG���5,���L|��?�"�$�8׀֨/�����pԉYBʲ����G8Oye�E��L��ɦqa��bk괒bO�X~w`������~Iׁ�H𝕍>�V	���X���^��V�aM?�3	��Z��#�05%�a�6�v`��\v2�T{���!:q�]��}q��r����<̎�.�~Z0�$9����<[�����	�ͽ�w�#�d5^ �� �2��#D7`F�0o�*_ߍ�h�2���ͯ,ip�?Uj)���T���$������H�
�R��+����P�/��c)-�%Ή��@!�==|L�T5�N�?� ����90�\�zP)�9|��!�����Z6��I P��0��u���Z���js�i�Ae�t�0V����L}l3x���<%q������֌&B�^�-�����]s҄�U�'$�M�#���ǿu�q5����	r��j?���5�)�����R�Ə��r������b
�m����1 ��) �A�M+�Y;��2����I,O��>K{�D��"�4�L���D��;�y�4w����vW���3���PǮ6���&���([
1ÁA0I�eh��E�:i}mv��H�.b-�rN�
VI�o�X�Iq<f��cDͳ�$FUxLEA��Җ������\�w��ӈb�E�MT�ߪ&����J�u)o���K
w�L�wE�c�d��{5�֨U��F)�}��J��Ϩ 
��������+�BJm�ڏw�RJ���	�pï��4ְ��NK�&�O������6��o�����WQ�=���	F�ǙKD[	ΐL� �F@Z&�(t�7��&���9����J�n���ͬ��o��3�M�Z=Y��t���<�i1#As�~�%��X6�Uרu���ǒ��Em/��C��ҏ�=�ϛ�d/U���(T�*W��@pO���z��Q!P�l���"+Nzի�]p���[��i"}�*�@�p��=�WK��`F9�t���ɘJ��+�;��]5j1��\;�����pV~��t��]-�R�e�2Ev�q�q����]`��ep�6�5kR#r����'R�U�Z{����Ҙ-�$�a̲V�����L*���7#۳%�5�`�d�&F,bA�����s��GÚ8N �p��6��=�fnW h�S�gv�=)��������k�0֩ڬ˦� �����Fd��nE�E�.7���En���I�R�(P}K�� �+:�@U�f����;�$1�uLFO4��v�mj$a�+�=d��iX��4R�eL�q2�L���@&��W�D�������GKKm�{u��쟧����=_pz�$UD������TCV��`N�����~�X���'=\Y*j$%t�	���T�_b����ꆏ�񻞂���Vk���#5�:��N03z�D�v�^'Z���U��(���w18��=��N�l��ɾD�����Ç�|�f��b���\<*6#�n�Ё�D�+i�͡�d?��/7�Y>r��E�ah��r�'j�ߢD�b�� ܓÜ?�O_�s�wUX�t�T�(+�p���
���*4���@�g:W̪񖄗�qO"V{r7��^ϥF����-�������>be#Q2p����H�ɷ�[x��v��AߔKK������Iʶ���9�c������c"˯7��*0��S��?�t;l}�}�z.��[b�g')@������A�����*��3~	�a��Co31�x��K�!��Z9�1>�0�q@��wm��5Gܨ@I��ow�1��T���>�g�KҔhA_�v�6q�|�3��k���NC��$v�}��+��(�nc��K�__��(w��v�2�� ����^���wNG��2Uc������憤�J�O����bە���ۆ���dc��R��a�Ɲ�&����Q����ƕ�3@����D��O�f���b��C���E�Ѭ�B(`�v�b��*���_i����Pz1�9#G�\���﬷�b��:�n��ߌ���P*�������s�Z���7!���[u�-q�P��{��F��R��{�>|d�����(z� _m���h)D�y�����0P��Oam	ފ4�ᩒ��Jt5E3�O2� �&�}�1�H��j1�k�T|�����t?�֑���]��>�Fo�铈&8�|:�꙳�@eM�L[�h� 2.	���� �Wt�>xR��M��V���A�QN�L�Z��?���� D�z��V�����!��y����6|	:��n����M?�#���̆�?���C�w`���m��?�Q�n|;[������PI��Rt刧u�/����#���\�ڕ&i7MӜ`$m�w'�P�kmυu���9��r�
�*O�?�οo �_C7$u��_�$e14(��� ���"~.���X6�z�W���E�И�XJk�yqq�7n
�.!��>��q�y��ǳm
r՟"{[�9ǁ�ޤ�B˄�+ݡ9*��L�ch�"��)����A�K�hV[|]k,�y�zn�!�#�7ŧٌ�<��B����icB�vc�R�ڍ�q��%d%�)*
a���<��JCܸF���UD�ni�<��-���ɥ!����7���i־[W���Jp/�'�8�~�&ÿ����@W�㵹2tn�H��j�J�
3T0 �-�בl5S��d��E��Y=9k>�)B�� �P���6rޗ@!��B���)�W�G�)o\v~S.Ǜ�� �:n�6�ʀ�2���"(�0>WPg� �仹�7��Ϸ�ܲ	��4��"F$e|���j�2tY	ha%�I�f+$� ��9�(�ZG#ί��*209d�t��M���g���r�H�hu�(~Џ�c��15ő?L��=*��Xwy19]=��6�+eֱ����5�W�d���kc��tÇ��-��"Ȑ�̗Wh3���Ӡ��YK)5R���|�K/�ϣ�=W���)���`�
4�� ��A���;%M�`�,�l�a܁���J��fHy�5l�'k��EݸuGBR����������^/a �|9?�@�M��ig�*��0�0#��Z�����˵��{Ɋ���iXg6;�L�<�UӃ�m&��&	����d�T�p ���u}���E;�w�L5_q�,����<��!t�%m�v���]�#�b��?��J�N�K�з�iyN&��ާ��+����2l`rf"Q��oq���(�#�=�{�X*?t�VNCS��4���i�ж��!U ]�Ҭ���`D<�2�eӄT���#���pj~��mP��,���\��7k����FF�S�x��[I)c6����{x�ۺ���0�����7�������,xq<r`?K��=����ɴ=��mC��w��%�y�H���X�EL�ʠ6?!��q�\����b�6���]�,�.L:a��ՠ�b��x�����opJ(�+��5.p0� 424��y0�[~�@oڱ 壱/3�Ova�p��:�$P�u��K(Vs��P�B�K�K�B�5����Z%�?9��O	�u%c��FG���ܞﲪ��o_I��A (�*U;Q7ᮯ�	[.J����I�ݐ�y�.�H���t-+�c]�*024J�R;8#����{���s�yX �x�`������jvA0���M�i�c�3�%�Nj�"b�n~��|(�a�
�4QP	ԗo8��`Y�c*d����F�?�\9�)g�u��8ܘ'�٦7%�����jݎ�s�Ex��wE��b꼭�g�`T~��'��#��t�˕�iZ�ߒ+W��vMEou� �h��/>x�=�Wֈ^�C	�E!	�����s���kyh�J��-5Q#��IWy��A=���cy����C�R���΀��;�֔�a�h>�!��n��d��QYg3��0�H��[�տ���"�ֲ�E��P����I9�rc]�Q]!�a���
����2��=�&�B�Pf�V�r��h�Q��zp9��;��2F�����Z4�Ӻ�/#�`Ų\��S�X}��`��{�53f7����?wq�m-}r���g�Ul�k��4�����?d@�a+N���;���[��E�<�٥�.��T!��/*.=6�����=��Vh�^�y���y�X�<�Ħ�IT��Ґ���1�5jV����Y��<����4c��m+�lY�I� ���*�l7}(���y�9��Z6�[Qf(� .�+��:�y&N^��j�*�F�h@q; ����K�a�M�j��q#C��/������TA���N wK��OX2�:sB$�`��-�������y�P��)p���WP��
��k7���{�\H�p�^k����.���ʮ�mI�e�r�V�J�� �RMbI0;���y~e��8;w�T+��u�����n�{���3x`P�(�(뢍pZ2�HL�R�Z�B��x����?E�%��<�`}����ۙ�]}�k/�Q��r���*$���)�-�m����r�����4�\$Tt���$���W�0ƀ���ۦtЌ#QdT	�[��)q��nr���>�r
��R.eZ	.�8\az��0BgyGßHKbn�d4ٓK���/��\ax^tM��!M��H���D��`����,q���0�� 	'�'�ِd���,���-Q/�R�DT/���cu����I�cw;'�t�����i�T^0kB-�`�OD&ceI�W��Q؇���⬊DU,��>H��&�w�IaF��lQ{^�0̨�>���Lݡ�|�z� T�@��f�Gh3.�1Cdf}�g�������9��MnD>3��t��e� GD-ˤʬ{���DR�5k��Wm��r������+=�*:j��5A����IL�o��CPxK?{sj�C	��=*�;��ڎB�n������T1GD�B�"ҹj
�}� ����C4��?J�!����4Y��x���rn�Yi���F���-�(].��Y$W|��Ռ2�V��q���!��=�S��W�TؘC��-V�2�q&B���^���
�����@$�`ޑ��:ar���>xx2�Υ��e�'(�C��BZ�٣����Y�|g���%#�_��aۧ�ܟ�צ�}�]�'�:�ʗ�=��"���o8�&���!Y�����y�T(@g`�(ezS��l�hx)�hC_�))?T�	��~M!d|o���0�{nC�a8~�ו�4�7����8�DpK��v�W���2�\һ	����c��c����:=�@{5E�r1�_�J������z�ڎK-6�N����O��vǗU3hʰ��O���Y�Wg
,���mP�@s'r�?t�m�N�#g�������w�	JW^����(��
��5�yz�c+X�V=���p���6��tum���v�#�{�= -�=v9Aؖ���3�m� ȗ�.��`,�|#�me Ⱥ.6�S|SLl�ֺ3��(�EE�,ԧ��ܥ�����ˎ8ͅ�4��I!��_�;Jk�I4;I�׆�ٷ�y^�hg�h'�T�ɇ�Js5�ى4qR���!ԇ�k�t�D|�V���|w*JF�bp�_WF�tH��k�<��E=ț�m��r�5rtL	��h�&�L=���ݎK�.�7�@E��p����U-�vդ�r~y�#����#�=ߢ��=d$���x=����2�;j"�7�w�Hἠ{ ���{������o/�dj�} �f,�n��iٽ���2�6�Gөu���y���Gt��14=v�r�����Q�����{ñ7�a����b�`O����~���QS�\����tʭ�_x)��YYUIXi�݉g����;z3
�S����˿�pUu�}�TΝL�LF&�e�����W깪X=��8W��殛�P������bS+Y)��p����m�N��٭9�XnG*d�㦇|TP?�Gh-?�!h+��`�dz*@��^�y,�E�ۂ)v
�\i9IYz��=����8m0��w�\��i�E�_0��=�=�T|�ӄ�rL|3O�r�yi���r����0�a�W�]��_��@���3���c�}|~nH�d���ӳ�s<jKS�T�7�� �9bf�?�~�@]EF<9,�LV�aY��bFМUJ�~��֟fԩ�V�>n}j_�1ƣY��5l�1c�e�U�D�|~x�Ln �n�ߤ�������,';��A�`]���*�]�.~�N���Ȉ@sD��`�#��������x0>��Q� ���Q�
�Ĝnm��+��c�۫o)3��d$��-dR����O����6�\Y�K���&.����?�-[la���PW�#ʃ�={��m�
|��S��ݴX;���Q�Qfv�pc}��q��XcG ;9��'ǝC��Y���h�6Ľ�2A���I�|R��	�AP������=�����Z��'I�N��On_���A\���&��R�|-R�+�m�R����=���N�R�.� t0V 
�e�:7��+k:{Ա��(D�q�Ϫ=�Cu��<�QOa҇��B[�;J�C�I�����9j�����5������:�5T)��2�x^ۍ��c�ή��Vn��K��d����^h;v�F:�;z��5�,��w�x���}k9P�E� q�Je10Dpv#t���TX�|i����>��}��xڌ׎��z���}��f?X�4���&�����/n��0F|OB&�mh�ZF��y�G�p"Xt����[�u�;!��3�f�0��4T�u����ȁ~kl���$6�V�j�ӰR��򰰇C\���ڕ^ļW�v�&x�a�S�5�ؒ��$߃FӰp������,]w<Ց!����>�Lfi�/�V?�c��)LxET lίh�b�W�ӝU���R��"�ˁI{���Qb�8����t����y/X�M��r�Lؾ�pͷFYi��A@�	�o{U��bश9�~�k�aO͕R���d��Ϡ��@{v� & ~x^�ضQ�v�n¦P��>tȉ�!���1b`�-=����N�Q�E�� �y 䪷���"�g����|�B$E����kK�"k�9�k7驷�N�R�@f9R���UcS����5����SO+A���틙�_;ug^J�T+����3@1��
�#�=��W�v�_zY��}]`�5���Ըh!\,�-�-&��UN-o��xG�g��^�9�˅Q���2��B�\����'���V��:�bԡ�<	 ��~�����`��k���+�F�Hq)^?���ט�<P�����J���׃~��#��*�X��C,��)8�1ƣK��тx�4�*Z�s�Vt��7��4v����dy�(0��4�hE�y�zy$�&�{<�XX����t�|͝�׎�˔�@�gT1���Z�*Ry�hTl�|���=cvG�K���R��{5�������������=>�e���n�4ּA$e�|� ��d�Q��
}���g�빦\�ri��8��UbL�����v�_�j'|����n��=��#S�ǲ�n�j
lt�9Ns�Ɯ�]�{�+y,d/{]-�v�!\R���6oU��z7���g��4�]�u��#;�^ڜvGZ���(@�" �gc�#���7@0��&���2����KTް!o��F� ��
���@)u3nx''u�l{��a,=�D�h���2-lT��<�p���7��A�n�ENʁ�U����3/�1x��i�;5�3��h��-�iYF�H:=��%�|��V[�r�e��.�<~C^b����z@P�!ώ�wH n���q��\P�La��W��vu��(�6&�51g�1�E��l;�aп)�|W��IA���ji�S��o��uV.�K��1�����ᙀ-�U��y���$�$�/r]5��|�r�ۑ�IX�)Y/�UPLn&V�4~ޞq��E���N]�H�FA �][x��s�>�,�zɸU_�v�4�&99gA�xr�r�eҍ	��뻥"p�Wgr�5�è��~D�G���Z�ec�'�16�J�� ��*��Ls�,�#����R�0�[���u$Q��m�"���!��Sl2���(3hC���x��	.}7���߄n�$�����EY�))���_u�hm�ح/���r1�1��ʰ{���m�P6�njk'@��.dǟT�Pe�de�͊�p�t(�F�>�RT���|"o�U������*,��2^�9�Sx�y�W����u��wd�.g�4��W��:F{�.u-�AJ1;��)E3m���_GOC�=�󷳥<��"l4�M��Q�a�{�=�KT��
X_X]W
|�" �k=ͻ]��6-ݐ�f����9�Q���c���3��{�N�Y�l�F�-��],��ZP�1�ל����λ�^��������t��b�!���0���w��! 0�B)���iL��09W{�5&�H�ܽ�E�Bb���1��w��" ���:D�ˬ?\}�B�TH~�sW^��y���x�����D>��&B�=6��� �ˤi1˱C���/��=�o�Ϊ�9��/�]�e'm���铁�>��2Օ)!£.�u2�K�E�	x���B�1Gڷ�o9Q�t_O&q�,&���Շ ��#�ڔ���=�&$}eG��Y��D׷-M}�QG<&��u5r�NI����.����w(�q�����:���������y��O�+�dD[�/<�x���6Y,���9~����%��f��+����i�u�Cm=��k}��7�����ֽۿ�����ϯ3�)b=�$���*�5Y�橂���
	�`܁�pR�I=Z���) �~F�5*�
�^�9���	D9y �k�)��9�B�-XU�B-C��4#�L���1�Iص�,��Q�R�Tp� %\���b�)�K"����<Oa��ׄ��ӳ�1�"�<]���������h9	���٫#��D��F�P��CI��-��ƥ���h)3�$���?W��O����	v/R?��S�����0L�A~��*S`�!���W��_�'_�o���j�m�w3�2��v����tf�@Z�c�����uސޖʺ� ���2+;�)Y�۵5�+��6�%�:1�U��I��� �������a�wWA�:T��q�t=ϥgr�G�4���㫞���i��`��4�~-V�y�"^��[�s��mqu#�2�42��ti������-8���GgUgȱ*�����r�N9�Ar��nm����"���U����F88�Y�{�h�|x��P�IU��E�+R03�T�M`q��������z:��yxX�F\��%���?|�|p��є�_@������ҧ�,�i��s���3;ۚ��vK�oi ���\x��?>��uȈ�h7i�:�/u+��y�G���o�2�_Y'q��������X&ҢF��S����ކ�on��]��	��$,YǸi�X�S&����������ʏ�ӵ+i'����Ț�$�ɪ�Ψ�Y&	j_:غ��b-�A#[�0��,`[A�x�`mr����kz�E���6�d�g�Ch��E���D�B��q�W;�G�����ѿS��r�J��������T8�%��fn#f�EC8��{�l_;�[��Q��n[~�	I�o���-x	t<(٧x��I=ҫl&�Kx�%(��	�Yf�7gH\i�Ď"�lh��@�`YpX��$E�P�"�z��X��9�#P�X�3��BL�B��U`3�1}����S���Y̺_����3]�@ �&?SP�aq(7Z�]��3�y�=��`�\3�\c 1��+i�:���=���" �)�����>x�}�瀤�t\X�(_�.��ꌺ�������	:�,dR��K�����i��-G��@kQ����+����D�m��c��ѕ��Lֺgh��[Q�QgD�U��.�.M#������� ��]�#Bn*E�a1�9���@�
�"E�0�S��]����D������/�0Š�q̭��IU���]��r~���
p��80Z>�^�/9"��z'E���MŐB���!o�J?T�Q/��%�R�h
������\��X��c�O��ww���q���Vf�aS�yQJ}_���DRG�N
|e/CP�?l�}V����Y\EWDL�g�W���فi�޴Ԯ�Y�K�/ڢ+��"����vq�7uJ�b}��Ez����X�5�YxT%�^@D6�%}"�x�z�	�
�`_EJ$� [�+�w]��X���*���2�1Y�����`w�d̈́�C{-��8���Q�1q��$9!�A��a4��)%XzH�j%gݥ0S�e�Dt���4�f[V�r�v��T�������1t�y9��9���� ��
)K�E�����AY X�n�c<ısu8~��BII�leMIʔ�N��_#��*�[�{9!�H�*Q�J��K��-I���$;���y_.���o�ܯPG��s�������Ʒ7� �G�e��dgma�C=#q�ꡑR*��fI�h�S��
3�w�C��Q�m���T�u&
�N��H���c~U��"[���} �6E4k`gx��E�NZE|�d�2*��T��{���Nq�ACe��<�9j�C�^,W<�Ђ�^v���Φcp�� ���ھ��S��X��ךԅ��qU�;z�23�=�ڎ���ӳ^F��nc��z��n�}[�.�\7��~
�����̫OY{��!�M4H��J��gBU{u�#~�M;F<����'j�^�Г�]'ReN[1��������
�X��ߍ}%%u�,X�~݊����7�v��@F<��?���խ7>�%�Z��<u�E��j0�kH�d<���Yj�/Bj�-6��V�fEh�hd����i���-��g�(���{�O�Av�FJ�1x��%m�f��4�)�%/��n�c���U!���ήT���u]��l뾅&��5C�;XZ��y��)�8��;u��P��A��
:$ޏY�ak§�1F%4��(��y�$�Ә�QE�蓢%;�K١����^�9���>!�%z�/~r���yv��I5?I۞�Z���&u��Y�߰՝ciR�?�
wtU(�	O�C��ȳ�3���-�
ÈR/](!A���=������������#���|�M9���nY�(5��m� ���{3�H�Ti_���ŝ���6�1&e�����G�$�s<EDaa�b�g����{"爱���3ۺ����W��5�&ݩ)��L�y��{6��Ս�
�Q�L���'k�&��*~�X���]l�ĳ��٪:�?�	�
3a�yk�L9�X�>̙bUhc�IeJ?����&�+/��9��2>�u9�65B,��ؽ��D��.�L��%�� �2}U�����>(éa	��u��rJ�0֎W .�-J��2�91����pX[wl�[LA�E+Ğs��w��`Λ�~RO]P��K�!�Ű���	K�2o�O �*��L��<$�B���l��%�LZ8bD����=���gC��$y�P
┴� ��U�˺2�\�*�'�<zO{n��L�~�ֻh81�zʾ�!��(��{G�J�hC�j�jr��dc�d]��r�ݔx��k�m& 5$b� ��1��>���9�̹̤~@�k+n�TʔN?�Ѹ)z��C/�6��R*����W:9�(3��2����=�����CMWzK�PF��\[�4��]CC��Ǝ]�q���xNNw 1������T��DL�	<'��0�3��`�cƚo�H��r�}u�[Va�F�o�:*Y��iĭ8L�u�!⇓'�X���Y�5>�S��S�����N6f*m+��95�6�M��g3�Z�G~GA~P�P�=m��K{�����ڏ�[[�W�H،�IVc��$�ta����n@��52
��d{@�9l����Ƅ�9b�ɡi����J�H��*�[�#Z�O��Å�w�,?y�+A��SKt4F?��xԜc�$�c� ���z���x�I�K��%��HuU-��!����,I0D��#�ƈ�[ 1m@�OZٌJ�F�&g����|t�`�xk����y�n��0^I��%v�mY�����z���"[��]�8�-9�H[N]�:�qJ_n��t����-�O��۶c -?����=�>����ǭPe�������;)2}����4�qO	~�!	�촂�2T��y���Jc�9� �	��<�ʫ^�Y���O(����7��%N���'�Xw�����3�k҈AF��\ï�
*���:~,,��vˏ��_��r����
���;���e��Dw���
����R��{�WO���Q%��=�N&�aO�j�p?���� c�q�a�<�F?Fg��P�l�����)���z���IMe�����"b�&���h�'+�|i�TД��x�M���Ft����2�Qx�TZ��)�H<`=v/6ܤ�� }/�:؅�2d'M2l��q� *�!��P�t��h{��槥�2�ݓf	g�?�.�V�K���<�N
�|���C�.��~M@��փ��Έ������^���u $�
Т�J"?�5k����z�����W���h�>�~)��R)����[g��ߏ$�K�K@9�4u Óz7"�Hj��9��+@��1Y��6�y����`Sα@�OB�^[����T��I��6L�Wl5��+��j5�ؤ�Ɨ�)d0�@����>y/�OQ�io�'�%�YI�$�jo��B�~hP�L�����O�����,A�U�]�v��~���
	M�+�ɾx�gи��d��,��쾝�&����a��e�"���Vy��u�"����i87�m�J��61�J����!qC1�m��Zv����h�˺%��{I��3��b1���5�L�������2�/����g�����R�87�ȫ�`�Rg�@�t�>;Rp��<�Ty� W*̑n`�i��!Ɏv��3���<�a�a�jV3�oZ9���Q�7"�{��j�n�$9hה��Tb��8�#X�z����������r��y��d��^�,י���M��6�MXDV��Q��G�F{^5~0��O�j)��^��9���5����"�](�P������/�60�w-�O�G���,i<+����+{[̐�-�9P;Q"�DŁ�$P��䛇�q�А�s1���m���o�|p�9�F����N_��\9��O�