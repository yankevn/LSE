��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?��O?!��$v�X*�y)�ޔ�$�m���o~kG{��cn�B2��d�f_~:���f&n�d"j�i�5�Ų�x�����U��*��]a��
5i�&����Ջ`�ɿ�0�0H��9���D�P04��M��b�/hrxD��%�:��xd������X܆��7Pk���I3�BB��OZ�m�S�E��kzw�
̗��8�C[S��a����;u��شJ$4)���>��Y�,?+��M��n������v��n���}Z�\/���.�Q���dux�U��L�<��	�F"�K����u�4`�����d?�zH���֔Q���ŭy���ֲ�l���3a|�7��ZӾO��c^yr��j�&B���W���>���G�F{���\Z���S�PX3�L��]b$��U�oy�����?�!%�c�?���_H��JgJ�jG] [q��8����*i�ld%���_�vX��,C������gl�ZH"׹-���I�O�n �FQ2ݠ�O��w�xn�nΕ�n�Ӯ#��7.��F�~z,[����⼴F��e��M��"z>t��c�1�����󌿿��$@��?X�j�7���p�ok����ö�Bl�UŊ����+��jR�{k�O܈���V�E!Sk����l�c�h�z[%f&�*קP;�����v�br��S'�}q�ZSm,s�$�0��7e���6ɽ��էq8�4�Yځo=*pH�Ӿ8C���B ���k�ˤ8V{��A��WDn���ϰ�#)�k��� ˦��O[�d~O��w�;*���JVv1�]UB� �0���J�/s�Umf,�Y�B������D:�l�5$�=���������RL�8]I��v��s�F1�6>�/͏���C��TH�5��#F�:�|�E�1��y��%��(T�*��˫��b��%
���7S73D���+s)Le-�m��?�����p�{^�]g̙�,pW���?���ߡ(Q���3]�j���.�m����✦�Y�%����Bn��56�u1��g��N���2���G�y���s���~9r���+7�<Y�
�qWٹ!^Z��pL����xDn޴�PQ͞��o@��E���������8�������S��$?İ@�Ϊ�M)fރ�m,`�	�F�,j�{�J$�d}e�gv-Q��$Jh�"�Z�����>!_"(c��_�/Hh&�HAD*����i��*���5�����h1Њ��Qf�2��Ԥ����8�O�ғ.�J�<w!�kR)���e�yfK����W��p?����
�hi�	�k�dޟ,�qiUJ��ؿ}ʇoa��]}��6[���F�0Sz���އ)'�hC��X|�]-*��q~�;��W�^{�RIq^�_g��֝�M.r��"��<'~C�`���R�`�� Ț��LXS.�̯)<WO��V��P��6Ky�gv�#�V}�;0�|��V�mg}��ɯ����)���@s2��o��D��<S +<S��"���ҿ��k���3�Ī��8�X�.p�$�'!EU,
u���4�>��U�
�5��� D��ܼ	�Ȟx��r$s�R�"�⪈�j��\����U�v��
Up������)��(Z�U$֥%CԦF��#���Y��(��d��9��߰P�O��\�Q���c(TJd=��"'~�`><P�M�ޔ�!Pb �b��³��뜓��Z�7Ȣi5��Va�c��o�-��KLy��믉�J����7u!^u�Om{K9�.�{���8m9�*��/���I&��%;#�*�=�n�|z5S�g)(�� �J�����'r�5?ø�׬pbE$�H��h@���Z�ˤ᤮��ޟq4��~�H0�!��@c�ֲ�<��~���E%Jxn�ܫ:�`�Ra���G_(S#���H�U���oSDJ�_fު�C�����;ˈ��Q��dBFm4D5W���]$�����JV�c�Jyr�N�>]��6�`pq�g͝����a'��`�c��=�J�o��R�@�D�I��B|��ǉ/ٲ��ɨ��h�|z]�̴���{�*f��Hg{w�M�����TƝK0�Ѻ����%i�ҥ�c]�5�"�l�Rn���������$��*@t��['� �xM�V8+�46dK�|����G���9���jHO�N\`��*�55Mz�}���4 ��θ����|�
�R���;.�b�S���k���|�V$\��r$'I�ÏC.�V�sӳqnX�Btm�e�����N���%�K�:j(�1)���8%���qFx�U\�������s��؇������/�3B?�ˣ�=)�����B���	����;K��
�#�O�W7�A�"w%U��7!']�]����k�v��F��$�/G�-��2���O_f8g�6yzGr3��i���J�z�hjf�G����4��=!eo�q]��p�z�յ�0�eF�s�i�c�ۢ�3� �������|�t��؇�eR�>ތ�c���hsO��?uZ�L�5a>}�8%��T��E�u�(H$�\�D�8�(�w���S7JV~�k@�kf�^�U
��q�J���7�g��aDx"�>/��>�~�NR�}�T쟚�흧��o���C��qJ�!��%����������E���\?�S����
}�Gsw�q�]��%-�d';�:�mjk9���',����?�g��T��Sm��̷�Lj(�@��}�T�����̏�	
�~ �]p�UE���m����Ge����j�X=%�ȗ��K�}�01��V�I�Z@�O�C�H�����Tr=$�կ����+_���&Bs2p+vԚ��&ɭ�T1�a�EI����a?q��t7���gη#�fv0ދ0�������ȸ@1���=����^
�}�u�x����Jq�e���^�:��1�ý(� eQOΕ:�ZPkx���~z2o/��M���xAݦ�6�(Ao:�I�E x�#Ƙgh�eg�n�$���:��Hq�/#�8���p��}����������&�2�&���f�H̆��ձ�O&&ad~NE?$@_�D@\�M2-b
Pt�> jy} �<��4f6,=�ƅjc�3�f��A�mS6I��wB�T*�=���{��0ўr�*��Xȴa����Mr����0�b�zH�T��cr�ly��7�ߟ��`;�c���z#�y�ޛ����L����*~��]k�M�� �{�/lx_<���Q4��!b&�1O3M��b`FH��6F֟?�C���:��i�߅��&l|�b�$�X�M���C���Y�V�5�����_IA�4�ʹ�e~)< C��!�����8�3-FJ��T�pe��B�b��_�2׍wV֍�@^�	�!��4�ܑ�R<��zC�Oc������mD��[9�Afˀ��O���8�Q�_�mG��ğT�2�{�� ����$8�ODh��Ჳ���A|����Q�Ч�O�πU���_���:N���3d��mʺ�c%��	�����\�m/z��\T�o<�@p��'�s���}�Mov�� S|r�+��߽�jn6R����#��$���2��E2�Ƭ�_f�Z��Rm�*�fGk�����LU�����*yʩ�+�[!��3�Q�d��	���Yp�'YlUy�_?J�G���)�ق�#Z�J9�N�? 5CW�X7x��!)w��ݵ�9)���C�<������c\A�a{@����`��9Q3A��oI�ͩf��"�Y���~���ކ���xK���9��۷+ތ���u��?���򨖷������$:h/<��`���ɯWs+��+��Z0�
k�����ߢ
����>{���L�V.����4/��w��
���>7�oQ,u��X[�����k���7%�.P��ľy]�c�ߤV4w ϲ��B{/=7M<�k;�&1�,�50Jq����~��zgl�s�ZB0~}@�O���+��	���4:��\�a�D	CC[�J����g���G������O͊�p��8��l�yF5��i�:�}��=7�Jg�d;���!{����������,�2�a̾F�����h\BS"��k��*h���'�MR3ZxMΦ1)��KF��sI`up _�K�*F�#�qd*��p��e}�u�]�
���&0M�BnR1{��bQ����"�iv�{}�~�T͉�VUKLuT'
��4h�5	�@�ϸ�V��
�vE9�-_���T!����э۬d�
2��ތ�8[�����w �"!�8�i�IW�q�r��s<*:��{��xm�е%�9��Í�������'��	N`4�����Zj�g��TUN�rC��Xy�Sj�F�Q&:y����8Y��qN���/�L�ϼ�S"btdD�?#w�r�h|5���ɥK��l��.XY��T��9k�C/k!�&��3X��q$�.5��l|�!�ս>oa;�*<�o7��25�6��u��H��X�vDƖ��G�������/���<	F��&�c����t�ڱ\FYȲ��RpX�"��+��J����F��W[?}��X@I��L9�M��p��w����{�#s�N�y�!;�"�O���( 5�c�<��Q�s���('�IG��70�T�Z���w�1����/b�$��qn��w�!���@��=�4���dr��ُ��=��v�(��o*�7��LF��so��ρ�LqN��&�ph�13��c^lԆ��VMցPc��x�.R�p��F�v��5����x����!; �&]�i�4��^G��,�<�
PE��� C��Ky�]B�����f�D���=ʉ�ú�Zi"��w��)���K�δ�d����:_�Eۖ��Gp�+�����ȕ٩��Z0 �G�E��
����U9�pa-b�x&gT~�3f�X?d1.A��$f�W�d.HK.��0�����}_�ZIT0��h|���3� xW��/H'���.��`�c�0A�=a���ČE�O�	W��2e��5�O�k���L?x��4:~+׍���d�Ϋg�I:��1�]Qނ!�L�K��M�#��B��wg�΋4XS���ϋ��t��S� ���F�-�Mn���T�{&� p�Y���8������ӡ�y�?�[����	�.
�JP���1�b��4Q�:RE5�K$iA���!�Ll��+/���wpp���� E��U,7�,��l8\�0oe�Xs:.oJ�&j�.���5$T>%<�&���HTn,��+.�4*��V繧z^����B����j(��->J�B�7�mH@b�`�G���֢)�vW�JY�-_h��T|�QO���/�D`����X������]aA?��M2A��О"怒G�Nr�� �nw>�زG�����*z�+n�~�+���6xXΰ�{Il�cN�X�Ta���Κ}��9?Q G���Ax��Sa l�*��y��R����Xd'���:}�����U7o&G�#h���~�bװ;|}G'�71���0in�D
P#�!��3��|v� <��397�����ܼ&�������H���!���!Ъe���M��e���w�u�omyW�[W�dJ�&�__5G�EQIr�t�}̒���8��� f�߆���
V'�o���V��ZC{^[�n^��:Iy'C��F�ͷW� ��lTY�:I'^��fG1?V�h�����F*_���Pb$I<z"ǃ����S�i�2��
/t�n���h݉Qd
�kB:Ԇ�	4D���Yƥ�RE�jv�_��7��Co�{s�_`��JPE�07ԿTF�s��p��w%~D
��3��W�|� ��U�Y�}ݷ'e��E�g�� �ї=�ܩ_�ʎ�*��Vȍj�=U�C�I�t.9΋3c��M���ɞB���^Y�;=5ٿ}�"e�J��>��j��V`PY������W$R�;|�׳pV���^�}�,M� ^"��?\?��d�RN�y�sXF:�;�~��nXȄ��]�v�?6 �����J��=R��]##vle5K��Xli0��i�ov�BGT=��V�J�ժ�
�Y,���k}��bD/=���E��p�!�O��!$�şO�q� �x��ߞ�:ӄD�z@�k�[{t_��sA�Fj��͘��;_%�u���rTq�PL�^�?���Q(ا#���ڦ��˗l�^����������&{�KI��V������.r��ְ�ir�Y��qB�mT�#}�ҺxVOZרpgdĬ�D{��S�M�����]D��$����M��.L�ޜd�G&��>A��B�d���U��� �0��b˫AY�E�jԭ���1r*���z�0�A�F�^ؙ�<uOT��5w��oB|�&[����h���\
jȽ�n��/��JQW��v�:v.��I�頶l����=6��:��Q��ܺ��@��h ��.
)������B7%���[VfDO�@a.�h�_���s�M̄����3T;4����Ƶr�:&�h��.�{�~+���w�+5�RҦ?c��`�����3��C���\�؁%��j+Ʈ��(1J�6�ˠTx�����qU����7�[���iЗ�>Pny���g�8���R��j{�4o���Z	ôg����p�`���&y�ʽ}J���+�9	���� S�:�n��#!"SUt�@K%h��a�{�U��޽�r+U�A�b�my�B\�&���>�����.��0�4�;6ג$�	~ 7-}�42�A@�T4��6��>���\׏Z�S��V�A�r	b�$��1"2���:1�
޲���W�THo�����O�B�.j�e-FIN"gd���$dp��>�R���@M�wb�ښ8&���B��k�M,̩��(�_p���g�Q�\�P��WWy�4���E�N_뽄_�G?e&�dm�h%_y��T��_�V���Q{�f���@K:�:�O췣�K�N��
��';���E)����$�s|���^�Aucl,t�u[2�%l I�G�\`d�_\m�k�)}��,�^�p����~N���.�Ipfk-HX�WJSbF�*R�;��w��TTP(FW#��W���E�{ ���*x]�]�z��>�[��QNU�V�L���Y���şV��p�-�M[g�4�?�տ��|8��5R��w%�x-�>)�9�m�"$*h������}��9Q߭���]�.�0�@�*3# �����!K�ױ?^�����&�A�)�Kq��2D��4�5�W�f��)������w%��J{ᕩ�h��g����M�iQ͇G��+	'�V�ed�}����Z����[���|Ʉy�t�f"!=KaP����0������-�/����	T�v���O*�19F`���vS*�[�7]��8��5�\����F��Or�����׿�j��,N �/�#ۧ��̜p�y�М~�͉�xH��x�fL�&F��GS����,� ��,�)oG�fw�<��[�w��Wv�X�����@@.��Q@�*��8!�U'-Ҹ�@*<FWq�F2�?$I������^I7�~����c�$�Iq]k���,ƾ$74���	$��c8��6������IŊ���)�NB��JU��R����?�{=���vz����I�TdD�"S��#�7o�)�.��K}���ޖ�a0ǥ��+]��##�&RG��#��L*-��l(�O���`�!Ϡn<(0�ċZd*�`���
�ZU�.���]³�";�����VM��PsZ��Y�W=�sMMgf&(S z�
�'m]^'C;��͛�I%��f̲%��_ė�b�"!���Rekq3�BQ��ۯ�&��DW	v���H����3��͠��Y%�0����~�C�&�n'�U��ҏ�է`�j��S:�*�Hg�����u��Xd7?iU|hj�s�v��X��I\�Br�x���V�&Dj�p��
&�LiyBH-��<����Nw�B�J��CH�����t+q���b�U���pg��O?��\�"k~�A�t���3�x2(^r�f�%�J�k�y2-H�%ug�
gd!"�Y��X�����1��0@LZ�<B�|T��ΎU`�E>�L���1W�lG�q�z��h7��8�K{p�=���Z�����ݖ�B2�u�MV�A}T;Jo,�������N��@�R�	�uQǕlDLJ��I�`,n�k�`(��w|�̖�7�� �o{��Ƿ��'��o1_B�u}�3M���P	㙔���S�[��e��\�z�O�2�����p��Y|/�>����7�m-/�j?�CU�X9	���F�.��g����7d:��!P�����WC��cc�S����Zo��@�ȼ�]Io �wX� ь�k,<O`�����x�>��5U��'r��_��+T}�z���}s���#u�޽�=��;����ꪗ'����iY<_�oh\�X�'m`��Yr�{G���O�����r�����kqK�|��J#��ѩW(�&��KJ�L"�/��� ��J��5W�7 ��`33�J��!y�ù�W�f6k}�h�����,�p���j�n�XyӾI�p��{�L��(8�������8y�P	=MH��ܴ+��k�����dyl:�@�aI\ ����?���DXl1��n��l���f�F[+��16&�ľ8`qWd0�_E�!�F�`���^@q�QS�w�`�4�+���}}��oL�'3k� C\�;֍���Y�]l�����S��� �R,.�rP�*���j���Tɬ���M`�D����='9C���u��d��t���r�1抍��ف�K���d[*C���l�j-�Q�p2�&곤ڒLL!0C��Ŷ�/w�]A]������}����Qs���OR�?~���N���s�����\x�4Fˊ���l�o��\���N�8ˏm��~�)樈�ܩ��%}N�ϕ�����_���p�/L�|5���Ӡ�&W���(�1���O�R:Z�o�QP�c��\��Rq�/Q��v��l'2�R.1�������e�J��)���ʨB��@G})19�Ҋ���/��L�h�Qↈ��rSN��Rm.����"�/��rCX�xO9G��\fph�ut>�̭��
�5�������YV��H�S,�s��s�\��tg�[;����*�2�h�@�z��no�ٓ��5m/R��)�e��Z�CJ 6���;�=R20xQ-��.<fD��r Y�E���10���魩 ���,��#O[5���CC��T�ݧA6DژNa]U��G �6�`ҽd3!�)�Z�V���%���m���'�[��H[��#Z�Tv���̼�I1CT�F!)�����I�K 26r��{�b&~B�-�DURE4Py��5������W��J�9vIv��}�Jہ��b�yi	��f,,���i�hc���oG��kh���D���Lx"x�z�G��y�N`�[JP�DH�ۇUIV6D�wgXu	���>���q��Զ����=#��>60$�����=5�*r;���k�m��E���潽�=�(���G7?������f�%��\�*L[��& �^N�e���|/��@m|�&pG�X
������ݰ�Ss��I<�}�8�N�P�`��I�{����l���)A����Ep��`�jh 6'.;����<�:���Dp4]�Л���*.s�����,�Q4-ײl��Ԙ��`�h4`�iE*�ﶁ�t}��V�:	=^TRx��R�/0��8�$7��4���C}�<ȗA[���u�;�>���(5���cl#~!���t��6)����w�`^z�����£#fs���x�D VD�����~� ����ϣ�eU���A�*�T�
ؔ����<"��ދ�ܪ�`� ��r ڽ����[4?��&t����z^�������G�~V��AM�~o;{���NUMb>sşhÍN"�uX�k�]����]:�|;�B�����C��[J	��E�UmR�b�jSl���I	�\�Ơ�2, �eѓJ!qJ�Xt_�'A&i�^i�SƟ��-p) 7�'ͦz��1x�c#l�ˠ�#���r�NQRŐ�Ό[�aV�� �q�I/Hz����Q�{3ƃ|t�T���eEK�6|Y�<`o��þ���	��W6;����Fb�z�M� ]�FH��Pk��J��˶�.�Q'v4U�͆�����k,�^.�ݵ��	R���}�b�E���Ĳ����?%9gY��Wq$�|���)Q�A\��� �ɐ$�;�*(\��RSkk������?sw͂���Zo�jn5�0cDlH���@�V���-�vZ�-�J2���_}?x"lȟ�T�gN��w.�h2h�Nܲ/�B�3�@�y���{V�n���a��ng��98I�R���U�����3I4Ι�j���ÿ��-}���6Bw��Y�"*��8#����:����Հ�)�fDX���IA�<�(q�Z�-g�%�ݙ�8d��%e��E��)���O"����p��w~(t�6d�Ӊb�1~��'j�7�Ӛq��������"ї _����`xɜW��oT�a��<����O��Iv���4r�q&8�jd�*�uJ_�8_� N�@S�,��k��|D�%� �x�Ou۟Sˑ�"|��5~�*h�u0�<���L�t.۰%���|!���[��bh��@�Hq,q�rsx0�!2ژXa<E8�u�y����J��7�|"�����SAd����2�P���F��%����a >ƿYh`�k �s�RGY�=�;{i
�[$t\��ڼd��i�U�~�[�W3츄��DV�dk�>�d��+Fp
�%%����#3�G�c���d�ǃ���Q;�"i��S-��j=ں���.E����&H�"�?�;d�b��q��8➽�h����AϸC����7_U�M�Z�n�.b�|inE�@�:�L}�/)�>{В���E�㢓��dKX���Y�*蠯*�V���øz#�("@q����8MZ9���3 �j/v���M!Q�"���H%tϢ�c�$:S��T� �KP��k�Y�s�]zԲt���*�S�k�$������x�ǖ5�:ȝ������+5K���\Ue�E ��k3�r��" ��X�.y3�]���}@:ݕ���\P�)�5 ?F��Q^_މMC��'���Ad�`T�枴�����Ӊ���V�u��:����a���RVY
L\�G߲4�AtRXX�Z��fA��x�H�t������:�fŒ��|���A%�2$��=k
Q|��Z��\�QFi��y'2!�uDw��R)Oj1y�6�����ތ@����!�R��]�c����b$�z2�����D�6��)��E�w�3���{hT8���^H�\@0���5��!c*�')��fM�Ke�M��	�Úg|ؿ$�u���˟�pC�C���������Nخ��(�N���n���vw���U�s���M���aM����_�ϙ��b�B�X����J��"Ƿ&�O�ԧ"��[�=V�3�{�
�12eM�:R�]��w��K?�sr�|^��^���(��y�����=(�}����a�$������7�`8?|`1?:"L��|��C֘�-��N!-��y�����D��]܋+9�V<�pc��K�c�a�tH�8�
�[��? �������@-J�6��H�N�{�rv��o2�rz6T���C(���;/G�5A(wF9��,��Y*O�p&�3�[� ������
���vٌ�V����X���	�zw�+]*��]~w��96�Fh䅯���*��O��-\�zt�:�Zj5�ye�xd��XEA%���3��6�@�é/�ao��\��ftsS�����%�4�p��kC08-�PN���`�jȏ
K��Q�Λ�NS#["f���!&PEG\Fwnk,��J�\S��H��e�o@���R�Պ��B�T�<`�KWgX)�S��Ea��h��0ɫ��r����P��P�`��%�����4[>9
@�p�A�#��|8 Y׎v"M���N�s�e������:8�yӔ<��%���}O"�����s3��8��3���Tu��R��\�����L�η Ȳ՟7��� ����U�\����xFs	��&����*$�[��Hȋl�{��D���ċ����,�v}�nu��	�85�3Un���ub����I��Z��c�{'��4�f�E�f�����\xV_���l93M6E��|�N����!0z�Di����;���G&�ıi}��[��~�h�rɅ�As;�p@��	��V����L�7QN6kXJL��7)�6�g5A<����<�F���A'��<�����SF����yA�BC\�)m�kt̕��$�5�>o�c��~����:��������|�nn��w�"�8g��L�f�@c䜕�g�{ڒT0�V�!Ը�|8�A��/6zvTF�x8f�6�/q�n���{��=�()�
�nZS�;�j�g���"����< ���_�p3���C���d��c�wv٤j���U(2Ъr�N7: �H*��zÅY��S g5VܣI��7-+y��6K�w��F)ףr����R�%z<M�`d�.{�\��B�Y��!��ƅ,�Uo3�p�d�pZ"φR;|��h(���R�������(�h5�đ������j$�I�f~�^�Ol��l���өQ�ד�!n0�-�#;���ܩ�������?��m0�uB��A�DgǷ�� |�,���V�Ҭ�l0�@������&���	�Ϲ�z�,�E2R�d�WX��R�DV߶ʰ��t��Rr7 ҕ����v��e���<�J�J�l�^����	�2Z��5���X 
 p�p�8[�Y��K��h�S��|��c�bJ����F��Q���ZW�@v/�T�\�5��}|�zZ����u i5���ԻP:���	���>����XXQ�� 1 �@�gm��?�� N���˔����k����
N���H�4������A����0�x�3僆�?hZ7�@GR�>�:��xRh��e=�⁻�ɒ��'����M%'�8k���xT�^4����g�PCP�FH�P�CPh���}�9���l{��������g?9�z�F����~��S.63Z@��&%�$�yZ��t�ծ|m��/�7��r�� �� ]R����wV�;�j�ǉV�'T���+�fO��w�0׈�2�뤊���B�g$!�7C�Ѵ�HG��\�<�p�Q��6}�2����Gv�y�hF�S�_%�c���Q~�e�x�~	3S��n/$/�fPk|�u�s'�K�Uب�'��ZP#j*�x�.x�pa�>{�(�Y���g4-��N��b�:]�b�O��l]@+u
�����ւ�;kɴ�4D�Uu�c�fd�(�'5�5W�Nv:1�����~�る��J&�]uǳ~ژ�j[-E�J���[��p&a,�@y��`
K��g�����WZZK�f7{�G�܇�&�2�����(C��)@hS�]�Уҡ?L����*?o̗{u�u�-���ogҞ&�t��4�/?�y���x1��z[\��zx�U8��<F�K<����\�e�4C��#���jL# �:y��{��D+a�#����r���%IaPU,V]� A�	5[��Y���������&d�#�!��U�ؿ�3�p�/m['=y}�g���.��Í�VjsG����'����ݤ��q�Xϟ��'c>�*Q(nf�J 
����iu�D�6�<�&*�Zm�+�'Z��^׶K�����j��7����YϺM�~��� �ӛ|͍�
��O�y܍"x~S7F��פb�6K��\���(��w�<5�����A�u���D��I���wCx2�Xz)��$d�⴬=ߪ�Uɚ��9moDv}�ș��2���؝��kf����EX� #�`�6b:��Ӥ���RI*1���n5n_��`�Y������a����j�
��.���22�uG��1�,y���;�gU�H�V�/SH˺D�[�h%eG)|�q���d� �b��MK,ܶ��񾮞��V�yk�<-�^��w��c��xb<8�B��,'�c�"��ͱ-�͓J��v��eɸ����;BT�nś��,�r8�f�[�^Q%�٬D�� ��]��󬗁ԉ�3B0��Ԫr/�
�O��=���W�=o�N�E9L3xH�!5~�9\$�5`m�^+O�W
��;E�1�p�\��	Ō^]ݨ��y�'nv���cVtnt����J^��k�hs"�ZeH����J���+�>��W��w]�ʥD�B����Bx�^F��U��q�qӝ���d��J�Z�$�L�`��@���H>��9������^dS면�\���lG	`�Xb8�6@X��i�f�/r��Pe������[��K������O�q��lCo�e��څ�/���w���\<���/2�udhۯTm�63q��P�:Q 6�&�o���BX��DL�}e������:���F!H&<�95������~)�R���� �1o�GkɅ��xȦ�$�0u'p�X�D��ӭ�QɛH�h�wz������F�х`�.B�o(���"��oe�4��8.�?v_���I��O�X��r��.�a-���� ����6�W������˛�I��� /��r��߮��}]X�i5�|�qqݥ���f��W��VgC�T��st��Ӱ9pǌ����*�tLS,�q[��²�i�������C	nM7��\f���WL���+�n[�"�Sk���N��arF���4�l�@��� �	�2�&�x�������O��V6M)��/���p��������&T�ĥ6�����-L���x�2Ә\�qɸ��M�g�v_郾��ܚw���'��>ݴ�Ru�[�x���'<d�;����&;�WQ��cT�4�L�J2�g�����&*!+�P�k��"9E|GE�x�&1���̵�������uc����zy�FA/�I����X@�غ�k���4,���~'�+�g��(^�I2��.�|�R������tչ6�0u�W
݆��6��fX|�H��x���@�]to���XH_>��d��"�q/��tY@�&?wb�:��}"a����P�&�=��a8�j����F8�	��b�ǜ� �+��`*��C��u�-���:W{�XO1�a�ɦ��	�lFF�&�2-a���u�h����8�W�q�J{D��Y��U�bρ�nj���)S�t�P|��.q�t�%�e��!� ��CB�����n\g��������#=�4?Ou+J�;yc��Ҝ��u����*�Ü�N��Ҡ1k_�!3%A��4���'���l��K��mxc7�Tg$�c�Z+|ݔ�W���~v��%[�����HX�ԧ�mDV��8rNm��p��a_/3Y��I����e1[�j��I�!D+�d��C����s3Â�u���j#Y�,�N	�.쫳Mmxf��Ś�4��� ��A�H30]�g*�;���4�;�vj`L��7�j|9H�=�!���ا�zO��K��uXa�� �n6x7��h8t֚^~Y\��w>��<�~Y6��}�|	_��4C�fg}�}:��3�m8�MX�r4.��<�]����s�l}֔f���/8����?�1��
�zR���먼O�����"�(+���7���ޞ�cTo"�������F���`zǻ��mM�v���l�kp�`p�^5��	�b���5�MB�@�?�!����=m�c��V酘����\��$k���`���DP-�f7ތ+����s�TF�>�|���"�2������T
r5,���,���º6��漜Jy�M���睖�/DhS��L��B\1��g���AZ{�<�Z�|l�^f��q����ܧ���U{G�ƽZ���	k�_��iO3��Y�rl�k�k��`�ͧ["�o
�*h�,�!V�Z�>���k��>�pvW;�EzZ�΁���n��[��i�ي�̑#X�ݡWr�K� BN��*B�Qv�D�;�CA~���(�@o_�{T���n���=��J��h��59 ����J'����;(��j�LV@M����3I��;AP{����p�O(」�d]����<������{���!�H�ɛ��M�Y��`���Lo�r�/rֆ��rp)�Ob�I#Aa�3�wl0k�A²
�rs���M�� PM���s�/ �D���$y�Ր��0�҇�1�q_��&�$�3�"*���H,���p��^x!��̠�u���'��v�Pzm�_���7^�6vpȚæJ���d'����27w��`����ޠ�_�/��!�l�d��q,la�>��h�$ �`�*U�$��Ŝ���/)w�TXfY�D�WB��W�=�zDƎ�	�!؂"��%�~�s)�=�MdΫ�0�2z���1���7@:��X��ߙTO-`�<+����ar�Vk�*����4L�T����F큾#ȟs�6N.�xg�����E��{"c�b�mY�����q7x�C�)���5eϛ�`��` ���Ǔ�e���"���7u��X@�� &i���viz}�=�y�ɥ����,��`o��A�^W�qi;C�䘩��'��y-���7�::��9k�L4&Z��4�C�~4��u���%'���2��"+��:,�(�D'c����L�q"����^�'��ו��K���[H%�Z�Z��Ԧ	|�T�Z�'���b"pH�\g*
Ǣ۽ZP���BV8�Ž�CJt����K#���kq�~��H�S@Y�A� ��@�i��^o�ܫ�T�������Qu�Z�`З��R;P��H��$)W��$]t�������ܙܰY`��Q��g�F�erX��j|v�C���OoZ�5y�5{�Z�tڳ��+�!��ɺ���:5mJ���]�i�f�
KLm�rM˖��~�&��	b�"T_��^�'����	��2E{��<�S�Pޠ��m�퉢3Pd�c/,y�0lf�=�Gm��զF��Wu1������q�C�K
�ۘ�1*N��=Hu��������x�"&�3��9֫o�?�Yp��*�ռ]'F]���D3I!�?%�o?�^�ݭ�p3Z�`�B�J%�-Sɮ#H*8�뜬�ÓA��'Nsk�*��˭:C��j��^��4L��59��.i���֤�HYľ(�7�͡%Ԫ�'��b�����7)���'�K�	p��!�?9�1���b���b�"��S.�������F+:����d0�2��@�󓔣c������C�L�m�ٝ��yJ�b՚�Z���ku|0�1��|2�^�?2D�1D�M�-�sfF�|�O~���F���{�ϼY�j��#	#,��e�n�>!��b#C��˔W������OQ�6x�J� �<{����SDv/:D[4�+���Ѧr��S��$��]�[S$�8,d'|Hk#��$s��ԓ����A�o;����֊�X� �+o����0hC�P],�d��-9�������$ٱCX�	X<k۩t#:��Szp�]d��mP<4��y�#����I��BG�Os1i~�oױ��=�>�o_Mw a.�����N���by���K��5Dܽ�}s�60��	w����+fF#̢�G)
-2菄��	h;�g�ܹ6���� ����B�3E^E���66����$C����*��$�����I.�c������;�
��|��o��?�;�'
#b
�˙�Β��
��u��d�1GЅ�(����Y`�2\�	��D]��kq��;C���k"��Q>�������$��n|��]Tz��ٔ�r��Z��^i���D֌�q<6����[�#�g5(�]���O�Y�n�J�NI���O�S޴�S��К@Tz]�g�X��7="�{��<���Ů�?HS�G�A�U2�w�G�u���K�KE��^�w�#���("�"3���ؿ�H��P������g�0�<]�q�N�-Ӄ�� rl��/�K8%d�A�Ԑ�^n�=�� �����Ϙ���i��zAߊ�I��M�u�5JQX�R�-�̧�h����X����B��9���� pO�`����B�.	���k�$�l,�O�̈�lW�����Փ�{&̾L�)�v$�b�i6j������j�r�����Ѳ���~H��@���a=�|�?�G���8T�m'���&�aV.�EjI��ˑM�}���*T��h�7���A��KR��A����!i�1G�l�����ȇ��W�N$;�L�Kk����� �k޵��ʅ���r��Y�j��S��A�����[��-�+�L�{��ZpD����H�J\�"���ǫ$XI���|K�@Gm�]o
�6�t]�L7�L��?�Z��x�P�j�)�3z�RkT궁�O�8yҘJ�c��Tx�����ߏע�k�%Mn�Q%xH��xE��u��܌�_m�5��M#��oyM%�5�hLV�N$���`�)f���M��A���:�ua��3�z	j��jn����ʨ�H�0��w�2��q}���2��2u�2��I]���mh��q���ݖ� j}���N��JSl�U����L`�$3-�U�
g�SEc�Ѱ����lןf�.�Q/H}7"������biS�-o���ť$E��,~xy��m�����on^����g��/0Z��Ev?��ʱ؊/��ˇ����)�2ԕT��[�/����'�����}SX���-�W�;e���A�C���T��ð�BO�TKK�)�q�i�Q��Xb0�`j�#�K�x�;�:Ği�BraU;�AmF���*ce|��au�Cv�;�u`pWJ<��q�i���gR�w� �[�9q����e$��Ĳ���,w�N�es��;L7v���1$liz�Dfʿ�%��2:ܖ��\@.p�&��(WIԜ@�AD��xz~#��18D��e2т�&��Q����_|�sb!�~�}w%�l�!����pR6Ւ=(}4T�lt,���
����{1"��߀{��91n�TL�ZQnn�%���VX�`ܴs���z \������g�zOTI�۰�h�{�Q tk����^���Y/_��`y}�=��:x�m��Z�<1mZg(����t|rBw�dtM.�|�B ��旡9�#�Y���X��װU��cy��F�@i���9���S�u�ԩv�<�|�	�%T�zե���3P'�ئ��j+���z-ʑ%�o�{�]a���,aᯗМ/�-޸�(�%�����|oCDS�jn��m日��n��cK�4������ֆɬ��xZ��&�����EDG\�Ȭ�%F7�Mf�Xib�����e9 X�+�����)R2��$|5�&���c<!Mtp�P)>�H*���C�᨜��J��I��uq�{�%�ڷ��X�����w���X�q��m'���.*����nb�m�ΞE�']����t$]8�g?������TCk	���4J��,aW�a�^\�BRg�M~\��-���oz�����Q�1�z�i3�+lS�jSA��W�����mSj��S�����<Z���e,S�c�D�U!��$��vRd׳8K�]e�ݿyz��q��if�OB֙�dK�y����n0YIo|��b����Ƶz���Y6��s��6N���5��h �9[��b�j��	��$H���d[������6�*!�1h���m���
����M�-����7Q��ú,$�̽4D�''��3=����h�[	�p�ǿrm�uu�����E�m�4�5�0r0X��v�b�����k���w%	���d�6w��Y5�K۞F����$�]/��ܩ�,�,�lx#O�9&1�@�y�=�Ľm��z�m�i�����)C@R�,u���[��mMAhV��+�t��G"��&Kc��J6ֽʩ����(<jF��ʖN��ߟR4���7M~�������Ri��Myi�(]Gq�Jц%e�Z����,�N�{�%��ɮ]X�.��	��J�P�U����e��6�f��\��dF4jkY8H��;����zl�m��NT� 7���w!�b���;��P!�h�,!G�SmA�)hcm8?�"�uK~W� �~�Nߖ_X��I�}&_��@.�n��m�
�#���S�:HX��PD�i���w�<@�?�F���q$u���;���1+$-֖��_S`��N�w��Ѳ�f�Q��F���q�|_�o��l�lS�i���!�e�:2�K��1dN�e�*����o���{D���zUpn21[����8��>{��n����Hz��˨�Z���N'��('��L�B����Q-�<�?gS-���[a�6|��|�N�Ҝ�G�g�g	����&�Q���i����.�B���)����y�:�$t7�^��g��ʰ��	������)p�ϒ
Q�'�P&�^���JҪt_�@�|�@.����G�Pv��VI�g tT<��@�+�{&�l�?��j�$"�X!sɒ3��o�Y�i�FAx? �P�ً�V�s��0E�WI b�?���y����P��{Z��v�2Y��^95����v��+�:�%}'#2��)2&��tR߾��M�.���k���լÛ0#8��ך!.I�8�r������u �F��_j4M3���mWٜ#�d����QK��Ғ�lM���x���G���٤�{�)�c�e)�E'ຍ��Y������@�1a�Q�Y��o���H�aڔB���^?&n[�N\o��s*7��	��L�ՈK@*J��j���%�����i�$=����u���@V�4���:����C@児>.���Iq���Y�9&�s/[�b,/󤛢ŶC�D,{��C�S_��� �M�TI���T����d1��zp��q%��lZ�?���CE�eT�x)�K����y퀓��)��c�s��،5z�����0�C�I��2m��\۾��*�JN�'p���Ⱦ����R�C�y��Fmc:� ��{ml��!�^�*?�����i�@�W��6 F���dd."��"'�
�>	u���~�K	2ԈšO��7�u�� ��f	�c���O���m흰����k�o_��$A���G�(����JB S�5�C�_�ƑaZn��Y)ӪF���L�a@nOt��6���D
�G�3FS-LN�I��U��C��ASH����$ڜJ��Τ���Ǫ�E�U�
?N� ��������G{���Uf�C7�|8�鍴��7�O��a�����v��h��yhd[D0S���_~a�	I�2.~�+��&N��H ��	�զ��sqJ�������a���`�^�;i�z7�{%�yja��WG�"-�V�I(åd��4˞����i,�N�?�/bG�e�]txa� �lsjA��T�������nh:�ڹ��2HBL6k�b��$ ��T~��j��M)S2{+̈́E��9��us#:XZ	�%\L�������I�*FYT5��&g�#��BD:�9(t�&W{
��4��y2d�y3h��S@ԣ�� ��]� M�@�;~H�>��h!��݄t_��&�7T�,���8W�h�͆�*���C�ӂ[�!	��T.�ǚ�9j�G����� ��؏.J�,�/��̾>MCŶއ@��`�Q
�	��ᮽ	�9��Έ�@3�d����l �6
*�=�I׳|i���@ھ"�eQ���'���/��!��?S�ų�/q�YE�x�>�����<�n��	�o*ඁ{�6��f�Hɩ���,����}���ݥ^N�W�m�ϙ�KbQwSM�p��F�� u�'���������h'��<��c�`���-0�Xr���j�ôǽ������Ҩ��M0�̛NcZ��E���}�A���D�]yM�y#��eJ�~���_p���p%���ޏs谄x:�\dǒ�����.�g6L� z�iQ:
 r��3�?q�ì�MH�I ��5��Uf�`�YB5��=e�5V�ʂ��i����D��8��Rvpf�2����c�K������> t�םcB�~�)�Y���8��؁��-�[fv����cIp���5j��!mz����@�����.A�P��&����wK`b\a��l\�U�I���ไ�nm��K3��������U�AIV�&q6�T���W#'�),fQ��4?�gQ3[w���m@N�Wk2ɫp^�h'�1v7THO��g�|P<�'�yV&w	�V���p��l�ϯK4!*��V�+���<��Ȗ'��%B�_�+���&1D�
lv M���q�s�@2V<NbL4�M.R&�k��@�	�y���>��c�Ks�^9[������ap�=�<�~�;�j�y��C�D����3.5�γ��h���Xh]\ G�G��=�,��"F�7E�%7�Y���� ��H
�+�v^���Q�;ܔ@���ǧϚ��/{_w��ʅ_�0�!Gj�yt�0��4Uk#�"���XE���%u>=�*|��s�Ц�dUr�w�n��F[����&��4������%p�e,�q��_���n>Sʦ�=���H9Ӹ���2n槔x|�`;�R[���l��*�}��9`-<�w��/J:�eטqCS9d^��J�c;	���弰�m�|�"�ЁHq�rD���U�h53�ocG��ω�ýĜ[�p飔�B%S�\��x�,`W�G�S�EhN� !�<-FY&U�l7��c��0�Cӈ�4ą��n����be��7ޡ�1��\��3�d�^օs��R9���CC�o�N��=�0��?W��,0�!��A�o����44/��$j�mM���bE��r;�>��R:������`�(�t�C�w�Y�5��$ ��G�����̖�~����������_rxU��ۿ�/��?�a+N�NS �n6P|�b�?�Xr��(
ۖ��u]y��0���\o�.���;]y�湮�u��aL���$-���T��t���<
�U�x��|�5E0�L	^�X;��f�%�\7��M-g�Cy�SO�{�0����=ͩg_X�ѝ�]��_$r����h7���5�+�7�L�Η��G����4� �ťw[1^̽Ä�b㪴����3Z���.J�B�r.�U�w6�ƭ-�^4��=�͙5.��ۃ�H=���A����kۃ04Z��{���y~�( I�]���r;!�l��ߘ�_���#)ҳ$�~�Z-V��jWC:�f}W%�yB�,k�eT�\N���D�� ���Ǡ��+��c$7�Op��Ҏ"�NlN�A���*xnȁ�* 6c�s�{��+��6���sPb]�ԥ�����!�ӧ���D�X�.�%��YpUژdz�ZD�����G�u��w�7��9���MK&�t���c�Pv�C#������O��a�~!u��|0���0/Ax�K<�;v����蠯1>4�.N�([O��i`��u;so��HX|�ތ�q���!퇪�Ȣ��� gmƔ\-��İ�m��p)>A#�