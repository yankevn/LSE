��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf �d���]��c�Ɗc�U=_J�	��w�5ޝ�:4(��ݥ4FM���8�(��	t�6�/^�J��G;�#h�����,�JB�V�g{�|��q���17Ⱦ� �-w2�1bfۇ�z��*�+16�/�\��<7����-���*��Y�����8��+�.�(��LE�#߳�2T������.���Q��W=Hp����JϿ�%���j���ԫ�����k�Q����%�F�����򿗘�4Q����p�7u�4n�F��W&vA�‛n�\�N^M%��OEԬ!I�졭�����D�=,�H8�K�	�U	T�9q5����qJH8Zҙ���m�dXm�'b�9!��润U>��h2�$�y�t#���5���-��[I��,o�}�ڪ��3��2���#--�憏9S��;Z��U4*d����T/q5��䱩'�Fb�i ��U�X���f�c��Ɠ�����y+,�b>a5¾L�7r�4nd�0e�w`�9Α�# �z���sX]h��N#��V��¡�۔��q��p6͞�RS�c
2GM?�o���x�F�2�K���ԟ�0�����p��X��A]�*-�Ǣ���Yj���*�WWD�ܞ-&���ZՈ�����Y�S{2G$"��V�	�q��y-��58=���X�� �J�r�C�^��U']F���y�r^h0+g�&3J�5��|]ˋ������!�G*�i��C�W}b��Z`�3U�����|WzN��&��$��fo`�,��2�iS��6:������Ps�6M]�KNJƺ�V��zm�����������N���v#��%Qn��n�G��n_{�:;��勋AqQDl�%�t�i6���!��P4C$�y)vc�9&-�\`��4�,"�W���	LM�.��?�@�琲�}�+�V�����.�
�S�O���-zHU^0����`"���#�iv�
t�<�!9v�������s�z�f�BToC7F�����98�L%�Ya_}D=K�j_�B�z��j���Q*<���V�'3���i���1��bM� ��O9:G_�j�l���^˞]��q6���wyg�,�xP�����`�<�%�/�wd��d�g\�H_���v�)�7fbXmy�Yl<����N�_�¦�����N3�bs�.�v1��˯$���$}�
0�pE, � ���%�
����u��T�?(�yS}!�n�=?Ť�U��#3���SC�c�_~���2G)(xG�M��'�������y8��r	6,i��	�$�&} W�`���V��9�n;�H�XS/��u���pY_p���B�)[`8�����Z���q3�R%pc?
q��*�Fi��Zc݉��y����ٔ/��÷��NW�*�OWQ�*�"�Y_z�Yx�6��M��	^m��-@�$���[����w�u��udkjt`�^q����b�h�a��$��|��UxEsxJ<X��~u�!���xӉ4޾�ʅ+��xDĉ+�`��5ZR�Aj��I��x�_ٕ��P���@�XK�Y��L>��M�`�d�,r(>^�ܤ}��g�7d6��N��À�O�_�P+�IʚZh�����y	J����S­_EӚ'tX��fV�羀��ө��uѐ�+x4���W`h�S�FI�}@Bq	z_�_�Q�#Q��C���K2���2����_"����y�}�_LC�ܡz�0_#�5����1����k���/��������}�F��Ř�v�\V�_*�K�j9��XK��?�%���D��\Q���b���%~�򼵹���ZΣ�L�Q�*�����ћ�V�Ţ�/BIW�4��R�\ND�yN������mp����O�{*�M�q�{��ؾ�ր�V&L��F���I$�[å�;�;��b�G�/��"�Y�Ѹ]�]x7k���(� ^f� \�F�q?{t��l�5��nB*<�qc�!o��r��