��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~�>:N��c|�M���WE=ҵ!���6+�%ˬU��ֱו�}]��*��f�]x�Zm�'.+=�I(aY@�#@˜�f�E��F��w��Ұ
��-ui�*���a�s��C�33��6i
 ���N�ό܄q��@U@��ȸ�Ӂ�ŢB�6��Q��Uq4�tx7�T��6�k� ��읻�����T}�i]v�G�����@*D~E���Yq����G���RG���LpV@�M�Oh�R��w�\�N;��(n�w�7�Ɓ�GfG��^�M�#Y����R���j,��B�>�q�~�D|:�ٛ�EU�h�HU�����w���p���-�L.{�׺#R�f�Up7q<�����֮ҋ�9�	~���Q����F�@0Y�y$�c��b-(䚘ygG=u� +C�N�"��./�����P���v��g��/Lb�50�T�(�(�x�-u�]5�4�X�[��f}�� ?:��=�6�JuN!sAe!�`tr�Y̗�HTF��E����<R��ft�EP2�Ǆ+@5;�v��l]��0�&9��D�>M�x�ȩ�F̍l�x��:֤x�~s�&�	�0R�П���(C�V�t{|�-D��X4]N\�t���*k�4-�3i�n<G#X�
V]:���P���7���I��o�3k���1�L]�� �@wl9��=_��yJ�����^�j��S�����l��[�z�h��Gk�L�N����0�kc���2��u&�=��������Y�*ٰ)��G��억,:NT_���.g"����.ⅷ���"FA�������Z�6"�X���0��z�H}6������O������ڕ�����Y�2�pf�xu8^��	̷�1V=�2E"-�ԧɶ���|Xy�$7�X���{'��RaM���}\�(��y7j�Vۀ���6l�q�&J!D2=%�,�5��v����K[J�Mr�4���B��n����P+�˧��X�X`@]7���ݎ�|��^]҇
er���m�Rm���Z������|J͝����k��	:㙰��,V]�v�_�TU00�3ڄ��(q[o�/���fz�����\�#΂ ���g�I�����y���M���S�������
[]nf`Şh����!�i���?���x"���Y|A�E�^��V|���!�
�i(+��PX7�|-�Y 9J�,�j��Y�c~�!��mZ�лO�rn�!�G����1@��\|�T)�b�?Z~%����v�3�D+K& ����}�&��3Dw��5�Rm���0e��Y�O�Ϻ�B��Е�1���IH!<~�\�n�.��gZ��#h��'겗;��rl[��Bq���t|�i{g�
.қ�a`2�����A.*q�J($uE�����^�-�i�W���c�H�k�!�I��1GX0,���e�em���\����Ua	��Ծ�vp�:��6K�:%�`��d_���Ҙ�����\c!�u���ti�l�+f���QN\2n9��Gqb���̄�NG�F�
��˻`j��!�Q_�js���V
�߮qQ�\ӑ,y��_� <�W�˿~�����3�\(���������L��%;�`�T�p�T$��~�ۖ���s��y��x?J*x�$��`G��K�N_����8d��/u�F2{�L����\n,8Y��BV�Ԃ�1��U���g�f�}kFm���o�$Y��!�J<�x[�`c����K�[�-H3ɑw��5pa���|g�W�,Cv���Ma�����;�E�}����@U����3��J(p�3�C�%���W�k���'�/3�4��2��myy�V��m�w)�^^m��-����қ��0!7٧N��v�=�3Nb����亳t���JPE�����t&�A�E��t�nɭO�i���\P'�������\BC!=
{pDA��z�'�y^��2`5�9�1���W-JӐ=S�္~���ѩ�W���\�'}�'�Ƭ�/� \�d�xN���^zf�
]�W���y�� P�m4tB^謇�pp�*T�֮�%�x6�t���
����*��@�=ӈ]
����\u�2?�ȿh��ط��ⶆ+b�G5a�T��j��-�e���P�oC!�4��'Y��zbF/f���<��6�c��K6]\g}sҁ/�`� ���$&��4�K%=�q�O�{P��5:�J`����[zQ�shFͥ��I��?��C��K��m��Q�fB]_��x�������ѫrP+�t����J��x��)�BTy�x���	������j:S���Ǿp݉��-���b�X���Buj7�v}�k����I5]�lҭ�����ַR�Yx�fT@0�L!ϔ�5[v��;3w5:񷌵�[7%��
s��e	��儒�Op"߇z�&��1�(�&�w0n��!�.#۠�z��Ǧ2+Y�r��UuW�����VF�k[h�P�
�5�*�$�ӷ��^�����1U�X�wEٟj�v�Nծ{EF��t`�2%���ϐ4>�fbd_��f�(�gѲ�P�Z�0W
H;Ԧn��q�1v��P=�Ri�P �*��Yw^���mE]�������[��&VI2c�D$I���Z���dJ�ت�Yb��B�V`NB���ƈ]�	�q�}ߢ��3�tI�C}5[,,�[	�`N���H�2�\�[�A��:GZr����}�`������In0��d�lc�E������T�-��g�].���>"N��e��Rt(h�S��eV�mʖG 7t7�bN��
�'�/a�S�Կ����7�H�����9����͈��1�^��-�k_��R܊������HH��B,�[,/�Q�wkU��5�B-$Qe��r�%�����W�I�7b۞���Y�7�x�؞|��Ǚ?
�E�����=�K�X~g���� �"cTwLѡa��w�g��B7,�P����j���`�j���g���hyS`ٹ
޾��Y�g m��j����?�ۺg�E��3!������N�)�)�,�Q�z�f�b�7�~���"����j�I)�ɯ�5Z��~X��ТϏ�#�FL~�8�U1��>�j�w��ܙz:b�/�Ӽt|jz���vP.M�u�9�!	��C�HUBxsb�Z��_/tf�|������ם<�$|�C�?��N���=+�k�`��;דS�%��-�x�ͻ�C�0��1۪�ι�~��,h��7鳤��s3��o4�U���ʀ�� �w�N~��bھ43������A����}��J�mӓ�Q2^�ȅ�w�J�a0�L!E�u�Q�+�:{T��ao�rúQ8�>>�ħ}��s럧���E����.u#&��X�S'A6O�*\���:R��/�-�w>�Z�(�u892EX�Ȅ�Ǒ&��Ϋ0���<�{wJ�*'��5��x�����O���Hn0�N(�������
��l+,��3q���@�0�}'ɾ,V��bD�nMՠ���j��F��=&�vK�7�N3X���.�c��%����_�gק-��j�R�c6������7k6�+���7G�<�ݏ��M!�Ds�����Wad�e2ԉ�U�:�l�;�%q]�!��9��%y�/{WDY���fSU #����8�Lj6����V�(�4@��lf�j�*�k&�Q�=sxCBƊ�1ObDJkv���G٠'H�i=�dj��վf*�o�$|�{:�#��=؎��?���(�H�Sp�O��
# ���⸌;���b�W�m�W�_V�H� ��_O��==\�����rG�6F���Rc��u��\�;rS_ܭ�SN�vp����Ze�"_�Ѧ,�m���:=��!y=<�@�X�!�E��������c�^9�@X���@��ٵ�5�#�ai��="^�fz8�"�8�.��-�}	�� �4"m� ᑏ���m�Ğ�q�cDH}#T� o�ٞ��x�@w���{��� C�b����m�r���Z��Ŝ7k��<�m�o��k۬�Ϟ0&Ho���U#M�>�g����+ƥW����3S��E�����b��$@�C�ei�(qpѴFhL�Ո�A��n�2uX�  Թ��Ht�mKe��?�ޒn6;�M>:����������贎�;b�lգm����r�	�}�Wϓ�֢���<���A��ѭ0)4��}:����@�0A	Zݢ�҇����]=����7�<���'���$M!e�p��RրQ��Z�����}{���} ��B% @�8�����{���X*�e��4�k��R�|����Q��|Ҹ��M�M��*��jͯ}c�P�BL=~�s�(�ـ����d5�QM}�Z߹H}BbN���Y!,U�/�JLu�ٳX�aH��I�������g�ޅ�C��G��T�+�j��0�����)��br�J��L��%#�-��E�~-�,��	)>eݕk�����8�J��*(�ִ�ôz�� �R3�%f�c���+��۾
����Z��V���B�����}�j�N)����]p�)�����}l),��0k#�8��ʴc��ꥂ$��A|��$��Sܖ� ֤)ޝuG��W?�#sJ��Aսp�N�R`8cx|IW0���`h��T�QΥZ6|��d41#�q�y���"r*�$ }�L�a�2~��k!
4�8r���K��1z1�s�P3`�R��$��v'�;-�B����BV5�H�K�~0ə�v����|!���pw�����LʖC�o�Hi|:�������n��W��\��>��qrF�ǾPy=o�3$v����Cf;�aW���2���ZxH�Qץ��K��S<��q��[@��̂���c����Tfkf��T6�t�h��j���{`:2��-Ɇ
��	=�:����
絰���&���B̌�j�#���=q�J�	�T̮�P�s���}l�m�s��U��\��~ȊC��.=��d�v2�W���;g�2M@�W���{�+Gfrc��F�1�D�����[J���˅����Fe0����+;t��qg�NM���jG���g��?����r��j�ȜN��)A��Z_PF�eA:�jS�&/+S�Saa
�T̓�"w!�QP���~�����R�+j���q4�g�C�F����rPc�~ 1���E����d��]>�l2�[�4S�ms[��t�w�� n �FT�I�\8q� .6������MQ4�H�Y\G�g��xy y��c���0�'J]	�Ɩ�^�B>���V��T��xb�;�j�ecc>�@���!��\H���!>6'&��7�Su�y�b,�X���n��RR���-��v� �,IR�n֌%A�I0~���Ex���❉��b�M�{n�Y�
��{w��]G�펼�n-��x�Qm&�7j�s����bgQ�[7�},T��\�WA��#ڂ��
�uK��)"5⇎b�(�?2��!�~R�K�1lx����V4|)bUo���&bֆ�Z�*��6R�0;Me<���t�
~�U�<6~큒�B�a� i���=t��� �N���|�A:ܭ8�T�����t������6��7o�P�Sb��bs Z�����V�B"�>;�<�[LF�Ĥ%W�g�f���p�ex�9���Q��?eU T;]�<F;`�í�j�V�~ld�H�ζ�)�V����'�r�|@���*�J�����v�y>b��(}I��]N�P:q��z��6� �7��j�pYaٙһ�,q�R���{iq�G�Ƽ%�s9�L�o�We<����/��\G�RR�xM9�T�����O6�����f�z������˷\�;(�Խ�V��l�LTʊ�Yp�"�cE�4ȿ˄J�%��Nx�4�O���IF�@���gլ�eV�"��_;0D�r:�
��z��:t���|�^~�cgy���>�Ʉԯ�ѾQ�qD5ſ.d\j����+�G�VG�ґ�!*#�P=6_��(8����ٮEt9Fc�w�׈�tHJǉKh�ŏ�+�¬&6Q~Z��LSThY�U�]
�'{��#$��}w�Lz�-�[ǯ����7(��s��OF�J�/Z/��tT��
C���#��w.p%����t,�*�%����D'�J�����vT9rY�� �э�O#߻:��ד`�|B�(��2M5�E%;g�A�s��w�']�Ǧ����)o��9��+���vLT����f�M�n���_3��Je7�2*`p�-y���x�@��<��O7�;��!�q�bݏQn\��>�Ƕ?s���\���/4�z�R�M��R�*�����k��1�"��<�a=����;{�w2jY(��Z���琻6�q�����#�
d1�x���.#���V������C-�O�ӓh�+IW�_���S���.Jd��}�
�Z��M�y|�z���e���7R5 #�Eɓ!��5;���0�/_i������ѽ&��(Ђ:�A�"������"�� :�Kx��W-����%�FP_�-����j��b����&����R�����lPAS˙v�&*�i�*4�;��֓����I�s�zц�
�#��g5(�/�6K΄"$ٝ��hOi���h��t4��+��zU�y�N�����uV����������1@�V�$Hc)K�ҧ-��^�@���3�R�K�%|��w���N\][˕ۊ�D�����m�"��5���QJ��K�V��.�r�h�#��?6{���L �[.J ���gs��lGM�̺G�Q�L�=�Ԇ|X�i�u;�k0�o���t�l��~�v�
��s�a�L�|�,h�g�t������O��w�P:3pOB��Q��rܔVؒP���GF�LSe�s9�`OǏ�'J���'�߈�������4��ͫ��2����Ñ�!���p*�V4��j�"Y�䦉LZ]_��u��T{��
��h�?v�b����(�P\\r����H9�ꐊ�R�-��D�qw��)��_!�r�-��(ʆ��e���G(N�<_���bu''�c����#�r� `�`�+mͪ������ +i�&Z��P�X�ᰦ�uG=�P��X�8J��N�8��kV��-yB�z��7�W8:2X%�T3̫VH���T�\b	^J�%W�?)�Y�=�i���=�W�ߴ�8����qL�Fň����1��`Z)��攢.o���ڣ�zb�T�4�t*�H��o���%`3=L�u�����Jɍ��έ*��p&�k��m�� _z���uE��f�C�