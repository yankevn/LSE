��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S���!���Ӕ�4���ǥ��,�%��F����a��Փu�!Ρ�'�h�|g@�G��v�����#��t��$2n�"��~"ٙ�oT�C��Q�x
"�4^���z��bˠ�3���>�/eG�<X�{w��pKG�kX���fí��Հ�trl� |̍�˼�'��>���Yƒ*���y����::+�_T*�:��UN�C��
��vD�_�Y>Ksb.�k0�k5�|�~�3�N������vtU���r�(ӛC]���Ѽ���'P���F���|�MU�y��y���q��=�J�1�y*�c�4)d�X+���L�����L!�H�G��\��e�OS$��S��\FL�ҁ�Ae�k[әs����b_��a��@���W��s�?Q�G�T����;��0��ʀM~�(`n�eu������N��eUk��Kg���<������	�,*�p����	������I�s�;�2|�B��O^M�<�(B��[X~S�pjfD�+����*�F��N��l��^l8��x��|/����bŉ�@q��q�k�PU��xpa�������c���F����P�훊k���6\�<�L���x�aLUs<y�딅�����@��6�6���82[Bc0E�D�3��5��I�������K��棢���P�H���K}%��<�7J�Q*��?����)L��FQ���Y���&D�u�%'oQ�C����|�q�R�J<���odLO4��xmN-[���*���t@s�<��x�n����>�j��\�r��@�yW׋�(&�S3��l�,�g*/q��C��wUfOi�=*�B���K��H��?h/�n��DYxǺ�.�M�i�1�͢hFe�g\*M�p(��bL3�uz�jp���0��K8n�F?�1|-�4�b�B�EY-�����21����᠗S�Pv�;�h)bc�'C�9�O+g��w�*�����X�a��x_���>�`׏}?�[hy�y� d�5�u�~Gց��;���:�*z-�:�n`��}2��wt�@�u��F/���x��J.R���f��N��i^5�n��e��L��&�}\)����m"��n���u���q@����E%3�@��fhi�EVg�<���hR �9}�����U�Q�w9�b0��I!(�\���w9�VqC�V:�mi]��h��.NéN��Z[���X�=����;�[�4�˃:�~xtp���n~f��Z�u�錮��8�H�O��Ճ�T��t�Z�˥P��L��P�B�)���K>����Ab��C 
��fЬ�	ucO�˳��k?����&�Z�E<*�Y�U%�^:��g3���a�{g���p���ؾ�>��iM����V��(ZBNi_�B�
5@Z��O.�?6��4��ܗ��]8�%&�r'��t�9���SDב�S�5Ig��H���;@�K3�mY�w�6f/ȑa��%�*=L����e��E�lB<H[����@}�[����."Ba,���VE�p%�.^���U