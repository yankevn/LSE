��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~��j�w�s7�����h�8�w�D�&Yma�I>����L��n��S���j	��	��i���W!��l�	m�m�zQ%�yݓ�c�r$�hZ�X�C^���x�s�	��ua���%~��t�ơ�����R����~H$�pRv��*S�
rD-��aS�N����̙�ARvnE�J�f�f���#�T7!����:�I��*\,*5��D��~@�MakCN�z>	�t�0����*��>8��l��-v���ԉ�Y޼�G�N8N&o���Ɗ���xe���;|�l&(���&<@<��T� g����Q0s����C^l�:��C�Bש>�
��;�$�)�s��L/�@���rM�mI��O�7yi��JV^0⇥F䰒b�|_�򭢔1LfވŞ�ք�ғ���1�ph��`��o���{�ں3q�O���@5���Y��q��T�M�9'�����0���%5�C�>�HgT���F?�6v�AYa�p1C��x���xfL�t�o�/B=�>�"j�rH`�ٸ��b��k��4�었��tø�.~���}y�`�:�jϚ��,���W��tŦm�ā�AP�*9��d����%CR�A\<}/��}+�Pӫ1��$���1�)�HPˍ��1(�@
7��U3>w�@��A"pvl��;��:���;V *�`�y_�2����h߶S�z"���0����'�y�S���7�2z Rޜc�UL= �4*�17r �s_�4P��&�*X�}>�\8�7�琽_�wx�F��	]�k��a������!X�#���`�Y�/�O�h�4�Z�9|
��FE��S0qxC$P'���{�o���z�15Y��l�KIݠ�����Pm�Q�0j�|�JWؗd<���Xv�F��."�|�_O��6�����Ba�U�jLC�^+���a=�A�����ƴ������w<'��N�Xq��֏I��D(�'�Yd��si�9\�sE�����"Y6�/�XLz~v�1�7���������:\�\�S��s�"#;8��)!*�e�X)�-
�+WRs	.�hZ%%��>��'R�, �6�m	��9�"����vO2��=�ܭT�Gc [�����$�t9���A����%�6�$�L6Tv�@/?�*�^`��El�I�q�j�v|��G��>L�#;F�ċ.86l/�
��,OD�1\�i.��Q�i�x�</���]�믌��3��{�l�PU��U8�D��)�A�3������ˑ��8��,��B�#� ����Þ>�J��2��.�؎}œd������EM�Y�$%����i_m�*;�gV8$�L��=�&�aQ/��3��:���5��=6��w2z4�N{��i�����gܲ��O��K:Ű	���"�h��U��}���$�FYϷ�{\73�R�~�zS�N�`��:h6�V� ��s�/}��x�� �V���x֝R�oi�X��~�^B���FďS�L�t��žR��V8RF��a�͟��}83D{��HGO2L���d.�.�K�l�I
9L�d��F���w�x �5b:G��������UA�Ωǩ�Uw�&"�:0ܲ<o��dBE��+�$u��<�z����\�)<B��\�0��e�������Q�S��(b��	l*�mT!��CQ�$&)H�{�^�Ѷ>Ca�b_�9�+�3+�A L)����L�g�5%�7��tM qE�DR)��s��d.8�"ũi�ݺ��8�U��u\?��u�7�^,@�����y�Kѹ�)ֈY�nKd�����c�5��ɲg���h���&b�`�Ĝ�6�Z�!�Ŧ��F�(�%�$��f�{��N[4Mm����<
Iݼ���DD�x�Ŗ�TFG��� >�����G��*��d4����1��7t'�-�����R��>v''^w䁞b����ޟ��<��y �I�K�	߸��)v�0�NV͔d*]�����p��Kl�����ޚ�֙�Ĉ�hz���?���5(�Q�^�x��ƒ#�)(}�^UCr�L5ڬS�߈��5�.k���/J�0z�&`�T^u~|���T<e/��,�@v��zK�SF*,�"������Y�¸��0WڐŒDQ(	��y<�U����cE�a���}G����o]���n�J{�-�R��iq(}��)ܚω�] r1�^�l�
�bE�f���Z�������$E�q��R��,�
�66��� @)�������n�e���'b����S<������������L.�`	5�g�XӠ§%�����Nv �@n��KW�����\��]v�gfSܣ�^�Uw�}��jf���q�0O�2���,�� ��52l��i�D��٢��u�ZVM�����0�aV�`)�\��,K_W��+���VclW��*�I�kg��8L�)A�?��Բ����6�)\�:	�<]h)�wz��'���>����mL�S��b�wC�s�G>`�HNV��ϩT���r��uy��6�^R/�|l<����ȳI,hݮ����>kE�m�ީR�\�,\g��>n�3~���ҿ��C:X��!�vf�D�8�
�jV���Ó/z�� u�t7�J� �y����	�a���������P%i8�!��W��ۤ�D�?Oz��=��������#Ӗ�k��J�`�Aa��Z֥��śù�4@4��O� ����IFspǫ�]�;����yZq�/�KW<��fdS|�z��P�Aɏ輤����K�-��[��R�o7Q����$'Jშe�m���,�$��/"�W-�S�	�/6���FB���/��7I&��_�"���aϑkHPf�G<��XSgҝ� ���t�!�W��r�PM��Áڴ�zF����|�h8+���+��&��#))y��/#89�f�X���q']`'�nmƗҖ$e��p�H���!��i�g�R81lr�q��;�R�\'���3�~�,d�N���`Z��ɞ���O��ξz��K�x����U6A�*�3��e
B/&�%)�.D�n>�c�ｸIJ��p�5��q3��Ճ�Цd�ؖ��ğ�-����T~��1S��S>P�{IG�݅q6^y��$	�#��n)ɰ	�w��7dO���)瘔��X;��5:�eL�ht_l�L=pH�-3Ȝy�^�X��9,̹!��	��^ Its�h�(�j����v�x��U�v:q����op��_J@���
�n���}�<��AC�i|5	�������w��x��V?D搪�����;0?U�҄m"N;-Y|�`C!|�72�Ƒ�3a�,׆C�n�(vx|K��BsIdjf�Ǧ����y����-:0f&��W�*��wE�>�0��v��t����s��HŪ��`���ɚ�hk�L P�a���p�O�p��_�[�߿�)��R�h�����;#鰩�ڍIq���,���l^=�� ���H���G�@86O�W E��;N�
p9]dpi��v��:+���:u�D<N���-�y\�|{y��n����E���q��/a?�m{��7f�hk�mN����3ho��=L%�~|�Z_��PY^�����*m.���Q~	VzӊG7������]%�)0�ǗE�+Ʀ9��{�����59��1���l�ϐ�@�;H��ԫ�EY�Y`��W�#���*N>֐����Z�@W�Q���	(����>��P����i�X�_���p�`�R[�w� �~����Z�5&-�2��N�K����V�� 7A��0#�jN�Oa^����$ɯ�ޑ�m7d��Zce����n���/�t2á�0���M4�ĚU�[�.ի��@���ً�n>*��0I��|���i�=��x��wS,]��>�����]Ʉ' � ZG���J!م���2���@L���ǝ�����|@��e,�����T��ϕ@�-fx�}o��!H�-��d�ѰlQk[d�ᜣ�r`���4���M����f��)��&�z��e#-��'����z2O1�`�����g�"��^v{�kh�/�N��
�T	�/�~D�f2A�3@����c1����A�!;��KS c�`�\����/<y���}�/Yw��Ps�vBbTvp���^Gnto�C:���T�Q~ݱO���ޭ��� 	���F�DU���*���2X��AY.&=�<� B�)���B����2�Bd�o�Tt`*�B��dQ��R�����*P�&��J�Bj����#�T6�����:D�.����,d�!=X��`�MJ�O�(�a��%�U0n��#����:w����zO(�rC�u0����p��:�S���U�<a��x��V�(G�����<1OX�y%eC�D�%ԁ	�Y~�Pt 4����e%ZW���V���9�	��r��p_+�w��|��d�Ķ���'rfs+.�%��FEw.j5ڧ��7��/�6��Zٯ���q�؋����xO8���72K��ߢ�|�Ͱώ#�Y%���@J�~�.��1Z�zc�b�6�����Oěc�*]o�`ߴIϜa<D}�
6U�_U�u)�]�ޚ!��j�cY>}���u:���n��djdg��<�kH��'f\"�%���Q���8'k�D���v_���5
�*�^�af�Qۮ������R ��%�o8�=�竬���.&���_�\c�y��p� �E��A��/�-7�l]���r,ƸD�]ߐC�:��c��1��L6g��&l�)��?�y��4�ENɓ�(r��l~�|OI�Q��par���qp ��J�U�Sh+@;r!�yw�>�s��tr3k�h�V�m_��%�ӭ�7��_%R!��r�b�n�wUh 	l�h��(4����^�*�7�!>9G��J�4�c�6�z���1z-�$�7�2m�FC����飫��`l��|�f��9�d�A�TD@�
Z~��knm��
Y��!�;C�ݟ��c�Cf�CVU���m�n��t�a2-HL��FaxRL_)�W�K$Oo;
h:�q�Ѹ���-���)���q|]�C��Ǆ1Ua�5f���o��f,N(��8y�cŨ]1��7r��`���Nٳ��\a깞`!�>��N-!3@�ʰ[ٻ'��R�๓6~\�X�XX���f�y�7W��źY��,g5	�Hl��59�>7P�Ļ��5��]�Z9�</��O3���r��������K���-ėb�Zw��(R�yD��ia�O�7�#I,2�
�Z�����B��D��\4��Z�<F��~�"Uv�@H�^�K;���29m��C8��q�L����I��Ay/������/V�M�����{�_R��J.G�O�gZ�K���-Ľ��}�@삘����v��+d]~��c\��4a�����zz;���N�[�ى�P����f�2�:1��Tf�L�`�GgT�7?j�R�}W�|H��Շ3M%)��J�)��l,"���ٵ��:dꏍ
����]z�<�oB�(�����$oL�� �p����˔�qe%�g�9�DM��)ˡ��jr�y��=މN8 _�5E��,ARI�|��4w��c��Da&^RG�p��K r���5B�4`,a�/O�A"��u�񴶒}^Q!*2CX��,�\n��xn);zb9{ə��Z�Y5���ynƓVB\��w�'�n�I����zN,�~��+ P�M�z��ԙ��I�����_}z_UG �X���XkHQp{=�<����C���O��jcF�Q~�+ßK��T~%%b~z1ks�?d8}���:��������9�Xf����%�b�*��1]�P��瘒Y\�����>�ɐ `L�]J���s+����� @<!�h�;��2 �U�2h�l��ĥ�p�.�0��<�Ok�:�o��8t�N=�с lO@���ۿw7���� �Y4�𭳜����(�,�w�nշ���K�J&�H�0�Ko3����#*�_Z�?�������P�Q�x���+ak̝���hy�7��h�_`w�����:����A3�J7S{.�Y����`�z��t�֭����q�d���~[ߴ�E�A����B��b71�=��x���t5��fre�����Q+�0`z'�#����"=��d}�Ͼ���)-O)��$�r�
{�q�2��t�;E�K��k�Xq�e�=��+�P ?[��_63��Ƹbs0� ����;���%�bg6���[9~�7*� [&J���|$����F���t��v�b1J^ "v�����	�3Y�X,cv&">��ɇ��!��fFvZ���3£*d�B��*�y�᩠;@��h���j�<�0]1��.՟�Z}���ˬ�e��|�ɘ�����Z���7U*��\����z�N(��*??i��\,�q.��ɪ�� ����Q	}S�Ǘ[(�U�p��k�[�ˀ3�5��
\YuA�OpeK���������A1�ơ¤wc��W�x���e��â�������n_U��!>�D����2b:ˇͶ�i
 ��@�p}�˞��A��5	6���a��	�k�΀�>I����1W�9�)_��MR�����SU���ۓ�4��{�G���)Q�@B}����H���(&$:��+6$���oA�f1�ڵ>�����F�5U����u�# �J�8�%�.�|D�+���>�����2W	�X�5��lԦw�?���c�Xe��c���;zy�t��r|��+=I��w�j��s+��~�?�C�#4Җ`t�D��G;T�Z��L�������E&��ۅ[�ŵw��(5Q)�ᣣ��MEK� �|��V>� �.�2���_���F�P)V[�8�f�o0��8�v���J�r�P" �H�#W����I��
����C���Pvn���RJ���P�h5�N�B�9��*eUF|U�G�I�DF��}�4c.�Ҕv����O74�ϒBg��}B���r�ޥFpE�z�^�`�OO&��2����l��Y���dA4�j/�P���k��hՙy��:��x2�4e���Cq�q��~IJ����wR5�4&�X�b��#��+
���C����$���̉lhӑ��DF_,H��q䢕��F�q�0�)��d{�����rUa���<5A�j�͕�7��d��m?ZP���Js
X�J�J��'HZ͖��8�-�'!���{�	mcN����T�i!�Wi���*�Gԝ�;��~�|}���%nu)
����f;~���}�!nIՆr�˿^k�e5m��+:�[7{��L�e��⻻��|�<�<��~�!s���H����)J'8�g���g¦�n[5���/�!�r�Z�������|B���X��l_��(U�v��
�Z.�|0M7��<Gei�ud>5�#�������!~gȔ�O�0;��:i�(��g���^�`��'|V���6�%Ʋ�9�,K-g烕Ȋ��[C�=S/�M�+&"v�9���L'��@<J�/:���]m�t������:;�mS}��W�Mւ�9�tI-�px�T�=���i�g�Co�)� GM�/��)Hl�ŀWq�}Z�@�^����a�C׉4܈��t�I�s�������ǃ!\&9��
��@3�$���k]|��~�J�O��3�3�#�|t:W4H����$�n�V��x��K���|�M���l��5o�D}�����Gp�dlJ�N�N�%|����� �/��M�su�f�	�c��3$�
9�7EyD-b�ZVYb��B~��`y�wf�w;�4狁�5bg�Z�b��cĻ�.��V���`NP�}���x�Yض�s7:�^m�l�E<z�Ut����H6�W޼�h$.���Ǳ��}���*�S�n�MU�{�5�\���l+[ �wD%���a�����y}��}bڎ�7�%X�Sv)i��SϐPF�����v�n��`��Ka�:�����t#_���%� �_#�������
v��ȧ��i�}�^q����0皟qG{�aCG��X4�i%�4�{y��J����vDk�Y��C���qt�ii���n��-�ȩ�\U�ߊQ�`Z��A��%���c��|pJ*���(2���1����IY{�;�2���4%~�lZd'����ӿ�|�U� (��k�`��W���;�P8&�XJ]	�O�.�D�l#U�w�p��'�F��9I��o>�t/!�U9E�2/���u~ʘi���}�~I�kB�P��\�E92<3w�`/j�1FQyx�y����4t$W=�6�V�'oH��y-3y8����$��2�e;�"��j�;ð��?7��Z�-Y�����S�¤�	ZK�"+�e"A��d����GkCZY�#�Ci}�!�W�u��2R�UP�ҁ���[�K���~Ul��'���u:�	@����×���Ҁ�u�5�'6�,{�M*NU�d-S%��勰�,WQ �?�܏�n��(	���ш�*��������l�
�ut�U��.{«�S������~����F�!�$�O�]슈�^�a���U2s�lC%�!6���<�wټ*[�N���&U��lY�Ͻ-��CnV��B�!_����e�^��q�X�>�8e�����#�x�]��j��ʶ�2v�)7MC
N4�>��?��՟:�W��}��t`��9�a�.PH�Q��&4�: �_�>~�i��.HW�6�ެ�4��c�-�͍𸧘d:�aS.=HC%nK;�ڃg��M^o��+kb
-&�(�&r���Q�D'�"��d4VϞ�P~�Z*��B`#�a[�h�dMb�+�8��=Iq�c�n�MjƔ�w���'�Қ��94�gA�,E��_��
P�JҸB;kk 3;�>.����^^��O�Q��^�nw�&'5�}�,-'��?R��ϱ�ʿK����df<G4؍���N��Qh��T�|ԕ��j����I=㫯3.� E���>�SMՀ"p�:�5s��S֋e$�JI�������[�`O�V8Cc31�e^~�>��^����:
K��L'<_���Z!��ud�vi�N���7�"������'P������X6���į�1�E�d�T<_�d(*�P��c�M�*����6-���&�%�� [��S���@3m2��k�c\DSL��b@%��3�cΰ��oc@w� ��MT��_�*H��G���k� ��kR�}�+X.�I����	@�V�<t7ư�4�qp�.��j/��kY�z0|Թ��~d����h���P%���H�_�?�BL�$S^JZ.a��4�IhP�֔�.Bm�^�'s4U3�M��6ɆqI�������so 0hg�%;�o��H����7_��ԩ�.�炣�,��2��'�O���.�7PL��Ì*)�<�C� �נ�'��2�c[|�+����y�.�e���,|;�bb[��H�X?�5�8p�44��F��w��I1�Mʸ>��c����^�#����g��XX�N,���^%���ϥ>Hƶ`I��ތC|iX���?�:s�+)��k��Ex(�����ܢf���F����8����ocV���j�"�i��aKx>W�+�&qt)7�:T�C�7p\� IŊX��6��bU���Do��[�Z6lPϵ��Ddr"�6 �W-�Kڸ/I��#�F1��e��ʹ�\��?G$%^�"F�@P��Gl�1� ���-W͆�x�DV�4˥?p6�h��A�&�Q��LU��RJH<��a�����Ż� �.iؖ��6f j�����?۳Z���^s����C`m���I<��4l�=�Y�Ja��Z4��ER�ء�hb�H��d��f�{��;���D�?1癐�
!ЩLK��\�o��u����+^�*��i�oU���f��(0���]�{S<a�ؒռ���t�%�[x��Z�ڠ�>����!S������ [V����� ��#�F��Tlc���%����B��l����tq�����|Z;e�������h���mBxa3�E-������/".�钵�PW6ƆEú@���l�G��w�1��Q���(��Ӏ�>�/�L�[um��h��b�9�R���\�l��Y�䥟�J�6p�J�AN$;r���[�h���-���B?,�!�L�Ӡk�Q�`܅LXv���-��!ܤ�?�)k�^ԁMj�N])�^����1U4ze
T=�C���dGd�aa�����HTߝu���8�&�b�R��y\q�ӕ���eizy��lo�P�V�'�;�K҃n�C��S����M��kT[��K��&�4��P�����<_��K�s.>Э�����DEof�D������!�}�1%�z�ƊhW�'���8^�E!��S��U�;�G�)o��i�L��>���l����(;s2�s��0%�����M^n}���ݿ��8V:`��Y��'է��F�|/w��i+�H��ۺ���=��(X~Y�		Ժf��F���j˷4}?��/A����*��#����u�l�>����*�/1f�%��ॆG�"�:���,nNm�����H}��oQ��s��ܐ�y�YEn�H6v$J��2o��$���R�`|�&eh�r�>�-���$�����(�����Ppe4iQ�wo��@��1���{�Oq�)捄}���_uI�]h��7�������ٲo@��;��[&�����x�+Cg�S1��ߪ�3�S1��
lQ�.�c%ƥ�����UƁ��ӔHu&#��"����n0�F.�
�m���p]��c�&�W];;�ݗ0��f�%b�֝2J	�����= =d�
zզ�����.�җ?�/c�i�O:FC(ݤ�޺�|3�(M�w�4�4˝��[`��Ӈ$������������A"�Rp
T�8p��Ұʆ9�d��~�@����'镋��gK���&��Q���B�G�>(��߲(���B�f_�����jj��퀁޾o`����X�] �S఺�{�O|�y�����͑�	d�&��)��[�.:��V>��q������>bk5��1A^�*�lOF�[�T�a�]X�ԉ��`��8��}<��x
;����]+Ȝ��>��3����\D�N5�B��@�"����Ff�S��(��Jw��W��+�tq/׍k,��	��S��'�$u��$`⿠�7����i�"z7�����I%~3�,�Vx+�[�s�&��څօ��ݳ��7�j�ta7��S���	Т�e��@�S����2q��CώI��O��^9K2;�g�s ���..���fmFt5ƶ��֔y�v�"� r~W����T-���0�i��e%�o�v)(��*�X�Ҏ�l����y� �I����NH
�+�ƫ-Ұ�xIh�<��1�d�~������ٚ��ꪽ�iv,�����|�3�#ٔcI<��%����R�Y(Y@�!�7�/�y�0���a#�zo��ri��t�vVy�W�F�i���["���|�H�kb�Ӟ)�Թ�FN�����xm�yJ��"��9��4�#��|�|c���-��<�Q��q�L�
�c�4����� Z�!%�:�$_�&4:���>�$&ˉ/������	C�����/J�J�0��քM��W/<�d�"<}*��N�q�l���G7G,L��-�jXT���9��X�E�O;b�9j�E�����ڐ�KmIͫ����%!+T��ow_v�g����ρ��u�<m�	/��2��.���4t8%��$}W&"c��"^�$��L�X��׏7����c���v2�:�:�'2e�g�l?&=��-7x�'�Qߢ���cH����i.y�t��8aӽ�FC�v�K��jz�(GgcA��?-�+��ldj�T2-%��Qӑ~v�?�R咅�ЊO�r�
RI���� R�8�v�b��m3���Ύ��nOyf����޹���i���|g~��>/$R��P	��p����H���K/-Ξl�3���vӖ|�]����t��x��`�������:>�	Y�c��	���:�Y:d��Dp�)x(M��	g��d��k�^��
IV�"����bܐp��_f h��%\-�hC��L�zxf��=�c^�9���H-��E�:_��r�k�+j�3-a{�F�5��&}�O	rJ�Gf���������d�F�����d@���T���n�)���D����}W�������|�u���g����B)$p�pW���O[�u�U�Y��.��z���ݿ�V1�t�l8�-l�q�	�O�.�_~U��P�iϙ��F_�����7U�V��ڮ�	�s�.��9�&<��&�S^�,�A@�����<��״��H���\��% ���_!�s�}���i�_��!x�C�e��@����u�s�t�-)�O�,�i�39{!nR��V��Y�}cR3��������6�Yp��8��@�`7J����{�SRT�
�k�F��}�@m��R�`�p<�@�JR�.�j��A�&;"T�O'Db�f���FN�������2T�A�ׯB�AQ�o���P�Ѵ����l]Ǧ�	�viƶ�È�d��6������`ˬd�I�!�-_�y��t�fV�qE�42�PC
w�`X[A���{ߖ�"W� 	�Lt��� �<뜲���Sqh���soyPj�̸�̮�W~m>Y��N����S���>�{��eH[C:u��	e�S�d�>N����������}W]�.U���$��"ξ�콝6�� ���I?)�e6�8�B+�uD2��y�W�IjEHL���t�Ͱ��$��B'�y �%����.t�vШ��QxF���9˞�ɺE�ۄ�H3|ۏr�,�/�iN_�K��a�I�.���̴ۘ�Hk!��AՂzڸ�v�|ۆ���_&�����Iǈ�SO�X#<�N��XԛP�]8�e��A4?bXA�I^g�H	�n��sG�rr��[F��@�Py���<	���v���Ee��P�lY��b�(#O@�L��"��l��Ʀ���e�� �mQ�GX��}�{�u���B�hN�ԍW�9��������@ˬ�:.����}~\�}��5�~���A��m��I @s�H���[��R��W���AA#�J68����L�=�=UA���m���R�H��ԯ�!�l���C�@�)�{h�)H�f�;Vk|�/�4����q�b4��t
3*UP��F1��Ղ�'���
cA�P��Gݙ�m�������Q�q��|lN��*J�0m�Elp��Os2kb���]۶"��Q8rE"Zn+c�9eA���_�D�5�@m�ZH2Y	�Jac	ɺ4��q)s���j&�+^j�� 	a����gk����C�*K�p̏�DJ�?��*��<��m{��o9p듌�&��E��Z�m��]�T~ɐv�ڃci*�8U+�z�J��`N������� um�)�Ƴ#�r:���l<hj��y��(^�Ʀ�K⩮0m�bͽ�1Fi�f�K���D4Tբh��`>*�^�_jh�%]���H܆����]Å�)D`�H[����Z4�f�Eq�v1��µ�>�갉�ճ�B)0x��L�~���JRX$'jG�j+ҁrI���2���N�������j�*����`
g�f��5לE!�ڈ��2�-�?�n���>�������F�ﲙr5^����a��X8|�~��B�in��X"�-`�֬� �^��aW�`n�AE�N�'�J�l� ҇�3����O��珰��Y�V�.�P��w�u8��UG+�}��f�5��Jrʭr��������Bm/?DA�ι�Z���-��r�z~�%��`��#`>�������D�g��d>�!���07�ңUZ����ea<���aH�ã(�i'`�$�i�cy�J�:<���:��S�J�2Y�K讘G8A	�b�t�qJe�ͩx��� إ�|������$���s8~�h��2]&�t4���U6����4:����nݠ�T�=��$�{��|�NC�/d�q]lTw+�߲��`<��E&gFc�C�6I?��O�6	���W��^D����hˍ��a���&��-l?�o�ޕ�0�po~g�(�
��u�{�O�-y��/�2}�ѦUg��W�g� �������J�(�J$��\�Ӹ���=�ڀ'����r���aozX��'�	׃t/�p@V��rۿ����oV�
�iB 8m?��2����2�3���@�y9R��`�ђ�|�����QRd_�fg�~�*-��"�����Nd���i�.����1������o/ U�"h c��
s�?����3�9~�����+�.���C�?�2mD#6�R�Y�C̽D�L+�\4GO�x�LM0�J���f�:�*��{�Mo~�N�c�j����JO/�L1��Vm-g��X=d7e,;��|������u�J��R i{.��r�"S�B��Fl��~3��ڱh��	!TbEmf_�7��$�3�b��n����>-�=G���u�H�͊`X1��l�uA����TY)A���AEc�
��D�:H���w�I���%x�%0/��	�-�x���-�vU���Ѥfz+���t��8����X@d.�3����r:\��=g]����0��<<[�_ek�.!�P��y��TaIC2}�����c�&J~�cF-��܀y�X�.WL�E�����,F��q�O�s�(7x�M/��I��z&DK�^V]Jܬ+ "��'�����&��K"�F�j�����i /e�懘$���NSW��fr[[��/��\������ 1�Π�X�=!�h�lҜ>GU�$lA0���V�7���=qz��¬�dǰ��׃^��5����#���wG��#ө�2W@�m4���S�5����C! B�;cU�������4��VO;ݲL�d���">�(��  ���z�`>�X�@�i�p.�����ʩ����i�0�ĸ��N�;쿁	V5eyܺF������}�'����&��-W���3F�,7ZQ�u	�S��l�����}�W���HEA�/\XH��¹M�/5b;'��`��/j����$��I����=I��(�Km�I\�w�
��]�`��,�R����Hi�-h��u �hX����H-�:h��Y
��#�~x���[!d<�M�j�o�K�p1�"[rRʨG��$�r����������[��se����c���x{&WUhI;~��ބ>3ȝE���ņjE��O�QC�ks���X�W������V��\p��r�Q!��(�I��ge{.��D�"_��-��E)X�c~B}��������QA�:\�3~�0��Zڣ�Y� �_�h�����O����_��(�z�Ceu�9n].�]qs�UB!���	\�q����oM�� Q�h���S�;O3�\Ol� �~rL����E�����d���@�q�ʁԒ\~�i}��L�P�&k�� e����h��m����e8-Ӑ`����3��|�M"��`;�����c٭��_(~���"��S���+c8�?�ʅ�(�q觯*�[����Ψ���t�>ɐ�St�Q�dW9y��؞R�c	�M���đ���q�H�a&�����kj�����D�E w�� ��`�܊���_N��㟣��+=��A%�a�"�X��N��n����k���%:�>	:g�r�Q�6_]��̝>6�X�֟<'�o�MJ�ʿ禕jB��j�k��Ԇ�<軧d!���g7f��h��s�A`�0����w�
9����APEm����
��ߛ�C��8��/&C(�CA!�T��8��M���ꏸ����/��T�p��G�����\����&��D<�@�U���8+z��Dz���p�g�"�棠�����ɸ5�ݚ�U#����t<f���锆8U䪻	L5@�(�U�*��0�F���S����H�W��&E(=��z9���/}���z/�$pb�C%�0OT��@z�B�9�T��!�m��v�h���l�"Z4�*��[���E�8~R�@W]��������rH�3�/��WK�>3e�>X	 ����v��ox�֪n�^��ׅ�j::�Yu��<���R��L>_����<�n� ��ӸNW"R=���*��?<��a�Pol��j0��)��"Iö%������U�s4��3H<t(�E]y��	�Ku��Dq�7�n��hS(;ZM�$��/gο�J�뙎����CE��d��/�"?����S]���c��\�K�5�>��P1�=��φ��HrD�K�N��Ԡ�ͪa��KbT��1�T����Y"�48�Z��P�J/�G��gx9��4y�0�I�w{U־�|�!W�9�3q�F�A ����):EwxJ��ꎘ	�J'�+��_ϹLq����,�Zd▭ɣ��"ɡ�N/�By��Q�UJC{!���t/�BFK�ѯ'�|+������f S�+�+����\�5����R����@_�e6P��=C�	&fDw��]����45�N�z�dË�P�(��	��>��t�g�E�'����zons�S�18������I�5�x1�%̶��w"i��g��w�hzr����1��J�8�5�"0����1��*H��㒽�P�`)b}#+[6��Z����*n��u^.�L;	��tj��d:w0�m��2��~��B��m��WMa.�B��UԇV�	�X��
!H���m��Y������*��O�Cn�m����8�DG�|�.�(�Ve�c�m��g-YT��$�{U=��g�;���t�����Ȍ�������wa8h���:��Oqx���#DP5�͈:�[d���ap�A�=L�C���I)��oa��@ú�1�W-�֙�ڐ�-�>��y�$`�>�/O(_�P�wT�4�Iʩ�*��˯6�-5��@(����v0;ޟ�"�|h�L1���O:
�M���u��Uqr�>R��OMK%��Q/rC?3�l�=��!wS$2��.����cm�����8�p��D� r���u�/�I�}�f���W#4Fp�&�"��.�D��l����x\Đ�J���g#t8'��*(��S@^��k(��Je>�9}�m}�9`���[�*)�3��Yj����P�������v�*
��[!�Fς~��!T�$q�:^�j�!��Cg-���B.��y�/�!�rXWv��~Ye��,�<s�.�sV���U����f����	�;]`<z���pC+�h��:�S�'kv�x�w�)��\����#3a�rp�'���3<�Oh/X�KO�e����#�:Zm�4��������+Qo�f�)Xl	4��|�����}��:ք&�I�9SJ�_^f�W���Ĥ�����Xl�+�	���[u@�U�E{�)x9��6�刨��<k�u��m��ڍ�NO��AЍ/���-�[P:v�pD���V �w�L1���l2�&�����(�4Ns���Y�"E���=q
6);IBX�9V'�'�F-> x��	�Yi�L��̛}*2��c�F��N}@�S�T��b4v]?�8�K�!��l�?�EkxP@��>M���d��I��ˮ���ĵ��9[e�����|�c
�lx�Q_��G� &�7%FǱ(��h �s{�#_O�Y���?�,s�ՌC�3��"(��C����HaK��:V�(/���d����/�l�a���'�����t�q���Qd�N�M�������k���#��=��(��8�5�	gH�"��*_=��!T����[0eW`��7C{�,�d֞|f�w���n�?�S`�>���{�1d��fg���p��SU
�O4K⟜�c�ˣ!C�-4�U��$»�|�M�K�{�ȰT�ћb�s�3��֣������\�E�W���+���/�
RF0�lZ�x�*��������&��zE�^\�Ϥyk���Q�ФL����V�Ed0��~|���x��,h����!��܍����\� �Թo�w}�ݵ0d�}��E���L�/o�Ӛ�X,�if�Q��Q��6���GJ�ڏ|a�����ٓ�ÔaFI�3X��T�f��'�߲��	~��:�:�	ìom��AKa���xZ��h��"�L�OFL�֣�B�����$$Ԋ�g�
}����;d�>X��}�tJ�� ��ٔ�na��՚t��]�r���!aW��gW���go�l7����N'K��?�&��<2Zl�o9����d�I����i�&�L 0i9����Ue���*��p�	w��L��Յ���Ts�!`���k��`�����0ϖ�$��0�4+����|F�e"���׎Ό(�mhˏGd��K�~��B��"e�F�{@�0h�仪:˭����Y5�(���.;���%�/���F����i#�Npe��<��������}������
\r�O�􎃸�&�����K�!]�}kS��C�[�A��>��Y�VKj��iZB����8���YV<C��J�IÛ]�A�=��\��	��KϼE~(b//���e��	�w麞��׳m��X��XӴ{M؃ܰ�B��� /9sr�A[�;�v�'e�E�6�F��٨u��!$���L�B��iPqȺE1���6�agmϊ�MO�w-Y��8�O�b�y�v4�b����*L�tl�sU��I)��j7)�WF��7�Gtk����9J�Q�+�+�wՠ6��D�~����[��
͕�i3s�����Y����~ž��H�֕C�dy������<�V"��"��'����W�������GjHD�z;��
��.">?W�D6��rPG7R]&��b��� &f�z������U�i�a������#{���%��� ��[�9�D�w� W�%��Dl%��veC>�Y,��R�� ֝��7�{$
�U-�L��z�����E���D��� �1����)B�n#�����
�9��J"���l΄�P����� �C*fz�t�@~�� <7.������=�%����,E��z�v��[�;B׬���U7������c���� ��7-����j_ĳn���A�own���3��˞����[d�	�hms�k��e�[�"����Y�w[v�v��x��BV�%��2��_����֔7�9\����6� a�m�h;Z6Y�p�x��R��Pݑv�
����~3�1w,�֢Al��
!�~u�� �y���{��OB7��?��~��6W�W�nR����.�_c�a��ĸ���\ʨi�l�4I<R�hF�qI|�滆�6628(����VahL����&݅��wI������bKZnn-�LQ�_/��EZe�#����1!���I��&@BJ��y�l�e�����6�g���=�/$�ڲ?�� O^J1� =o��[���,��O�>���"��\1�Sw0n�Z1�u.\��p;h��ǩL=�W�;<���m�]�왬�4��3��d�g�zJӾ4Dy��R����n�K�lS��,�u���Yn5̐�am�5[�����:K��$'lג�~�z��OǪg���z%�Vx0��E����c���Ո�B�L�N���tFɖ��/�f.�p \�:���'"�1��~j���U�"7X�]�����{��Ƅ���`u��n����&9��A\a��@�#�b�j���C���$nrTE������D���d@\�#�=\��U��?�ٛ�2�P�S�;�Z>S;��Nkq�j�X�)�����MD>��T���zχ��^��Lnz�OB��P� h�ȕH�Oy��jn�%�k����R\%�-�B2]
�����Ǌ�9���[����`%c��z*hQ��OT1:�!z�c�@�?�}�E��p�y���GC��a~ó5*��I}�an� p�(�~��2��,Ae ��0����l2I'Hż���s6D�@%���R�ݨF���=�z�"9j�+�H|��Tx�LZD�O�d�gv3��N���zG�x���(C3W�;�[�NF@0��W$�+�;&�"겴���HKW����R�NR��J�BC�u�f�8�ॄ<��`��V�4�V�8֠e�V8EsZ�Dԧϴt_��2�
�xVF�ǌ���ٓ��ufrX��ͷ|'�%r\?]��Q/a�����c�&��HJƍ��\�����%�=e����r�����_*uDl����s&'�:��J�n����.6q�J��P�٘F�:�t�w+>n��>5�������R8ӞȀ��"n��~1��We.`�!���,l|4�@6�b0�mv/�A�?H�6����伒i�5�iƍ-RY�)���wK���i$�/k6�0�Yb5�]�K��`%2:��Ҵ@9�E������`����I��|��,� ;
J�s*��pK�g�ۼ�� Rro�*1��N�%d��F����aR����ܣ:s�{�h���0���PYO�e�R�>�����(�·�hvH�X̱�����C�]Y�� ��"���RgNѓ�J�P:����`k�4���)��������īu!f|><�DS/��l[�1��۹�ǫ��Y����K�Ԇ�G����b9C���!�z;�:���8�z8IHd�c�<-�H5?K�G�386q$�D��*������Kt���\M����9���=��b��riH0"]����R'D�1O���)�F�v6Xj�:x��'�AuF=����� ���@����� ���^r�%4����l�D���LG.�Hq?��J�)�2b�Wz*g����|,yK���&�����w�$����χ��ҔM��U!���Г�R�Q΀TH+�)AK�\�����s���έ��ȥs<�w`R�n�: -v�k��"����NU�kD�ᓧ�ﮎ��<�Φ��q���"�25H)��Y���,�k�ul��Ky�S��˻�����*
�q�N���m��>�N'0F�?=�pK��V��n���� ��1��Q����߻?a���e���b��mZ:0]aoґf	4y�B�hbӉ=�^����	���eorO��e��;���2B�T��4�j`�Ol�r=X36�9t88��|�4����CЃ#>�"�%�.L�]�x��f'#��H���D����/⾙�>�D�#����7��i ���4&,��Q�
Qrz�<X~�k���d2��F½�E�6�B�]��p��Χd��ļx�(����ͷUҔ}T����G�n�-�e�X-"���n�d�LO�Dˎ���@��Bަ�̝��w��/�&zQ���LZ���%*�U������*	�W�b�c4��9��\g<�iI�����#����旛^̈���n�V����
ߺ��z�7�2r�,>�&8�g��)�d+���i�68�����U?k�Σ��F��!(.�[�_�i̯Ğ<Z�m6+�<��)A�5$�ن�ح)S��o�N�Y�I��=V^�*�������{O�CtbL�����?������L��Zi?���2WZ v���D�(g������h7�i�"��������8a�5��0�+~mr�b*/SX�bT����c~*��J�t�Q�ˈ��w(`���k��@���|���U
B�I/���/]�Y�k1g��5 ה�T�_�h]G�9
ne� +E�\���hsv������9L��C���dr��*G�U=]���ƈ�kY���o��}Uo�I(a�6��8�EF�4ѝ���P�aZ:�j5�g{yuҼ�c�ϳɗ�˝A%M������7�|j� �L����wY��X:=����t'��An<��դ'z��T�N1m,W��[z�kUޫ�`�I_7wh�U�A���'��
lh�r�=�~� x߹�刈��'tͩUv��K�g�{ �~C􏤢���R����������$�a��㲉'SN--�0��\,,@-y�Q����/�%Di�E���, ��?�m	��&w�u��^��2�k�֡%^�]u�	�����'����5�{-�)�%�no'a��Tޣ�hAB�VnZa�b�0`W�:ג�+���ͭw%���>f��6Χ�d���L3mIk` So3C�M75�U4ԽHFŔE���<V)�J�,���`'Mc���H��R�\�EM�uԒ^E7���T��2�$3Ce�$�}c�0�!a;[��!���4lG�+�g�Τ-�B��6R�f�y�=z:�����ɳ�Ek���%��[�D���n�j����T���r�O{g�%D�� t�7�/��rz�G�ɝ`U�B!a����@����)���M𤓡�9�6w���u��]1�ړ�j��}���2�'���������W�Dl�$��M�a�D��q�|�n� C�f��/�8#�8��B�,����o���>��^�am3"����;����LF���$t�(��>�V}֌|���=s�_.*��K.~=�5A�����~.�=�K:�r	���	Y��~Gp ��B��y�B�(������ :����7S�ɭ�)qk�`T:/NG3!63	��⊅\�	�X�d:�X+kû���'�g7�R��{~�����o����vu�Dҩ�9q�ٳmt�fћ4v.�/S�tI���4�R]א�X퓋��]
LT��hf��jӥ�i��4����ƫ�2��2���f7">rm�����G��[���
�� l����'4tmi{�!��_a�)Yӊ'`p��5Y2n�
���65R�����q:o*�4���&��v�O�	�gkL�]G�
����		�<�U�����BVa35�vS��+EXP�$N1;�N�-����%,��� ���X�Ń4�b%QiVu�St�����p��𔏾w�җ��|�i�i:4��܃5�`�l؀"����A+�HS����Y"�ǹ�x����:�V�n=߮$O�s��%��{J3�ې�[�\����ߗ���ܐU�Lg��dT�G9�G&k��;�N񐫶�$bP1q�5�X��)��K���b"Kf!FP@������1�ĵ��WB��?��U/��P<�1�1��+�.ʪ6�>�Q`��4��H��mgwr��:�VT{)eߟE�m-�헾�N���ۮ�i$%���ؾ�ែ@h�w�s�tUw+�W|��YAXk q��ɗ���$%��ƪp�^R���+������,�(��6��cR�1oj�^��L�9v7�����[��[�ܞbJ�\+H�{A>�{�k��~h��'�;����wX<�������~��d�ޡQ�M3tñ���ǉ0�*'/�M�mh%	����
���i�;o��BR�=��/��� ��Y��!N�>nÎ;IC�Ҥۡv!]��-6�_�w�~����l�O���� ��qV%z#�i�k\�7���;�֚�j�(`	�������Y1�+��-.�JX�x��v:�@H�S�D�??�~þ1�ܡ���1D��uO�![bL����{ׅ���޵��}���f��&�� �s��=�x*���̓Uv�#FɌ�VE��T���W1.DXͽ�6y/s�l�{>���'i�V��&��d-��o�ʁY2td�g�C���Du��h���ngWs�@��貄��Xg��0����GҏZ����x@H�9�Q��ҷ��#'H[�� `bSN]��M&�)��5��9eΌ�=������}��a���V�}/���KҔ�{�֩�2k,�ѳT>dxS�[Z\��aWJ[)�K|ۓCv�zڳ���k7!��M��=���Le�V9�D~�bYb��� ƄM&Z�s�|��N�����No@%S��a7l���K0Ygj{q��n3��_\��߷�Ԩ����i�0-�W�\�K>2I9�
j�ͩ�[�Krtc��E���=��{V Pk�zXa4�$6a�
o)���1�(����=7*�L;i|���*�k~�"�~�>��[�vry.8`������A����O]y����TKv���{���a���s���	�- G�a5Z�De�o?�2�����"� �BK�8B�Mz@�M�zƅۑ+�(W�:���;�IJ鍕�E��
��U�hݭBE�9�);v�m+�n���Wh��4�2���KwA0�3P�y�w/J8X*��g ,���"���U�1-H�
�eeӗo�Pb��ڳ=`B�w��Z�{&{�v!g�C�]�O} q� !�N��Ig�H�^W(�����K?-8�_H���>H ��VVՐG�����e�`?��|��Y����6[��=���TRՈ�а��l������gyW,H��O�{@���m^���Etq�P�{'���6���3+�D�����'p7�A����I�T�
���j?��n+��l��l̩�:����,.���Hk��t�X�iz��S�{�ML�f�~�ִQ|����Z��ޤ�1
-�6�e��2Ʉ"�`;Fvi���ܦ�m�~�ˮ�M��ͬ$t��� �D�	���&P=/W\'���	����$��Y�:�}���Cʘ�g��9T�s����,��82@�U=��ܳr]�K�>��� j�ZWq�\��%9ﲣ/[ҕ��MrO�f�Õ5�D�uـ������(�	���L�v�4��N�V�GvyG�G�S�'�)~&�Ż)�j`j������H�4�f�����<�'Չ��\+�'�����qH:�(��ss�~���pe�k�� �{T8������.��^^�)8���D�ßP�w����d)*�%��)"�3yn;,z�i��ܬ��6&�O�B+�JK<�t�~������/�iB��\�ĺ��%"H8EU����`V����=A���l�o�j�e�,a�,O��P���;ϙ	�W(����am���D�-k®��.�?�O�k5����{<�@��҃�]���S�T?2�)�������r7`�7ЄæCy�I����I2o��Q���x)]""E��u!�4���&�C�τ˶�\a8aN�lK���_�Z��*&��ٞv�m�Ʋ����X��׷��L_�F�9ڲd��l`;�|{٠)Py���Z<���6�B�A�M1q��E&�=b�Cg/`ˬh���%	�Q(�o��:��eR�fPg�����l���#�%�OC4�.�RO������+N�Pb+JuB�59҅ɷ��E��;o����� ��#��|L����V� �5HNIג�>�;��o��̟��A��F��c1��eΒ��^+c`��M���aRd���ĿW|�4�W�+���@jV�8LM�}h3
�	m_n,�C�FDw�^B�Ƈ���qS�
���P��S���{At���:�N��H�1�h��z�K��5R#�au>�Q��9����o��[�
ir���{��β�b�4�I�ݘ\�x��蹞��,��
��`��H-���������Z��P	�O�k̬��Տ���)�[d[�_d��z��3YS�~��9Ia���W�]�"��v)X�ր}M�̽�����'�#Q|n�Q�IC�� �o/�,�A)咏���ޖ���cbO��K[�>��07fmh�E.����M�uVlEWa�!1��W��"�uqm�]����#zCy4��hU�XW�j�� ��V��QV�C(f%�߾��>O�v?E=���Sai��5Lw{��T蓦�b�������N��ps�]H�;��~<��1���ג�'�^oM������;�Q�х5��kh�Ӛ��u8���.�t��4��CY�MV�'2Y�6����u�K�,N�Q���'�Jg��p°6z)V!6HހE�!׻R��'�=b�A� i��t��}�6׮�|K߶ݫ���p��-;h�[���+�pj�j}��am�I^�9-���گ��W�wS�͋s�(N�	+o��s���8y�7�
�f��6���ų6���|EH*kX�D�%i��=z�GǮ2ʜp
:��M�>��7��o���^n��N���i}�~4��!����VE��� ��I���z2u^����x�0����j�=�#�i��,!�&c�j���PWz��ZR��r�0�W��Y���ch��
d'}1u>�1�8a���2��J�9E�՘�Z�{7�hg�wIo_r�n��R6@�����?���3+��]#�<l�<�p��]X �9�Q�$rm#�r�H��?�<O����JS��}�č���^˫g>Ί�����֠|G��%%}�7�rT�SM�QC?�BSa��H#E��Y~3O�_Б.oe\�X�חʵ�V�C��V���(����St��W7�������/���h���A�"-	�}�ݳ����'��9���$ڕ�.&+��3�TH:��.CސJƏ����� ݧ�u:<fs&����"]|��D�͡EѺQ7��m��!%@��u�B�,�g"�e��E��Tw��|���L�4o����f��-zBdp�uM�@͌��#�.���/�Z�o�r�����5���&l��[F-,(�3�Q>�F�֗HY�����jx��̃��}�wGeӷ�_ú~Rd�&��y����s,�]�쓦@�~�� �����8��/�d� iF���&)p��6Z��@q�+-�z����L%;�怹��I��y��9{��&�і���Km�R��\�I��� ���Ml,�+Zn;$߰�~0�(��]�k�`�N!6�j!��
�H^GQ��{,��pz5آ�'�C�'���Rw�O Btz��`4��hχ��Ǥ��Ȩfm&E�OM9��O⫆L�����tޏy$+w�,�X(k{3����-�m��N��w��������f�݄3�ߒZ�(��v���+L�h���;�f0cw�S��}Q�^#�a�]ѯ��ht�}�/b 4A���S�u�*VpB�m�)?�� x�8�t�z3���M�;��\æ����x�g@�dP�A���<��ߌo5HT�<��t��V� �����2�+�����;�S&Z$p�&A��J�����=Ćsͷ����z��\@M���b1�6Q|�8�֞�O��r�kI��d������l\1�H���ހrȝ�.��ћ�#HNkZ{�6YK����S2�b�ˆc �.�4B��b���r�l�v�Ի�"{ɲh֋�&����^����s���$��%��gy �JO{}��*��[�3Q�V�@	m��G'M��ј'�W&�N;J��J3f�H�").�`��G�~��*���g>�O��la(pbe�$��Y��h	���M�,�ZdQ�'�HPy����$p���WB3\@ıD��cgR���mj�&կQvNz�� t̄��Ug����#�$�zcA�%��bFP���T,�~(��X(d�#�F8:�%ۓ�����x?�h�V�-<�����]n��D�R0���G�៘���d���h�K���rR�0d��<�=������'�ãk.��\�����Y>�����)��8.����q~. Fp_F�7j}�#c���%c>��D�ggKaR�be��-���<�Hw04θ�&\ۅ�oW~m0J�Q�&}G���lЊ!����������	H�Ʌ#ILB4���9�?>:�^3I�i(A3r3)�1�9]>���É4>7xzC�5���:���8�#�ii�[�jlVR2,UԡqXGA [�ț,k�^w�ph�Ւ(�\��N�{�C`���F;9���w�$�x�QX��;LV�ǬPr{Z�<%�(�l[{�K||'�Bʜ��cZ(��DH�ώ��[�Y��ن�(N�%;W�)K��v˄��,�!�&V:buK����E�	�8�:�/2�X�<L����l�n�*�i*t|��T6� v͂/h����I�{wؗ�0�L����}AE6ym�K���f�$�t�������M�~�<Ok���Z����j�X��!%S�]mN��Rv;���,eɁ��h^���!.�W�8��,� P��<�
0�o��d%�Z�:�`���|]sBfb��%Mn� �X?���ե+>O���V�y�*�ԃ�X<��z�;����[��3��(�y�� ��
���x����vE��u��քk�y���A�	�4���̣����ha�	v0SqN���Ck��߈�7_X�I�ħ&���U���.���ev�
�4��!J�]�-Wч�>c��4�ZkS���택��(�� ~�{X���,+�x�-�3�Ø�,�Ȝq�u/�䥬5��N����[�(�j��˞b�@�^%7�b��yD�����sT���\��A������O���� ɵ�{�C G��|J��@��s���^<�T��=��i�d�z�~,�#�C4 5
�OKa`�������[�,@,i����>�z&����Ìy�Q��Z����:���E�����a�`M���UU����j��"
zNb빏)�\�O�|�����P��WQE�V_�AP!�mB^�8:��2K)���/���� �]7/��p8��A��H�<��Ǵ���br�3*ҥ6
��WFa��T� ��e��V�yq�w.2�n���~YŖ��~��(z)Wv����m1>ŬG�;¦��c8l�Ks�8�ؽ��"lJ<�Sh��^��dօe�2�v��DF�F�^9�w�DOb���$T/����u�by�Z�d:��d>�)��A�`wc�Ģ���2ޅ�c��&�X�j�"XP��W�Eΰ�t囆3ZC�vA���Z�&�2jL�T#`n�>z��i�@��E��0�Q�Ww+��O��g�J�l/�������%�Tb���j�)���?�Փ��r�Jo�����/32����}�HgM�f}�5�ś�Y-]ED�����r��G|��ciyXo��O �RV�8D�F�<7����2�Ά���fi��+fD�S���"[��y4xZ],� �b��D�F���|��$�܍��f�cfsw����%�AR��hхWv�Q���"�ݫ��Էn��ڷO5Y������#�=�[X���o�#Ej�~R�!d�a(����^�' ���*��wLO�r<�Z�B�F�8���.k�2S��ؿl�#s.1xP�m@����ysI��<
eG�������;x�"_��x��3�Z�q{����:tdg�x�+��6��ek��Q�o��a�Q*�t�v�k�V����}k*C�'Lo����e �^ӳ�u�P�z���w/�����[�ɥE�Y3��7�fg�R\�6c������"�q�T=���@N׭�5���O�J��U;؄�c�ѥ�BͺN��� �j�����r���jPF��*,�uv��f��LqKzq�����%��O��	8�"t\��=KU����Dȶ�$�����n�f�$}P뷶00�ْ��1-��i��5s��f���I�����!�� r������U(:(8�{`z�Ѣ�KO��J��h����:T�S�%�9�F^�E���=��D�����YΌ�aݦ��U0;p�&�-Ws�)����5U'G2����'�2N@��X"�c/�5� ��/0`�����Q�>��)�~5�NkyM�֡L���z��*`p�ɚ����Z��Q��{����<�����m���>.�4A
��p��oc��_�v�"��ut$���[�ԁ,��i"���'�;�SÙa3I'4I�0��_M������>LOX�p`O�ɟ�'�^+��p�fji��{���G�V���ʣ� �����-��,��h���OC�V�%
;T'P+S���9�LG���齐m�[]�n6'L�SSC�,Z�>2�Ta�~�=�ܾpS���,����qs_	T���&R�![!q����x&x��̆�*�^C�5��8)C��T�G�w3���������ڔ�Iv�U��h� �UL������Ӱ�&�(�p��ٲW��k� vi�1�U[��?>�V�;Acv��3Ӄ�@Yِgq�$����`<g�F�i�4Bxt$����j8{���9RPľ �+ߪ���X]��Ȣ(�	��̥w)Z�R ]�E�[�]���4��U'δ��;G�tC(��`��(1�9w^Y[ϻ��EP�E[�/<��Q�+���^T?m��>�Q�t�ޯ�'�s�x�
;�/n�RD},qݾ�AīQb}*�z��w���o��E1���sDsu�f�����|��8��~�~I1.�$SO���&7Z��V`�u�_WL4z!�� �׎�r���c��|���?���'�}s��?hc�USsd��=��f(42|�,���n�G��U�k"S�~!!̟0+k7�&� ϰ<�*ίn{zҮr��2q#�����]��=G����g+.�Jm�.+�,�~���:XDkz�Μ&l���e��8 F�@MY9�݂6q��&��hS|��SEM�åZ�s�ۡ�kS)ȵ��QLx�P��`�mUa��G�H�o^s��4|�:���A��?˫�<"���u�5uSv}D�H�
������*�a���!'�g��ޭ�&_S2w���aG'���B����,�uݬaL��@�����}��c��uG�psX'�����������^*Eb-���L���-9@N���wa�+�@�����"�\/�.�a/���KK7��,��ے`����q�?���.���?GN��Yo'�������O�P<b�;c�L��X�F�o`�ˮC4��%e��D]�w���?L�9�΢�w��4������a�����Wd��YR��7��me4��j�U��ؑ���i��A�H���鯃֢|I�Ѵ�}3�Ӓ��<��S�>6̀\�5�iAr7�Q�C�)_��o�L9�ۄ;�����z���Þ '9o�����ԣ�:��K��t4ݎ����s$c�� P&��cީU����aZwZ� ]��")��q�O����f{�P�,Ҹ�um������4g�������{A&6y���Xb?[�$%��R�)��K��	N�Q��x����qɚW;=����~�rpNDoq�W��r��m���ȩiQ���KѠ
fZOЋ�A���	n�;�5�5��~KΘ`	UĶ`�f��,�=����I�Ycb���?��E{V��_�@�TT��ѫ��1.lb�"���������ÃiA�����d���5@7��X��H�Iu�����ߦ�����FS�if�ȕ���Y�_YTʑ�Q+G��yTi�W	O� ���Q�52F�L��S��b���XL-z��ʟ���f<%�M<r=zH�diZ���~Yb���s��&h�֎7�q��8��Ҽj�D潑���E=����e�"٩���DU�mv`S~�L���f��S`lG�B)ѫ��jq�I[`
a���>�ۄ?pFl�/�tԆeX�HQvK���Lk���'A� �T�3��.>��~'���+8�e��K}�ԳM좱�<��bT�5���k�(������ğ$�]��Bq�F`�c8��z��)�ꋙO�f`iM,�r�T~|�D�ӋEkma.`���cnNT��w��;��;BMb��u�G"�-�%�(x�5C�$��T��~�8��}�Ք3 �q׉����d��#[�	p����G��W�k��VЋ����}�m]˗4^O����sђkv⇛�A-������j�>s�`�
5\�f� �,�B�c�@�T��l���|1irKn��V���ߛ"��>ډF��F�'���\� a%��´jI�2�r���Ɵu����腤x�#��e��jz��~�0���CM�8/�p�v�ּy�{R�8�Bߠ�M��*U!����Zrr�0['d��9�R���ki��03��]����H�K%�j�Ќ��Q�|�l��Sժ���gv�j
)|��@`���KTZi��+9:�:~�E�\� ����ծ>���l+��=��3�Ur�.����!沜����{�j����+����ueYP�M2��R�����D�ݟ��3 �qPC.�hSY�Y��Ii~�r�t&$�O���g6+f@��M��Dõr�4ā��%��]x%^�
�`qb�OYf��'��rf��tп�w�j3��S�O�bc�9J�8L8	�HC}7.:	����-A�B��]�PO��{u�i�ɜ�'�6�[HoMj�D�/�<���^�m�b�@�:;M1Ȯ�T����)����w"�
�����6|H1Cν
��sG.c��6�
䝈*<։@?�_�*N���JM֫�g�a��fL(d(�?`����`��ihk�mJ�4c���gČjN����2x3�
�ifh�͕�cbnx�W�ɲ\��9�G��L�c�L��98T��ו��z�Q��^�v��~I�Befj�d�?-?��۞�"Q*�)��S�rx-zb��b��.���z��pi"od��`;p? Ĩ)H�֍0L�V�#��٘N�:�/&$p��IN�s�����uZR�RP�sX���S_I���L?���^�z)���B����]���Z֖647M�>�ɧ�����P�qG����y�^\��Ԇz:.Š/eGڥz�	�H�#��Jc-���
]��1�Z�}CCMn��!��t��]�>+�a�>,6�)�A������P,~̀��̱n99!^<F��� K�F�H�1�5��[U`ZmM$�j��
�B����^�m�Ig��s�Vq��	�t��7K%J��Pn�_ڇCC	IlI�0-t�JI�����,��M0��I���Eum�.�>�����iX�tc�m"��9Oo�;��{�M *�0.p�_[~��N�3�G)�Ԣ]0H:�eQE֥lus�!=���K|}����\�@;�;�A�����Ξ�>�l�V����'h��]>|~�Uz��c��j�Z��K��̢iS�d��y|��~�^m]U�	��]�z�M���q�{O�bw-�O��a��Y������υ��4���V-�R��٤@�j#Ӊt2S�ݍ3�\w$ʚ�Qb~�8wLQjI��bt�pr�Й�^_�s*#}u��e����ױ�`]Pi��у�fs�/��F�u�[Tw&_kW�<����R�2���*�܉��0��ޜ��*�_y�:	�A�����ɇ�lA1�r�N?�YfU�����Yx�;V�<H]�i�H�=�*Q�8X=u���\�ǣe�u�!��0�[	��0{�2~��C�A�%=ﱲz�Ď��N���gL���c����[�
\r��c7�M \��S�^����ʦ� O��!JG�m��v��h���`�3#��@�9��j���T4���hd����΄BZ���W<��q�<[�H��U
�YD-��n�=���\=y��Sb/�*Z4i��"�B�=�C���K���*��T���6�M䄌K��.q]�TV���R)�r���؞v�v��i�d��x<E]os^��GO�E����j�C���p\(���s2��g[�����p+�,�������m̛�Q�-zN��c�6=�6 ��
2$J+N���Z�r��[�7"r�b�~bV�����)۷�
V�WڝTگ��[�>I���7�ޏ��9��b;�`�+���v�?�]�Cq���Z��@�R�bK�P�mhg$�	Ld��t�Yr���̭� �.�iG �ӫ5]+�^��Q@n�a��YS�j�^�a����"���i��"^`UT!N;B�/J<��ߪE�/���?[o����d�g	3��� [)����ϒ�%e����.y�ya���2o7�4�,g�N�c�>]eD������r��-��ULW����ak.��!�uirc�=�AfP^��9�8JW
G�%�F?�Κ�9�ߢkmo��v�&�W��6��=�����f�[�,ZL�B����)�C�:��{�+1e6a���Xٷ�Q9E\��^ �ud���-�݂�)��AZ�0y��Ү�8[.�њ{�?Z���zgt3�oզ �]��xt�e����(�G�-Ŷ~��9'�Uo�1�4}��RwT��6��Y���H��Y��I�֖�N� ;�B���XB�LcSPN�F��/�G]��Mv��i�,�G��`�u�]���}N#+���Qa"��f��AY��Bv��)�t�9�����v��ÔL�qhD��B�
������y L�]�W;P����N_�|�I�XKcQ��YY��]T�aC"2Pg�h��F����+�W��r� f� ��H�������q[󔺉��SmK� �Ō����6i/��j2qݝ3�*m����c�;�&�waǃ���s�S��.�oa�x�Š]��u.�0��^Z�{�ӏ�Qaӱ[1�z�ր1���\��`LIe�c
' Ez��&j%�s�M�]�ϱ��h�����t�@�~�{J,��($UK�<��Z��Kp"�'�g��+�qq~:BMK�&A�0^�V�p�4���pQTd��q��	(ƚ�>`��H'7��x�,�����U�V�_hD�zX��4���狋|e����n�aw>Ȍ}vU7�֘a�>D�K�x���W"�9�Msg�~�$5n�Hp�N�NI�ۦ�=@�5]iq����	H�$�����P���60���-Շ}	�?�ft�1�v>��ś��<�<kE�WI�J۬��Z��S4<=&H �(�ա� �\7H��,S%g�=0b�ɹFM����=p^:|!T���x߷���P����W�}��o:�;�������
i)^�`c���� V��Fmk��j䕕֢�P]0;���!3�2�H�ֵm��t*qa`)���v��*}''$̌���;��~���_������2ie-��lྷ�2S>6R=�#���v�^�V�,�h����މ�
��DN��\B��*��l���5�mv���� �F���� e��J}���^ n;�>ݻ1���#�8�����ҙJtVA��2a4��]-^���\y��eR���B5�8�9�~`��L��'�T_ sH==�#�r|�L�ؘɵ��r���� ��.\�W_v�ҩ���T�u`��vnJW T5>=����X���[���l'g�W��]<�؃*�Y�:yt��O
��~	��&Ӂ+��=?׷n8�^t��%�]�{���.�M���s��."�	�JM����ƳǛ�>�����>��R�f�c-�ٓ�=��)����-z_�5���� �/Q^�&f��(�B�ya�e�.�.	�\��k�6n&���Ug� ��0����1��J��V�h�?�O��<�l-�P(��U�1��0�:Ȩ>{�M��t�7�^՟��%p�f
�$�7p�l����0ם��ٰ��ȱh=J���ޥ.S3�Q����X�E���2�X�8�|s�rn o��u&�F��w{4h�Ұ�Nсr�[0�}�A�����m�D%¢���֙oD!a՚ �HtE`�$�QY��D�30[���(���$���������Q쒯|<�/ �lhSY�BQd����7W�6�B�Ko�l~���'�[�sY����n{��C�{��������6"��_{,�Hֶ���6j�v���x���q�"G�:�k`4����P�f��h
�3ߴ(��yY�(�!M�I�YأY�Ԛ2OExF=���m�Gu5�L���:_w���[����{7�¾S/�]K�����]f�`���m�c��	̹#~�����!y�e��S=����d���͜A&<ɯ��Z,H�Ⱦv�:_���[�0㮍1�~�<f?(�$f����xR�,{
?Rd�XD�SU)�������Pr���r}���V[7���,�Bpx�e�ϣfӞ�],�Tq�<6y_*��$�@����#hB!+mB��$�gؾ�" f���̌�3BAK����9��'m�4�̳b�*dV:���+�bt�'�z��.��qI�m3�1n6A�˟灒&�{V�r���z���VLyb�y]�)�|�ä��a�ɘ8br�ϱ��ւ~k�m��4�v9(���n�
S`L,�Y�~	������S� W"_�F�������0�h/�bϰ<c��wi ;>7������#�橿
'*8����&��{3쵸p��51h/��Ă;k	�c�U�c 	r"ի�&��W�+X�ZH; Q�����a�'�0��(��L��C�G�T�X&��q^ĳgq�<��k��xFq3G��V�z��-�0v�H���; y�$TY����/iTS-�d{�`�{���(��9k�[���L7ny��N!g��2���-����{|��5�oDMF�=��J�����8��K�҄!3�ܵ�k"t/�^7j ��p��"�G6�I�·n"}n[�f K�aD���C
�W���0Z�J��-�!<h�����;�l�h�Am����J?��o7�Eu�g��+�'�%-'7��U���c�� 	(�'d�H�齎�(�V�4�����u�Vխ�o��b⨭U/�j��C�~��� �PpF��'��o�d+2?�YX�X�QP�	'W���>�<��o�����^J����Dco>�.VR/�mz�i��s����ءϖM/-O=|H*�N'/���x�;�Wư�T'~�)5" [��9�'�DY��u��s��c�#W�~��]3Ʋ��� {q�A��	p<�)�� _jQw#�I�L
G2߽g�#�W¥/��	n�LJ	0,�p�-߮�;�y�����ٞ%�,w�#�ho[�����侄�(�^޳㉠�j(�13.�_F�����"�S�rObP�O�T~�Ͼ/�S~���N_���"��0��"g���)u8�݉
��V��ȵ�gF����$�NK�Ԝ8��Fq����ߵ��8\V{��{�6�	'� (��� 2u�l�}с�.��D�	uZ�'�J�q;��K�+�c�(޹���$
~�q���U���q�Ѥ�J&[��D�xM;�I�/=��'�O���f��� C�e�K ��<�^nz��������O�{ ��F�����:k����i�(,�i�ՔYԇu��S�,۪'-���}�5)m��>�'m5�Ԣ�d��
 ���k��6�G�K��m��!R�׋�.ɲ��Nhm�NyC[�pH�>�����̘���M;|DQ�",���Y����\��(R�7G&n���&���D�R�zb�?W�5=��-�ށ���0�r~�𬚻G�0�H�\���'�����"t�:3��j�i��v<T�ptK��3�ś&��TP\�y ���6�P����Ha��4�$>Y�d$�3LV2Ɲ&�,ﻱ(#����H�y����O� �%�[�T��<�a�y�|_be���S5
oё�V$t2�F_���U�P�x������mvN�v�vܓ����ˢ R��"�\%�t�f�kvxC'�_k=� `�!R,btQ6��������l������*��H�,5ٞWBs��$k����nJ�=��8q�*Q%���,���'/3���(���߳2a0��_�t����p��ME+���AYP���0���[܀D�Åo�{����$9��!�(k����;F�~���0�����im^[2��iv� \�X�,?���W�$�߇�ٓa�\�9�3+%�}<ulQ8��8;ZX�j��7q��n��^�:��Ì����K[s�A'������L���05�(�b��KT	����h�G���gvmeJpߺ6M��[�T����\Nƌa�L�n��A����v��' ����0�r��'_�v��4�i	�1۠��aB�y��s�����r����jz�u�:���C���t�s(W���)Jz��D��y�ݓ�;<�"s-q�k��NKt+��ޜB.`qW� ~���S͒�%K V����P_xg����,�ST�Sؤ��L	&��ˇ��mfJ*�g!$a����
&Q���r����H@�Þ?D8�C�/��Ad�Se�)%����8P_~g�d41ނ�ܓoyC�_E$E�k��� E���;@���iIs�����|��o�Ԑ����w�Kn\��c`QD��K�~/�.��=�3�c��j���p�Y#���0�[+��=3��4`�����aFiz`��'B�l���c-Lt۰I�zY�������ռo�M3��k-���c���0A�|[�K�Į�|�YX�1���)���� �p�&n�&JA���B���a�,��ic�������Qܭ�"}�<�+��� m҆�EҘ`ы�9���՝���H/̜��b���3��9^�ӊ��x ��iǒl�~O��S4��ӳ�yñ%�%!1�	�@c�19��[�����uB?�T5D�C@��,2��$���O:Xs� (��7���>��o`�˳�/$��;XF6��$��P@����]
nqyVp�bg-����
�(��K��Y�ex��� H=��F!������0�w�ꎻ�݇?�ȵ���d��6�aB���뎴���|�sOf'�	ύ|�?��aW(F'NCc�һ���}d����8��F�#��S���$0�墉WR�Z�SaX1�[�[�r�&��3,$�	�yyS��2V���uW�KnЄ�dýe<AN�fz�w�O�:��!���:�����"���T�,�D�ע~	�i2hD��/������&�PGo�'@�N�^D��}:6�+T�4||����O< �Ls�LH郪��+��8��Q3�v&}�����.�d����Ѿ��j�FL�TS����9�{����r�V���O�WH��?a���I�=(��qY ����Om�-��7z������@c�6�-
16�L�jW����7�{�ѫE��a��8ֲ��U�7�@D<JP�:��|JUF�~I=?���z��(w���ݾS���S���5����=�v6A�_�*��½<��Sm
�#����m�43�%�9���tFZ���t��	|��2����؈���}n1�C�!��f�ީwx��D�$����=�@h`q��%N6kQ
��S[���U�f��-z�$Q���a)�V�\|p�A�L���b�R	Ȃ�~���ē�7�K�g3�������</�{	�y��d�%8���<��\�o�G���&܆��L�f�Ǡ�ad��� �I�wG��p�n�4T��K+i0���-������,)?E��;��VE�(�EK�E�g=�K�� ���$��%���c�¤���m1�K#�D
j
�?�A+�	��bڋ��p�G���9�1�1\�Ӎs�2���ym�M�L��Ҩ/�DLB�~�G=�P/9��՗4�(���	mfp����5 �2[���C�#�6�]|fi���Z��z��߶b��25�<���Ln ��H���9�NrW�la�aU�P�wlg7m�/���_�cV]��$�\��<y��	��2V- &{?K]�RAN�{��-`O����	D`�Ӣ��X�^i�`SsC}�dRQ�|�y�=����I��=�]�/��	��|z3��ÚY`mYN�2�	��$m��ס" ��l@�%�$�I<8M`1��cCm�>ȝ⟂P��!l*��mo�G|���T�B�R����׈SI_K�2H���)�C�+F��)�/IȔ��>���6�b@Ix�ʕ�^j�B�%�xH�PE�==~�����c>(�aI/dsA����647�RW���y�����A7&��R�w�
D�ķ�-����{����Վ��v�u�-{�*~e�.�Pc5��o���uuẽ����I�L�o���d��p� T��f]��&��ϟyp�v�N��)�d�U�,�1�[����م��'C;HV�V�s��Q�;������ٌ]�sϔ){��f]��Q{�sXIÍ�Y�`�!��[�)��.��Y\A�լ�wP������p��{k�:��شppeL���AgYtsg:�[$M��״u�d�C��7��3�rMMgn����d�~��2����)N���c�wy�E	:��	^:�x�r��X���R#+o�k�鸨sPPT�Y��B�i��ގ�)?|]�hA��Y���� {��̎q��Ҧi����qRC�'����`|�1�S~�Y�+3�e�#y a�ox8v>�T���A��r:x֊{H.H��I���cA3��&r�j4S,����p�����bHb���̸�����w�]�"!��
	3��W5���p�-�Jb�cKz�4�Mi`���J܌�h2�(�F=)ޚ�RV�c!�)4P/�	V_鄨d_�&Q5��|�?ui�y|�x���]��O)�R�+o�����a�IU��S݋%	D�K9��TW�?�؊��|�V�[]���� H{���zg׀Hk�D�,�>�!�Y������B&��F8��RT(f*'4�Ś(�����I�X��uD���v֙wD��Yދ�_+�F��q��u��仑@��摑֮��V&=X��[/&�6E\�?,<�z�:�s�z>�ҿ��U����߬�v
&o߇�U�0�8�ZF������:v{c�\�-(O�-#KL�Ϛ�ki��(V����7�fQ�������(߽��ʧ[������>=6�a.�B5ҝ�m�����@�M��`)ٮ�|��f��1��C���^b��`qΔ��t��T���kl�4!�s�Iѳ^e���>Wc�N�V|�W�Q?�D��]Ӛ)wt&�|+i�����C��"�y����p�4Ec.�r�;4��P��璼a���!u�WL�=�/�B�x!}�6T�Z�;�&קnfb?�u:�����g�Y3N�^�c��y#�L�Jr���<�~䄿 �B�܎�3NF�i����L���+�|I�\s#�f7b1K�ֿ����)W��/C� �^)1sm2�o�e^+pm��v�t�X�V�4�1���y���	P3�����/���<�,�
��7�j]@f�ǻ�, [t9qҀ˂��������w����@C ��
 ��hҥJ��gW4|���Q}2p��y���K���B��AnJ��%δ<�l6n-}��+���y��ک�lk�����TeK�Ώ=I�����Y�
y����
�.p׾��FA-5��K}"�T�A�"�= =��p���l{���37���F��oƠ�z���t9VY�r����=;�n7����B�r�l����S}�[���/D�Q��d��pe�V2�F}�vt�Q����V��ЄGȽ�*��W�/�,�����?�#6�S���(�7��X��7���] ���>M��˔���<�Z$U�� ;xݓ���pr���Y�TH�S^�*W���D����q]���9�Q���NM�ňZ�_�/Xu@��^��  �h�b�J(6�BR﶑NX���O�Ns �� 
�Ӆ����-]���J�]��HV����"�K.bHa��Ն�q��i����y�!G�A%�82�Fh�T)(�=mN��۽���j����>}Ru@��gr����rh��_
T�E�&xA3�ꗈ�h��n�<8�m���YUfݡ�,��HaOa̙�Tͯ"*]uE@��� �DD��y����}"Q��)ZM:�_ �ö�ޮ ��ks�sTO�~���հ��� ����O��=*�F��.�V�G4�U�\~�O-�j��]3�q9]���9x E�nS�!ƹ%=�VΚr���|�ou�g1�~f�Ĭ��2������$���ȯ �D���/{(��G<�%^�* ��v�#_��Y��8F�@'H���+��w3�|Plk�>����M��sY?E��rN���U��=8e�	q
d,����_e�~�t�Z�G�=1�5�+y�۬�Ӣ/_] �)�����~�����\"���>��a #9��F�V�^������Z9<� 
�F����	�fn]��\��Q�,�u�#��Fa	<l[Yf#Y;���nvv��O�C5B᪚���LJ}�/}�#��:�)�#�~R��g�9'�uh��ar�αpew���8�N_�夃����@y?N^��t�O�93r|�uq���D�������T
B�� (+˸�n┭�����t�4y��
�KV��r���Sġ"�K8z1oJ�	2X%-��[o(}e3[�Ӷ�,��ܵޫ�~�=p���
� C]Nb��?�&O���kJ�wxz����~ٶ��`�������% dW�:�A-�Y�Ő��v.E�!M$��{2-�Ec�M������1�A��?���
�J4��NB�e�g+A��,l�]^�Zd:�o&M�ZW�A�Һ�\f/'b�ofՁ����w;���&�6�Uǹ^&H�� �L����=��&7��9�^cך�`m����N�=]��"�E�`mF'#���]U�Q�/��2Gu�<5�W|m��g$�#ҩMu�x!My�mc��|��"lwŚ�z c3�$��.��CV�"Öiӹt$�ϒQ&�L.`x�����/���^7�_�[�٫Y�����\���I��a�����-�1�ax����"_� �_|DvYH��/���Wǥz�u�y��:v��_Bٴ��W޽��C����ӡׄ|DD�Zb�UߒOV,��/�Y��d��Ze���\g�)�6�3�O֤iѐ����nر��,�ǒz����]~=�IX[�/tΒ�!d"�)�ͭQ塎Y��N{�l�QVH(C�S�ز>ZY�t��hկ��y�Z-=��!8�#_O�?/O��n�1V(zFH/c�|���<�?�B#��:�O��cQ�Q���AH��ꮤ��𠭞���5&^$�b'Aj󚵊�	����ߩ7s�b�ݪ����5��fP8��N�42NX]��J,�3���c'q1�@�C$ ��T@���]��L�C"�k���I����=�~_�=��v)�F�ǌ2����h�;?�"�\;e�r*��&�OA�Q]����X�dF
Ǭ7B�%�&N������)�d��A�%���]<����P�S��)�*��L̻bF�3ܹI�+rt��3����ցe�.�߸;?I;^�98���-O[�e��/7ú&�l�E�GK�1���F#�P����,���^F�OS�ŧ�×2�N'�}����tYc�N�(l�d��,�NN��\�M�
{*yd� L(�j��΋�BU�%.<"
��J�#c��Y��%���l��&"� �Q3^OO{��B�B�>�߱'G�:me�m+5!���`J�-/T� �,�]�A@qOp�Xmd���h�fSNHN}/C��B"��*��(�������x�>�ʂ@4'���ǘ�hP(عe�\�P�@nAu?N
�q�ku��nC3l�� #��<cp�����Q7s1����Cn�˔^�:|x���~����^�['7C���C,'�<Y�a+�Ǹa�9Y��؊}"�lsؙ��P�c�f���?�UV�P�����ǭ���GXm�2��Y#*����[�h�f�Yf�.WAú���Pg��:b'�D�IFk<�Օ>�{"��R���]>���0ǄAc>�t7�����i�e�;D�/�A]7����=��j=�^S��p`?����W�(o��?�n.��?�H���3���__F���w;��8��Sr���� 4i�i#�_�o2e�m�~�b��~ܰ�S���')�Ώ�7�n)�v��ț�%R���nkpxWt��LrD�8�jA)
����G��<XCq}	�3eGu��F� ��*z}wW��f��X{���ٰ�]�+�F�P����z^�r���	ۆ���R�V����'��g �J.���N��	��*���$ �����	�ĬŘ����ԿetkX+w���{`���rL�� ��z�O���O{[�R�x��ǍLr����sT�{3]���vF��	��0|�so��g19ם6�i�y�����@il���2�/�	�\�-;����g����n�͊`�W��9C���ֲ�0hA�K���'. m>ր�ێ�E�q�xB�csq��Ŷ��(���g^�׶B�\Lʤ��z��2���\򽼈����741GY��>� ��?Q)�����l�;�S�Z���}�Ϋ9��W�9^,ҵ�Ӹ<��-�۹����������a�=�)���:�!}�%^��}��!qA�d��:T~]���0yW'�=R��P��H����*!+�r1��j ���r[�D�u�K���V��Ig��ˬn_��Q����D�j�؎^�i�u���q��D�ȕ'a!à��nq�F���y��Qr^�\���Rpo��^��dι��݋I�?5��R:�|Ѹ.� ���_�����Qȉ��ϩ��!�5�'�!��g�.�����B�W5Z����@M=u�����L�#��9��?�7T�ҏȔ�
 �� ��l�ʠ��x�}��5����ACz�%���ݽ�l@o�Vfo�`��HC��4��%7������ |GP 릌3\��e	;��ɨ�LM;<k=P��Xo��Ts��rp�	�o�n��n�yz�T��-�w Q��L��wG�to������z<�cA�]rL�F�3kӵ�r�
e?��A���أ��L	�^���7rJ̇�Z�+�o�g�����Tz,���Pj�"81Rn\ _�q�/��Xl�Sco����Ԕ�����= ����!S0�
��`������M�$M&>�/8F3����v@�j$��<4���dy��"�:�}қ�6qʁ��ʔ8,C^�'�u���q�v~̮��S��O�h��5ܛı�V�+��Ծ�?R�W+;��m������ʰ8��ז'���A��
 �<��<�_�W����P�|�'�ߞ��G�����يi�:-�TG^¬��^l>�^BŨO|��V��w�h�=�U:�{_	�яQe��P_�#\�$p�"��\�Ȓݐ2;GKRM�,��b;j�tp&;g/�l,�$�Dxi=�
L�y]m8I�t���l
T�6*F�O4b{̰*\^�͇'�n�~��{��5
Ɩ���#y������Z��ƍ����f�Z���Kj��3}"���{���k!B��Ɥ+$&�������*��u$ґb�$
���ͯ��K�":Q��E��wHuwS{�$9���F"���n���
���\���D�ւ��	���i���q�=�3�9�k�����x'{V]��g��a;�bAB�gB�(ZXw�t U4��a�x���!��0Q�X���dǘ�lF��mD�O��/%�K���� 7�t�[�KQ��n �)?D/+\��v�P�����:�4���]��o-���t�$��*X���8�}�|��;a򄮮�2��=¤�z{�Sܰ0B0��&�xV[k��ѣ��pp�z�X�|>�V߇dӅ����g"���g�}HЉ�s��XJVn��Ңs�E�V���^Iuc�|7���� VF�֎�
M��rk�_(�����7lH�0�W`�Y\F�҂v�p�֖�ǥ3���L�$�)�=�ѣ�TĮ��.^�%H�Kc���UO�?K^��]'k�],66d���ƶ���1�0!�%P���3�(�G���U$��'�
�<1����,��"��F�r~��T��!̩����@�^Q��Wa	s��Y)d��j��s�Z^�{��oo���b����~=Z@8������j���@�b�Gq�6kY��OC?|�f�3����y�.��	�!\����};i����_J��{��x5;�����r�Nb�hl%��g*w��L��~�2�k�T�&���»���nT^�(�p�?wm�ue��r*R1�u̴F1������c�س*�c2��N�%;zj"@��٫��CVȖ�u���G_R�W¡X2+�R�Dqk�ؚ$���ov�?���W�\�䡃CjD�%`	��D�B���Ϗ����+�t1�Fr�7�*+6��!%1"u�؆:WXd���`</��;�i	 �.�	`�b��Nb�p���j�k��-��4��.{A4�&E���2 �$��R�!a/��*+�<Hl�������|�n�ӳei~�?�$��~Y`lfAлF��dP�!X�i���=�����p�>Z��,�Y9��?������,��ҹZϕ!�U�撔5a�Ȧ8
U#�����#��!d�R��$_��E��O���
�SLh�MH#�a��\+W��(Kc�D��;��`�xD�"1b �aB�L����I��o��~ʼ61��;�C;�#��sa�+�H2�c=^�3Um5ڬ�����,kJ���G�BS��5S%�J�;Umg��O��R��S�(?���� �i�P�g���"�;n���N�(1ZP{�}��f�6��%Xz�9�CwP�u1``'$q	���F� .�䊯C�B`��\\��a�W�x�vj�;�O��?�{�X��:X-��yɍl��e�K�l�@vq��������R���7����1Wؙ��cl��!�(g���t�;�;ܑ�B��4:�Og��&N�x~��\ށx�Nx_�C�ƧB�v���ч���ïQU)P��>Qy�(bQU�-g4������3$@?�\e��k`+����e��F���:�}�Se��nB�)^�t[��������q��5�������~W:=�[Li�+�P܍_x���>�� �͗~�a���aY�����m)L�<�!D�L&�B���R���*iZ����s}��8I"2�5�V�6�"����e=�'J�R}*Yi8�Ѳ�R�����L�!wd�M6vW^v2ʹ�7��L;�6�~��*ͲN!�?.�b $?�]�o��=��P11TR�ca�w�S?��q��'Y��ѳ��ZsH�Vq�35��N���oѨ�@x�x�R����fp1��D�n�}�.��	�\�����**?���¸N�E����7	G�I�vM�9�d�������� ��@�ʌ+O0)���������l�<�$�h:7�Q��:���<h?��[8��ӯY�VWm�{�c��"k�	V�(��N�k>���)�Ǐ��L�7�~�`�7��k�;м	bֹ>F�z<�q���X���?t��):���}����̥m�@:!ԫdd��E�=x44J���m��k�d���AfZ��9�֦�6�N3�#K��"�����c�{�x�ET&p�jjYv��jϢ�7��vp�(�X	}���^���X�6�|K��ϷY|�;*]����3Ŝ�O��A�~�+�hY�L�zm����I��2��!�oksc�4�:�Vq��A�g������h�z��V��\43�}{�R,M�1��(���O�*)'Ʋ"�� i��=V��z�fM`)|�~�G,=���'5	m_�N�@C�M莞+Pʿ��P�]�Ŵ%a�_o m�qP�S���<IA�xT���!�K)j�*̲��O�
S�тr��Ⱥ����(R������ޔ�B%K������QҨo�)i�������1���N� N��e�AeT�8?{����(a�N��p���Gv�ɹ�oU&A4LU��j�A��}P{w��^L�Dx[�G��i��֥=��Kl7��"׹��R�H�Y��MW�'�k�܈���6�,����Mu����l��ݧ��i�� ���8�\m�nm���������U ���_.҂���R0�k�WF���9ӆp4�o� &o�	�K��Mއ��Q�	Q/�MnJq�:��R�<��%�0�Nu��ou��)����:Z-="��0���֎ ��}�r�vw����?T0Co�D��
�oĮ[O�榟�E�05D|���%P�8#�a��T=�Ճ��� �{\6�
&_�{��/i��d���>�N�r0��,b��%Z֑�e��_����)�VJ��u�@�H�6c�o�l�2ilߖAr��J@�q���ؔ�:�5�N�S�xU.4r��\W�q��d�G޶��	��$RwA�Zb�O/v�fR5�ܿ�dZ��x�Д��F���*�NE�aB�>�R�XCq�����d�����I�Y$JpW�^�s�;Kp�n�XT�`�h�b���G�M٫
1�����kP�<x�K������Vm��1����S�ii�/���@�/|��@��.�0b9޳�ȸs�����9��v-��m�~<(�m0������ic�Ы����s�A���p�*�Ɋޙ�J�y��`8g�U�{���7�qY?n�p��A\�L'dD��S�_ �5�p�S}�˟�I�#+1���j�%�כ��?�h��0�׶�$��t�S(��e5g_���]��r1ۊ)0����N\�c�C�(��xKt)����ߺ5P���z���������h��ksћs�i9m�&�ʟf�|0�~�ЮO�n�T���2]]�&�de����2��J'8�g���3��֪}JT�l�������5�=���� 6_���灴XF?|9�\��]ryq�M%$4�3�,	g��QE� ��D�pj�l`��&���Ѧ5F(8tV�w`�ڵ���ʡ��5%�՟��=����)˂氡����fe�"��[�dV����K
N�\��-t��I�n�1s@�f"��x��}*�W�9!#<!�#ZE
2=�${�#hR���N���y�� ������gpn��{c��M�\�1�-+!�y���V��-G	�^�	�M�Ն��B"��/q���	�?�v�^R|����r�����
ѽ˜:��0��ӊ\�:H54}.q!��Di��- �L��I�CC���X�
���Q|���$��r�҄����V z��`�ټ�Ŷ����u��}�,+��ͬ.s{۷x�Hlߘ��]+���W'�	����[ZI3罙϶�����
��5�	���P�w��AlK�s&ibg�����>���s�����Xp�h�tU�y�Х���D:���$�e8��Nj�&�׃T��tY��x_K��F��R���Z�Lo��g�>��x<~0|A]�*��}� d���]d�y^R�'�5Hw2�~�U;.��\��C�^)荨ʮ�å�iG[̘�n�΂����X�1��#4�;~���p�t��آ|؁)����H�p�Z̔P)7[`��]q�f9;Y��(��C�'��;?�_���+8mhT�E���9���Q��ñ�ac>�]B��U�X=:$�I��$��z+����
[��!�˚΃B.\��2�v���@������)�\�o��%���i�<V]{Sp���=�Ŝ�eG+�j[�̏v�_i���#����(���֦�/k���Rt�霫R�����T�/��|uY�b��{��y{�hk��X�R7q��*�`�h\�@q
��QyI��������_&`:\�@>��FOW���3v�$�s���N��tC�ș���� ���4�$�ӄe�8j)��^���~����]���D���j9��h�%=�Q���nC����KB���t���sO���vB�Q��AP'K�b��0��y��*+��!��Gp¶�<���J~���_GA3<�v	�s~ONΕ`�T�;R;)k�Ĳ�T[�"_3�D۰F(�ܮz�:&h���࠱��tg�9ᮄ�4��������|q5p�|���H ��Wӿ�U�$T��&Bo˻�-�ӎt'2C$_��B
x�ݻY��V9��Uo ��e7�����mͫ��/�/�U�c�`e5^�`�W��N���Q��v� �ֹJW��~�=n���z��D����Y�R?��x{�;�:�yX�11�1��*��p}�2�%��E�.��������Yx֍�:ˤO�b�}C�BFR�o��'&q�2���!甏��0}���#Ja]�+VV�O�� Bq�v
"�ۚ�:3�Նd��a��:��U�K��E��ռ���L'��������y�W�0"5�Y/=���)5���� .�s�b�y�l]�h6fCNj	l��O����wz��)ԇ���.�q.��z�Mmh�@ޤAD�(G�i}���L<��r\/l�r�]S_�`�%� ޝ��$!�ĺ�b�l���n�Ʋ�0��_��+z�3/0~YZn�@��&Z.RyAi����B�e�u�V�Q��s�>7��ᡨ`M�� �ϳ.>g��i�����Q�PB���y�8#��0JX��}� ���?YL����
{*M�ԡS���ƻ߷d���b��S�.A'�*��zY.��\�۪ϓR��f`g��g;���!2�C3	=�1k���u�RN2>��d�G��.��L:�ηHQ��>�/������9xFx��~��)���A~^��[�� 	%��X�8�;���$�J�Ek���H����u'�
�tP��(/ĻÃ��%�2չ�%d8�-(�4_��ºM#��ǟh4��&��O$����z������Ѡ��jNs�C4�#�$2b���3�'Ӈ�=����'��7�G��wlĊ=N��$�?�Kk�M&�?���y�,of�"Щ)B�csY]�X\T&z�~�ފ[Ʃ�Ђ������X��nZT�}��e��m�ꯩ��/
U�h�s5�9S�ԃ�Y�9"�UCg(��8�rP��e�<Ep�ɽY�}��mα�mec�� ������NKA%���]kRl����>�����QW�rH����uڕ�`(5ݷ�SY��&'c$ߎ�Q�e胉�p �o���w.�"~'/�yշn����ž:�c"_�^�y�Y�������оGIȚ�-[Y=o��6�.!�Y��0C�'ev����A��b�Cn�3�Oz ��V�棝4XM�C<W?'Q_� ��,[r�KK?%?K�`n<��:����`!?�$,W� YB������QiY#�8��cybp�@�8����q4^~W�ߎ=	]E o񊨿 �9��>4ol6� d���$ͯf��;r	����L�&�mTc =Zun�)����nF̄R~�wL�]�4�Ѳ�˃\j�Щ�t�p�'4\<AE���ϧ�뇟k��$���7�����O��b��j�%9�jz��J� d�
��m�&��r��87�<� hj)�VE\� �wA�ro�t��_�����Y�=�*��勮<��@�*�'4�8O��oƗ�K�ynB,I?s`*Om'V�;��y���t�p�i�U��Q������?�-t���XR��õM�V����b7�NO�GlX�ݤ��4����#7����H4��Ĕ����#�vPϧWRQ��	3Tv������\#f"�2T�p��A�xz#��.��X9R1���~o����˚�B��7�sH`������\٘�����u��vH��X�X�ݽ���fP�k,p,�KWjD��|װx�I��߁/�_�����*6��c0�*�������7�[�l��s4`��(I@}����_�;��������������\T��j��=s�	��G�\��J~(ޥ���ga��4�v��}(d�N�w����h�Kvn�/ͻ�U�"�낟b��[(�dO���%Ӿ��$ �=0�ޚtǯ��:Rcy|I�����N�u?�̱�B0��v�%ҭ���P�Q�Y�9W�d�ӉHd��(�6?ymW�c:*��[�7�S�퍕Bi����wL50-z�9D�T�z��AIw���얶����?�`��p	�� }�ZuǺ�j߼C�z�R���*�br����~�Z�7
V�nL��/�|���ȃ��Q跁�-�I�&���V�t�����WT#�F�����S-���Ɓ�.�_��ъ��������8����(F��7�SK+�]�Lj+��`+c�@���Ҩ���Oq�l��y:l�h��v �5��� l����ַ�C�������G.��m�ۋF������~��gPӯj-�r[ſ��j�(�V����Mڭ����0��3���J��9�����+k'�SI��w�f���1&��¥U_�N^
��*r�	�k�-Dֳ�x�n����F��[��t�	��6�$U��|
�`���ǥ#��#-�׶G'�+�����(Ƽ�k�v���� ������Ak�YQ��R���U���׋��� [�*h�J(Z��jA�֬vx��7����>�Ҫ�~���v4�J&Fm��Z���-�K��J?�VLM5��3�5�e�b܊Ur�sx/	3+�LՋ&	�F��Ek�Um��U)mQ[���,���u6I;մ���c�DF�$�;���Sz`C��?���JZX�9Μ����)')�g��z�M�Kh=n&�U�/�5}{尩1���gxI�Ǧ�:e}�t��ڴ��ߵǻ��
�2�r-���q�}���H,f8k¬z�2x�Y��IM'��^Me��.��,1����S�eJ��!���^.���7i/�(1sl�N���ṣVw�������iد[W�������0s��Mc�zMB�T�:EE��Y}�Ҁ*ҎJ��pvڍ�u4����D�#���g��|��!)�MH{�ú��WB��\ߢɳƢiD�G��(Eԡa�}�K�A�+a���V�sś���j\oĈ�����I�=i�0���݅�����Ґ�{3���е?�)O6��˧�E����9-��}���b�\�t�`_4�?�%������"�x)K�8kH$(_�0�	ɒ
B�����Z����Ml!��IۺZ�,�ڟ�c�M�����{��ӲL��fȱ�PXM`��R��$PR�����ɋ�)�@~��>��hs���z�>C]�[؇�P
hB�g��C]Z��kK�amSx.�4��NצNEk�R�~ط�_�c���F�o���4`+)ʭe�-u�*~��+�f/]Cn����X���@�Y��sDd�0���m��VC���`&+��\��0�=_}��?3$�͞���������.�#ڌN�'�Uy�K܋������+��>����d%���7
��Q�!�s=����g�@�y����/����^D|��Zf�M��:=UT��^0��s�˶��f'XU�܃�I���c���r�v_t�w��|�����BP{l�C�8c@r��bkW�/�n��;?J��G]I�듀�#[�1:{6��Ie��ɝ��d�0QB�T�/'�g�W��P8��k�i@�T*��`�1ٍ0�Dl��<θxʑ!��|��t1������������J�.g��y�Ғ�$�ĔH�����B4�<�+O��ۈ�V�[;]�%fbnZ�yfu��o�u�0&O�jw`��V�T�ł��Kά������!k\�,�h��f[5�%��=��9v��	̭,�{�? ��NW��;�ph�R���|��F�����>H"�գm9(F��̵&b҄�^]v�Ěd��ը��Y�s]��/|F����} ~������_hʚt��ט�ئ׈5'�B9"W��v��T�G�'^~s7CmG|�GȰ��u8O+H�?�b��b~3����}Aw#�yը��W�.�1Q�S��V���&���yw��aUjiv
�3��)����Iiʑ[n���fEԜ&��3�A �7}����7"{��ʣN��y`6ۦ:7�Fc��|�Z��]�Ġ|�n�7a�����^0?s�0N�@�v}>/ɐ�M�IO�&����ҽ��}\�|�[;�笠�r#4P� �$���b�}��1�zi������Y��6���[:V� �40�1��R��Q6W�N,8۱_�[5}X�#00���I (�R����䱹��uF9}Z����~ذ�Y����k��o�*n
���N/��s�W7�\Qg���GR�!�	Ywb�]�s�wĺ@y�|�Q?c���f	��d����NIS��<G��Iz�k����?��>����rǛn�?N*{W���|��w��g���)� <�V��6
(x�[������U��o�3��flv���p���K�'�C�ݕ�6CB�����"�@���+JvgE�*ũ�R{pE�4�ࡉ�$4;��Ƹz���l��[�R����7�_&��	��W�m��F{�x�o��r�(@���C��A(V��ɺ��`Pj�p�x��{Ļ� ����j�:�U�>�ܟ��;$�t$�Z;2س�Y���H�`�x�+�R[�n�X��u� ufyX
�e<P3I �A���S�8'�K*�J=���{	��եm�x�y&`��!:,�zEcU�^�q:�M��P1��`eVvb��w5_����r
AU�*t#H��N��篁]���־�7���EG��y֋uX���©���Ns����Q�ූ��YZ���5�B�{p�J���FaQY9B;t�, �6'����"�s!��(X�GU8�S��Wf§��_����O׀�4%u0��[T�R�Pf!��/$'�P�e/[&�7eHƏ=W(
MȪf�-�~Bk����A^�o�g�FA=�'��2b�Э�S�u����T�y��	�x�5Z��9�sE<��З�F��!A�t>*.@�ȷ����HB
��3���6�r\��ֿt���Еb�L�A=H�	�^������H�gC05��W}b���M\}���b	hn��<e,	�4����&Ư�i	�7%'|�{e(��$��(�|Yw=J2���x6��~;ӆ�	�M�g�jj�VD�X����NV�8��t*y�@R2�NW|7���n�q����E(�J�4�bW֝p�$|�H���a���>=����)HF�؞a�1��Dn������G~��6�o�e~���b �XzCȶ��wɯ����n�t���M���=�u>����)�d<�4.(�(�2�d�*��ԅW��^;b҇���`lX��B�+:�>I�U�.S�p(�Lj�f�U��[ސ�%�9�w�R���Wau�,g�2��/�)������X3K��S��qU�;�˼Կ�ܐ7GO5 >�As��ɨ�m�W��w��ɿ��FE*�6����!��j5%`�9�Uq`�Isr���P�&�ț�����~B`��@�=�����sIw����CG�� w" �W��aze'X�y�
���?32����Q�w,�E`���2���
�3k3��R ��Y�|����Y��,垃�C�(���cg����fީ�6|��&��"m��j3vu� ��D�ĀՐ�^��!�^���p�6�o�ʫ���|ƥg0x��sv&r�.ο���u��&͇�e���6wZd�
�`;�Zo�P�&�����N�P\`��`�`�=������b|����'�K?!.W���w`KL<�Lx�Ξ~p��3�JS�`��7��FfЙaP2O�xN�8�Qav���2.���*U̧�?���̇б�Y�5mi&�c����G�:d^�_��*�F�s��� ^@�u�J����D@�\}�{�\�4�,1�E�*�+�rF^}�'�i���5Ӳ�E��?���B�7 ��e��2*�@��K!��j|�
��-�4�@������[xP(}�:!3E��5e�4�'&-�!�J�M̘m�_}�#��i¥X[7%�H�"�Ǎv��P�l�;�k��M>�T�qD\�ǰWf��a����NG����"%��Y�����v��ɴh�;|��1�j�W��F]�����ɸ�j�a2��$P����~[�\O��9r�S�K��N�PI`�iZ��D���*sR�o IΡ��:d9�g���h_�f�� �����?h/U0���Ed����Q̧�;n�}��z�i����Q��NO�bLp���Ն���#��^�$�&D j�fwO���&HE��Nw^&Gj5ϩ�����EW�Х��\f�����u����>W���M߂���߃7[z�zr)��b�Oi�f��d�{aB��9
��۞DBR��5.�\��؈TcM�ї#�7��fA����%�6OIX�c�5��SW��H��7m�&����8s9㨂S������/ǁ#d�ʅ�����Z�@c��&!�{�l&x���sR�n:�\M{��(i�Ůp2�#���5q8�?�PC�b'��d�9���O�؁�C(�F0?��9���O�ԁ��Z��o-���� �E{U��]Z�l
��3ҴX�
)��*�mf�3�vP����Zn�>��r�H6H7x���m�|����j�P��C�h�z��J���es� �l�!Q���8tp��p[C��\�<����8M���ϧ2~�f��K�k~m���Ϲe	���}�_��tg�&�d%�8�y�#��A?[�K�١�4Ƙ�v�LY^r= /���~��-oc�?�5�ӥ@yO1��+�	�LHx����u�
:HE"�ˤ�Wh-���w8��MC���~p�����fg5e[Q>�ĴgБ	��W����@	���^����d����|GMɼ�����qwb6���0��5�b����D�Ĳ�#�O�����g�0������;����J�o;;K��y�ܬfX�ּ��"�W��֜��:eO����t�#\�0s ����������r �keW��+���L �S�U;���|�!R��ޢ��}M��Qk��G"�i��1Y�^!^��0Тwg|a�����Z�v�Tη�A�R�TWE��l��v��|���P�hG�qf
K�]�X���j��xl�|S�WE�RX4�c��B��;Mk��Í��PČ��3S����&�EJ��ׯ.I@"n�J����"y���u����)ON s	!-�-E���a�[��5!�|c�"�A3�;����1%�BI^��L�M�$E5�|N�w|�s~��Q
D�Q���2^��l�g0��M��0P9D���&���[�������!6�+� �_|ECV�'��e=�&��<6�1�����Y�1�\j}�lrǕ-�;�D�$�QX��-)5��T$5��{�� v@or�y��^*��D4ż�-��;����^k[�;�P��³/��Br�P\|��`�m"Y�{?Y�s"�?���G��^��+f��kwk�D��"����u�!���(�D'���$����R.(����+P�KC`Y����>��W�!*x������wٗ�JI�ۤq���H4YO��_�V���g����y3�|a(��7��`��0N�ī�.��C�}�������T���"�-�Q�m��t��#xnH}�WW4�����=%�	�=�6�ګ���G���}�{H�ꋣ�EP5����J!��ć*���}��\����{oG�cvBx�����5o������:�9�^!��w4�u@ ��]���c�`�; ����j��R��}I#�4ˇ��5�/vg�e
�4����[[��n��^ǯE��A⬝��� ������?� �w���ކ�/�J,e�C��;���	�,�O3�S�An�FKM.���);q�^W*&U�`t��L�Hfb��e�p6���>�_,y�5pvFYLZ�)�>�CCCa�[bɠ±��0bj]�;�=���ܪ������W�	��W#�*��aJu{.���q�'�����,��%�ƈ�v�۟{�>l�j*����)���ga��VBͫO���c�>5N�X(���!>��l�O#��	d��=�UU[uC�P�Vu��ѻ�����ֽ������'�`�h`���T"ANH��	V�(�b��z�O{�p&�Lx��	1L�{�����}�f��0k�=��w�|��_aAA��t�L\��B��_�#M(=rQ��J�X��w�D�kk, �t ��:��L���Pmn��UV�8��*��6���ӶO���}�4Y��GR4����N���3O��[�D�jyr+,�a���9\�RW�d�2Z�� k ֢�#�L�_!�r8̢%ZS!I^�O�5W�'�d�bQ��k S�h-�OB*�S�8�O�ϸaR�Vi��8� ����d�aBm���L��O�ث�##�	A���'͏Nx:�\�i��G+���Xΰ�$E��-�o;5CY�9�l���E������P��K��P��0���ލ`�:6$�#c�&�KD���04'��1(oD��9"HT�7w�n_�e���~QԮ�c�(�b��]t��g��p���vQy��Y��Vc�og������>����;�fC6(`�]�v��˴��%^��L]\.�&t����ԭ��\
o`Zx3	ce60\��%_m�ր�iAf�0ҟ�ۀ��μ[������I8z�D��� ��u�D�@i�.N���BIV���Z})Ϫ��<��iy���ru.��	F
U�h�gw���1�%���\b�%��sƸni��՝���K�hWM �#���'�'0
@f���ԫ�g�6�ч���XT��(�8��$��&���8�w���Rrj�C~��P�V�buªo�50�a��7eXP2{n=�k3�-6��z��H��L�M�#
⸁���uԋ����ذ��g�-����z�w���i��i �8#��{����W{Rk^Hm�d�Hx�����О7~��+.��$9J�vh0MF��m�
v�k�f��%;�uڃ�g���H\T�O�>ď�y��W$�S7�{}���b�oa)
�~��-�6��T/�Kw_�	#ZB��%���]%ν�b�h_���Vz��x>��u�A�n��d�n��`�e��{�8ל
�h�޶vB}fa�uJB�,�T�,�ӤT�s�2WE2������"��`���XZc9�<'�����kG�$0)`k	���4���"�kBlZ�͔OI'3[�é�sj�"2۫�n�O}ݰN\N���!~ M����	�n�_O۾���N��t��7-n���#~ �%$\����A�g�j�N]����϶�G![/�����v����F�%���S���{'�A���CKj�2�k�җ(�M��-�A��sw�n���}�kB*���X�pG����=�U��4Xφ6�ez�>dj��u|!��|�ß�Q\�)O��4wY8u������pl�������BE�~1�}�m0�k����'Õ���)�S���x@ni����'S�Cp���/G/��z|W^�oI5壵x��/��bo�2ഃ�k=��p�������jimy8��n�������<?��U���zfq��X�j$Ŭ$0v4GyG��{�	ȡK�Z�}ݒ*�ڏ�.��wq��Q2<@!� cD�̡P�)`�Q."s&��L��Q/,�h�س�݋�����q��	ΣoOJ��"}G��[�TFX��qoR�N��O}��Y^�Jo�M]����{�{\�}��4P�e��d:y�Y���|P5�_wǥ=�$d�q���Fm�K�=B�$���k�cߘ�e@����2�����AsB�L�������S�)�d��ч��Z�Fs\��\�Ô�3,�vX�����⾃FL�IE�����~�${�f/���܆�M�@�����	��us�w��N�$IWF�ˡ��ְ�y�Fz�։-2.��D���>�}��B~b �tj4P��Dն�6Z�&�-�l����鵎g�w���N��i��)�^�P"��4J�Z��a��B���1H�<�;<�=� �}�T���R���?W�x���@�����bE�q�^��%f[��^��x	��}j#ӎpr���M��k��Cc��&�SR���q��4�	�}��<C�8�.�yt$y5�ʒ8]���S��5�;{K����{�&�� ~�u����C�ЃO��:}���5���o;��z�5���m����!��UykZ����ě��Ea��bhV���(�U�{��� .�>�b��1�~���y���F5���x��G�y@�p�I�h�`�C��,�.��gK8�U�A`��z>��Q�}U�C��V�<��*�FlqE͉|Q�u�[��`�i���j-�M��R�Q։�m���.Z�5/GDQ�CV�I�ao���tL�ʳN�h��F}�zh��2���M�e�Xna�F�o�a�Y�����WƬ��Z@eQ�����Q�'���?4�IG>��>�>�2��;b��d�L��/��L�sv�9��7�y��ֈNL�Cӱ� 9]8[|}��%������e�p3S�K�K/m�s���3DT��<�R6j4g�|�}��*��Wk����e4)��i��8�i�u�]Je^����U��-Y��=�����֐a�6*d����p_���S%�)?@�Q|RW�SV%�<���ս�-�.#y�~f �b��ǜ�>ܽ �)�� �Y���;��-3����i����Y��p��e��g4�����	�t�U�n����FH�@��}F�����[$2��Hle�o�rJv	=$�*5�a�L`QR�S��p��m*��C�����o��䁷_(�+����g�1�:�r*��mo���2�e�U�+���&����g�B
}
�a��1K���G�k������q��L~�s<��v��=�m����а	E����UZ��C�<=K˽L_���V�u�.���JtJ��(_��꒮�+(�*��[��G��x����(�ļ��m�"O�5Y������	t_i�O��/�瀟Őo�Se�5~��u|�x?O�G��a���u�R�Xo	@s��Oi�������D�`+�vo΃\7s�h�G4$�H�}},�v�pN?��#�e>_%n%� ���
P�C�n%7�����[W�@:�BL��f�x	u`�1m2x�
گ� �ш�>ԃ�|�@2�9�J�|d�?*�]c"�N���LcqQ���P5&��s��ʣ}���l����}6��:�n��B�����RN	b.�#Ψf_y�3���؉�#��z��uP^�AU0��H�]��A���'D)T>7`����5<~])U���IT�_�4����F��nlҎ��ω(�%j�E��GBv�M�س>+9�i���jl|���f>�q�@+(��L��P�P�f�@1�F���V�k�vtW�ӪW�K<-�G���u5m�4j�@�4\�����-�߄̲���'+�!ݥ��UEw�����GV^��w���X[�̖?V���W�Iq�|6�E�:�Y�3��G3�C������V��i�&�����l�i�n���|D��3N)�F��g��>`��N�o�b���I���W"P6�>dm3N4M� �F�ׯ:�H,uҸ���8Q��CŹ�	�+YLG����-�Qh���ng,(����.�e%�s��Gq��S�n���iˀ���u���'L|}�._
|�8v}�{��uͬխ�l�7E���)z�=��8[km�b*cz
���^xI�'��"v����Tğ	_�^	�b��f�%O�EHA���䂫Y�JPعw��U��#?�l6�a1����~#S`rջ�ه2���[6�)�z���Em;%[�o�Ky_T�4����㩗�	;�l���lG�mC�I<���#P<[HV.Y�\�L����װ\�s	�@Ӟ��S0)��)Wm���I&*�ۏj�"�js��'�����ic�=�3�����π���`�"A��
�� �{A~ùM�-L�#6��l�Hd�]\��[enq:��<k�o3@I�kGS�I��S���UC��3�|���ٳE �h�3)r ����6ү�Roil��n �1����2���˽K�����r?ҙ%�F����B+�)[L�؝��(1J1~H�Cm�&��!���)\8vSS�{9��a�n��7Ȫ_�gԃ���h���k��+�k��x^JP���Չ��E2�%��3�����i�T5�mWM�9Dj8+�����:�ʩ��5VGZ����_����A�hl�!���#ŝB@1bY^'[�
�t� ���g�dq� z�2��z���J"���=�O����j\?��.�B~̀#i%"��3H==�BgR޺�UmIR�/�Q�Mg�F��f�!����g�[k���l�� �0���sK�g��^��+��x��� ����l��9���^X_�s��ïkvXQ߇�v�l�G�&J�vkD
(�����+-���s`�,� ��/��	���{j�X�{��l��.0X�43x�Z�O�+ N���#OLkƦd�lRG�$��Yc	m�Y���w��Vx��JQ�nK��9�%�#I�,�~V���t,e��9Тû�.�obd��uG=���f�����~�'�����]��(��wlU�z���H'��8��9R����1��?B�:e�/1�"��0`���/���4R�H�:~����~̓3Lu^�V�i�c�> ^C�A�����M�ӃD'�qqj栬F����&0����($%��Cg�8�,�Y�ȯt656�H d�F�:z1yle|F�[[�(��`�s���d����u]��1U`C�h�Kr����P}����W��:��wEѨ�C����mQ#��G�m�˷E��0��q#��KyfsS�Nb{��Б�ty�8_�+Č�Iً��k�B���h:`��f<w�Ww�/~]��C��$%f�xXp&B̲K4�����uo�H(��%s"���f+���T��q^���D�_��xHk�Q���u*^c�]��"���{�19���Y6U;n"{��SU��Q'@��A�9��u�G��tO����^���!/�Z�t�a�hȪS�v��ȼA�%�������9-��M)]!J�T��� ��N���h�!P�5X�>e�	�Mg��֮�6`a�x�@GMϘ�f�;�f�����ҽ�cv���n������jR!|��*yس��r�r>���cq�(�wo�������6�8�O�L��z7W�����6��	P�{Rc͵dE����p�=�n ��Nx{�u�١c��|���C�m����;!*r�?����T�B��`��wAt4'�t��:~��s���k��S��7��0�")��"�O�C� v�nI����yp����7ҵ�����g�
~Wi��j��D��rH+H��K��,+Y�h�%;�,�������8Ŭ��;6Um�6����'������$��˪�
�z�ru�)9E�m=$t(�W��"����>��� �����V6�{r���5�CtK��~��w2xD���#9�^<�(��]h�E�SL��=�W=��ҋ��7����>S��{��Um���CuN�x���vP5P�´�6L��X*�tz}�&�nU�鮑�J��ѫ�Oy4�H�ϙ���������Lܦ���ub�f��[n��H����2�����40�h��mU_��� [Q�-DI�T�u����@
���b6�V����`�Ѷ�M_#%}RKP=��.���m;;"�`�6�p�؄��HjR��gİ�����o_ŗR�|��3/���*�=��\��ET<#��9��!������NA����
��WꙪ�Eo���1�f�5u	�B�c@R-Tߚu���c
 ��Y�=4�'x��+la�b���$��?��Zs��Ѣ�<��#�ʣ˔��
���1��LG4����`�9;�K�DF�n��q�r�\�l��p����ߪ����n���9�o
K+N�<(�=b�CG��a�d�x��3LVyϨ���(�PEB��>�ً�n�E�oar~I������/�"���l�m�j��q���x�`{�g�V]-��}p��]'Tϐ8��E���&�v���:"�J��[sIn�����j\�kМc�` @�Y����b
���Y<���NI1Lcv���~eV�<ǂ�2�Ҟ*�������'�ǾÑ��ϩ�*2��OM�\󱦤��>�§��U~��6��'w�� }��ș��_�mW�~<�~g�US�E�]���vٯ�=�N�2F��/�ؑ#��X��;�Z����,��ۋH���x����h�O�\��B۠��@'��`��2����ӭ�<ZUn(�0����5ueTV��jm�F�Y ��j^�I��vN�	ש�۸|�9��=3H�C�笌�P�'���i��`Ď)`�����^[��%`���ry}�%È�Q�:����-�zy�q�e�"����L��x�`(���f,��>����&����,k=A��n���Z�:�Q���<��\BLE�?��ly�j_�ʹ'�xV}ǰv�~ ��R�:����9�k`�)
�=���ϭQ�ڮ,�m{J�3z�S�,�j�y]�2�5O���R�+e:N{z+����+���x���_��B���n�|�-�~~
�'�F�ym��$%�Q����r���(�4k�:K=�knN|H��lA���m��f������j7B���]�t���@vU��Vi#���ԀI�a���A�]���)S���[}�Yt�.�O�l��@���%N_I�l> 3��1��"��A��p�ۍ$.���S��`7��`L��o�$�N�[��ܡ��d�˨D���j���U����o�0`>�ߖ�l0��}7d���o��q����k��`�|1E�sqb�s���g���;7` �`L竇����-�Hه��?PK��,q�^r�%�1@�:>���\P�+mZ��p����Pn]f~�&j�����B�.�93-MxK�o�C����p��&�[��o��䳙���0AB���zUjRsZ8�"��#���	�?�h�
ʜ�cc���:�H�D����+���X3/O�$
la��Д^̹�z����_$)m������i���vieb������4i�L�d�Rv�&�������%��{��&�*Le� �x:-�Q�K�}��ڌ���o����.%[$�*�&�n�F��3Α��[�������c��1�r�|��7N&)��+u	��!'�~ܖ��w_�l]��ݘ���"l�g�^�,��Qw#�=#򈓺Ϝ���.��k-�Մ�:�]��sgʧ�'�6Hf�yj.;;�Q�F�c�"� rA��snj���*��_�+�q#d��d�A	�;� ��9u�����l`�_S�r�w��NZTU� �8�{CR����3��h��I>+����hT�ʻ5�o�\���2)�U^� B�yl�yƹ���0��t.fBCR��"#��?ă���sՐ/OMT���ih_@�����A�`8���-1~�.k*d���k�'ވ-�w{8���6Տ�V��x���>-��_5}�UT���TI{��J����7����`�˞�(��(�-���F`yi��hO��?�̓�4��u�����م����vv�b�"��,�bU�6��% U�	Fx����)�|�lEf��H��*Z�F�%�1�s���n�눘��1o�����Z��#S��&^B��:���k�3�'�z9� +/m�m���y����b\aQ�?���z7�+^�.rf^����1ob)ii ���A�f'�lo3���h��TH��LNy�6���Ґ��ך�C������-T��y��~��.R�I��[S�i���nSO3�-���SM.�=��p�&EƬ�ƅ=b�& �pFڗu���Yi�� ��y�%)՜����@��X{�UH�`�����_#aY��E�>K�nTW��ƾر6��v�\$�p��o;?	R�:��V�9��^XD�Q�5�j?���������d�5�ģ�ˆ�!��}��sI�7�.�7DKi!�K�IB7�)o�BO�wd�D��u����ۣ�U~?�z���(F���C=���o��9Mg�(���2�����Hp�[<�2��:�#q��?����J����������^@G�{v�I�� �f��I��6�!rk{�s�z��e�n�o�:�"��U�3(�슔�Dgq<
\`Л�����S�Q����������~@�\�O�)�f�q�(K�ᑦ�f�V[Xi_	�~-��9�WY�"��U`��b�9L�)��օ����B���9�z� �
GzH�8�(���J�W�w�nV�G��k�EY	�.�t�K�W4� z�_�Wj��e��?��>��<��Fw�Rd���u	���5|^xfP�L>M�w�f�>����
`7�8������P?�@�����ԅg�Ӡ���g���3U�S�.���#�-�!"�~�o\�[D��s��J����;�V������C��x�� 2J�,j�1����}��UA/�h�'|[�5�E��Ⲗ�����]u$|�)��YQ�F}^�^��&6V������s�U���b*lA+�a�IJ�h�� &M��=$x΄hXXo71�֮���9%��3����	h�����X�-8<<� ���W���+pk�w�d~�$�?vk��G@���~��Aj7�5}ܑ7��\��/ �~Ñؼ����u��o%Z�+x\�݊�X�.���Z?o����r#��ҋ.�}�a�u�\��G�L����W�rpu��$��8���)t4��{�����	�G��H'4�������߳�j��$x��?'6�/ЋTʐ���~f��(�"�s9���p^�5��������	{2�&)��~��`��o���Zc����4R��6��P1������޺�X�7�_�͟���
|�dFIe,bjz0S.�C3^ͫ�8;`ƍJU�˔�z��f;�T�ےR=[g�eua�B܄[�DN�[|.����I��z���g��W�N�U���hϪ���1@�(��w|��r�֯�+��h�x��S��3_y�m�z��엟r�̝>:M,h/9ŝ��֣���K�AL��JC��f�"������{s�OcL�LG`���ɳ�x�`�6ۚh�v���PE�{��B{�8jq����͸��n���I��x�ț%�z��G�2@�/�_ݹ�
}(�<p�sn�3��Y���x�;�N��r��_R���g�>����#�x� f�A�'!�:s�g�@sY2�M�Z��R�g3������=j�	��{�C���N4Oݖ#�7x�_�S^��ż`��Gn��i�c�w�rε.���)LΥ�e<��t�j1$�0t��U�O:�2	��R�e�^�\��(T�ܔ��{$!����ȁ�/���inLh��2���!I|�Ϗ$B��[�~w�q�C��ɐ�f��NU���.���"y����ᴳ��z���h���-�rFA�vM�v]�ᅸ�#�Y��qt����-�׉e��z�Ȣ�����I��E���>j��ڽ,���*�	����z��x����rQu_M�k~�Xs+j<���a�޽�U;h������P���tNm����E�m��C�^4W0��j4����Xϰ�l���Ю��i�vgS<{j�I�8���6ْ���9э�F��uƙʳ=�R�_�E[=3��}�۵�*Np#Im���vx����tkZ(�Ml�u���z\^TZ|߿:�M���Zᑞ�@�����D��E��>�%���C��Y�5%�d�k�C�=������HG�2���5S��Mp�q�vw���t@��r�e���$����5���^ �i�Tظ�_��s0K��z`�lR�O'�ò�NX�G��'H�m
9#Ը҇���Ї���-g��r��Z�w[aK���:]�j*�yX�*�Mk�Œ�����I����WT:[E}�!����-��<e��C^^�6�@����:kR�ښ�zqvA��?,�/�	D?:Z����Ej~��y㩡,�|���؎��_����4�1qE�Z��W��ÁNΊl?��W�/~��M܄����Z���$�\ {�VX�:l˕�urm��n�b��,AK$��p^d-U��� �p	���n�X}�C��}S>x�A%]���F������;�\��A��٫���Y5�l����=�Z��Fn~�t�j�*��+�
xg)�P�^e��1AAF���٪5��bI��'O�W�VpiKkJ�p����� �B�0��9�Ɲ���ω����Ӷz 6�yߴ��0�w�
{.j0���{miog�r�,a��č�
� ���L�|֞F�,�g�Nv3��Hŭmc�������4\�����4B�U}��1���a������FX������$��Y�Q���P*�6�F=���z�*|k�o~�0���Tq��u��&T2����$5lo�u��j�nl���@���]GM�0yf:
����Iy��_�P��s$��t"�/� �?���q�ws��^Rϑ�z	���4a}���I�rV/G]F�x�^�䞥)�&NDl����
��wp1�lSx��.��T�1��lT�.qg�Q"IVV�@�H:�w��s,������1o�h�@�A��GW���2>q�m�D�h.$i��n�[�(j @!�+��c��tF�c�V,d�j?s_�=���l+�	t�w�O���䷣E��zV���^�/��&��]��x�u�b����q�{�������[+��5:e(Ҵ�Ꮟ"3��f���'�6;��k�ա\���E`]�!�����IV,Г�%C����f�Ⱥ�����:������]��ֆ�TN�A�l(i+ݭ���{<��Ai�
p��j�����F8��z��Z����p4��Hn�+����!����J���ȳ��aC���ĝ���GQ���n����i�īaF����]d���dJ�9��e���q���8���P���Ó��>��Ԇ�sD��t�R�#yV���}�CQ!��B�ys�U@�e���wM����D_��
R"���>t����d�ס]���ΦVAL���\+�t$SPă16�5KT����Ո!E�3*N� �OΞJ��?����7W��O@�3�Jkâ"�
NV$Z���U�&�W����՞���m��yp��]+T:���b��C����J��%^ܽ#(�����������w422�Z��zC��ޏsy�-Cן2�ng5\[�w�l_�Gq�s맇E�y��L�&'K��2�و=��j>Cޛ��1Z*{�mK
e_}T�Iȡ���5�k}�J�oH�<�X�����K��77]���j�	�_��g����^2��}Ӄ@x#}����9�j�z�KT�q�Ĥ����g/f�qqS13���P�į��¯�F�(~�Bn:�B�G�m${;P�U0��t�8�)E�4�aῴ�4�q5�d��>���#1/���$���R�8e��.Ŝn�- j��dQ���j���$�M�x�W}I�i����I��2'mmm��!\��%�<�
rA@�j^׳4	���/"9�s���K F�~�gB5q�ҝ;3���{�_�"���3�CI%b't
���<o <�ql]6t��N���*�_�c�RQ��x<�VmY���&��*{WϢY"���L�-�!�fw�'s�L�gL�n3�l���BC�sA�����|�@n`�S��7�Z�BF+�R����j�j���AHMQn������S�e��S�vNH7��b��$�F"� R�����UL�Qu7�4���2k���x�˦��6ң?�Bri�w�^��<K��T&��,]����#�h�\��1�ciS���+֚�'}��'�}��*�8��w����@���H[����\WA �K�����ㄎ
3��=�ٳ�X�a�< ��^L�=1H��F�!e+�����N�B"��2��=�e�GB$q��K;����uA�H�Q�B��*����Ү��R|�߷����$s�٣n�јBJ��e6��x.�@�>�*ɪ����p�|��T��3!��fK��L��.�J�<�\��r���Od��L��N=
��(t�E�)u��Ŏ%����y�Y�Y�_Ŝ�G�u���9{�d�i� R^�z�Kd'���XA2溦^�ms9�*�js{�9&m�>��~}�XZ7��I����ąYʲ���M�5��� �^�����Į&
���\�����`U�$�)ܖ*���i��e��j�\���C���_~}��ppHS�1��:�I�o�%6�e�`�y��ѓ�� Tm1dx�EW�=;�{>���|:R�d��oP��;T^�<A3�Ʃ��6�U;`x��]���"��͵�JULx�H��{G����I�
ݔ����7>���j�x��Jp6�_H7.[��5@|�wuFB�[h�T<	F�Uu"���0�*a_;>wG��ܫ�y�4��|H�ǁ�π�9�z�O	��@M?���)����A>����"?�κ�$�0ǩHJq�Vj���H�|�7���:x�"!?.�+�Ӛj�|�o�@�^��7���2�<MȊ%��&�tQ�N�H��L#2P���3u��C����"��>�|�()R#�(׮*�yؤ��oWf�Neu{h�\C3�}�u��uˋJ�Ø?SC<JdS-���M鳌-qʢd
̲
���1§{a����|l|�̥@ՙ��}�=���Cʡ��&��i�״ .mP��ZgW�*[D��r/uuK��6��l���LZ%�C5Uc!&g��5{���"��>��
�=p�/
AKz�缁?����G����&\;{����fݜ�<k+ ���<�ǀ�d���������m���B���wА��``0j���÷0�m��cv\p��My.�P�J�G���nԎ�Ŧ�8��T�C�@)f��.K��~��8����m�P*��j��<�iW�g�c�u%u�f+�� ;g����`̬v�Y�
̴�tL�4���U����@���
y�d.��N��Cͩ�q?�~��3���v��ڥ�ܞ@ǈ3;�� �p2L��Ꜹp<^�.~�Ef�=�a��Q�9�s�	l'�/@]���/h��̈��MVy��9���i,��i�5��� Mz����z�-G�$��=�?�%���PJ����9�����q����L�^��=��	B����k����P1��eX�?>�07���},lI�y��w���@�Ɠj�oIQ���	G\�8�<���@�� ���7k��ܩ��il�;����fJA��tP�>�x�Kd����[�Q	�&I4s�#����s��x�ޢ9�fH�!5��R�!#f-/r��@nh@���hX�ʚ}��������(�����	�,����C�a�i��"P��n�SD���kɓY?`¢��eX��'Ȗ8ug��Z���ƣ?7A�%"��j�}���?ܬGaey7�ɺ���2�cbW;D��C�R%.N�*�����7�c�%��)�"��::�pq�؃�����Ra����D�Q���/?m�s��.A2���,�S+I�X7������}@S��fv���~�E�RC��~�����kה�̳����Hl���~�j���u MO`����Ӎ�Z���T�R<�\׹l��*���%��e>����*�Lp���)c��Q2ܭj'��SDMj[,?�?e�|i�[�Ks[2��x��	��`'� d�K�IN&�i��`�E0^�f����sfg(��
��FR���ѽW��z��rf�%�j]P��D蛁۸*P�f+|��k[�T,#�������o��sx ��h���G/��b����T�o�a�$�t�(�{�">r�iV`kW�p��	zp���Sb��[�`?8&�6�H�f�3�9�� ���\�"p���
�ȃ�k ���PYs'�x�����c��-{�����ف�u�[��\b�G#��V­��c ��=�q����y��@]���n�1/� �M^zs�i){�e%Ъ�6�Tx�W���O�����3"%��n@���y�f̓�������Oh��Kn9?�IIM�qw�Z���/�B�d�j*�H�;������,�!�k(� w"%~�#9R�����f���9��g�>��!�b����y�Z��גw� ���74�� �x��1��]X*�d��"���4��_� ��*����7]�����ݐS��3��P��m�Z`àRě�Ho�?v�O���cu� %�3�jC �P�� B �i�Ok�� ������;���8i��������䐂6��?q~ �s1��[���hZa�W��1����fP�r5�� -Ƚw�g�2?�����v~*ʟ2�9��z>m����^�h_��_�V���ۊ�cL����>,���p�LP�8�E�@��6�B�ߋm h��b�����"+ײ�N�����D�6.�n�¼VW�\�2���[�TZ�`�m��E�&��'������ބ&g#�2h���K�n���Ļ$)�t��*�r2D�/U�X�Th�S�<�'����M5��≉��L�e,�����m@8���MB�^�����;9�(��m
�9*�K�/+|�^��%ҔS�Ը�=ޝ������6�}�U�<�T�I�!�FXX.
���n��<����ߜc����*M)[#;�TX�$﫼$�^��g�� Ҵ<�'�ʲ��0�Xpj�3+7D��b���_@i�z���31����\�t����f��w臯_D٭ն���w�������ٶQl���A,g�$���B�q��vX'�H�Սa�R���,l�e��:{? /�	e��垕t�D�t~�ح��'��C|��ޑ�=$��Q����v�o8��F��B<�r>��ē��%���0eP�C�1��gq���܉��򕹘09g]{��;h*c|s\$��-�q�V�b�y�7��6L��;��3��*���p�&��7��Ԇ��ba&��EI�sd�34��_��ֵ%��j��&;��~l��	�'�äA:S��[�h*��{����/��
�xo0D6{o˄��<�R���i,��o$����'�EPYI���l	g�!�!����wi�i�#��va7�8w�i[�|>K�(�S��y$�"��:dk���D{��}v>�9�$�e����u9�2�%%�8x��������ţ�S��j8e��達\����٫��P��b�X�3?����<���S���>d��p���V.���@6�&��t��k��Z��>	_3>�*a��ۃ���]���=�aaδ�Ğxs�&P�<����>�ZS3̴�5�%x�[����n"��[7vm��y��[�:}C�ʮŌR�<8���KS�H"��52�㫾��_�B��&f!,r��c�*�=4X]&<m{���xQ���tr>I�]~
���cW�S����1p�^cr�G��*wE�α- �	�*Dr�.��u1�*�}aw�����A��.��ǋja]��C��gJiJ�[�Lb	F>��/
S���(a���8�eB�v������{�y"S�J� z���p�[]����p>îK���U����'F��8����¬��q2�L��L�7X4��@^��=&���A2��I\^�N��e=E��f��Ж=Z�2���@�|���Ę#��b|�v1��ڙ̂זIc2�i�����^(v5�z�O���7�v�x������j��E�0�9l���)��;��� D&ã߄gC��%���P�s��GYY��V�����Τr֪U����=�Q$'>gt4�_��)~WXZV �%z��8�������q�`޲��Y#A�2g���C��/��'ӄ�����=�R�8��x�Z!�7�v~�J)B���=���V��$F"3G{Ȣ���o��";��(�}1���`��kξ��%	Bkg��M�p@�lQ�x4�h�2��0Hh����ٵ++��K��Y����i��Z8ޤ��	����Q��,~���B�9bT�4$�
JO��503����3�� �>�%H�F�0�u�O>�d;��y�4�_��,�<Z�Y����·
I�/�x�$��Hj���M���YF�L�lAH�8�5��)I��`\�8�D�����"����o/��l�4_�"�c��|�|@Ш�9��t=���%�>&!ϑ&��7��^���E��1���6�N��Yb�fO�Q�$"���|<�}�p���X䖄w�+%�`Y�t�|kk��TU.�a��qX�#�tV�i��\9�@a˖��	�5�H����`��Wc����V&��{�w8̿0H�[3$r�3O�D�c����`ց�2tr�X�5e���d�+�������i���[<�랏����߉%](@9��f���,����v����8���t��fM"�E=��a��5P�RxL�i����]���=@�z�N��u��}K3b�?�/i�[Fya�/���U����,hp�	�(�����s�b[LE��s�����h�����o#�g�=HU�u3�+��������u� ��HP�zN־C����?�,����O_�p�?W�V�&C���H���J,i�I����^M�L)pG�����_p�3�5'�������c�2I��p�0a8���{r.-�l>�2�Fub#Pr��6s��s�?i��
?�dz�8Jt��"1�6�=�Q
���\�)��%�|��EIպ�5�4��h�6F�����Ў��$��j�D��'Z�a�?�`_��x�&)PS�ׯU@�k���������C-�ǵ�𦰇�$����E��{��]jK1��3�R�"xo��Q�Y�G�DR}|���Q��`/�B�P��#��J�ѳO��e�|���I�Uza ����y�j�yWz�4����<]5�(��5\��R�V|���NJ&�A�0�.�G��� ~ ��C1�����	^�L��લ�_s"RL@͓�|�+�����Kͷk.����7�����˱)6K&_��ײ}��p����2��Y(Փ���?�����V
!|I�4����1�y~kKa�?�.OF�>G��D;�y#�n:a�Z�yzf�p��a�sSZX���TΊ'=V�p`�e�x�1s?�.�}'��:��(�O�w�+� ��q˙�S]�i�D��Pb���.AO��R�o��ʱ��2��~�hg��Ȳ�}aM@q�ʰ.,D
�Z+��l�e�&�sI�B����LAp�Nuߴ���A��.~��#��x��Ri�����9��"����,�^��N�h�_�#�
�����N�4�/[���u�K	�A#�*U�C�0`	~嚱_*�p��/C�v��ɑ�Dz��䅓b��QvHHW���OǍ8�_KEؙ�oeE�E��'���	��̣�7���[�2)Q�\���vA"m����������N�����_S�j/y{���e���$B�)Ɣ����(��-^�30�����
�9Ӱ��u}쮷o����ϐ��Ν��r���{�i�u;�1=�[Ih�W4%Lgؚ��|�n,�\��N�imoiMU�u��N�z���F���j�Ն���AuN�� @�!��cK��i�X�L ��5��	�~�P8\|U����!�� ~�Nʒ�o\&J�m�]~��:b�ı�����m��쯆M"���9��)�����Ŭ��P����þ(����ǭH�ȓh���^{��R�d �cuM[�X��Hf����h��u�ߌ��(C����=�w���U󋑿<����W����e�&�`�Fd�2��a�MO�c����v.���Ǿb[�`����5��gN������ᛁY)<p�V_P84zb�/��7&�o	���r�t��Iw}}&��O�@��4Ȟ��c������Td4�U�,}��	��✠�h`|�{�G�)��"�������:w9���L��	~��'݃@���D`���f���4��N�勔a,��:4�
QM.��8Z�~�x=O����[��-�܊�\�(�o�v��'T,ZH]**
)I�P!�+�H�+^���d|p�?��� �Ͷ{��ŗI_���p?q�O��"Z�Ȍ$�W��$TOV���2U�K���l�@pZV��������zbE�����õ)u��K>��|SvX L��CcZ������={�[��P|
V(/T�'Y�'�N�|����=̞"C��8�:z^���ݮ#�?{~���ĉ����M�������?�A�&L����E�hź|��u@�[`�ة� cN������
�'�MK�}�|�c_��1?��)O��2��q�ew^������U������g�x]l�e���z�	m�x ��/R�VƄv_�T༠gEV	���$k�8*�CY�=e��7����¡�氚��%���=��1zDn��]!'V���򙀞�L�M{��
0�������E���(͛'#
�����].Аo�4vUy����OoEZ�dVb�Y�)�F�˜By���ԉ�t�N�.�c'N�2��D�O�)��7k�Z.�������;��+`n��l(��'�C���[�����6d��"}��=���A��X�[<CϭvV���KA.��i�w-�����R��;֮�s1��<CJX��Q�o��]c*��-`mt#�J�ik��	_�'��)pm�w{&��8Ҋ��&��?�`����G���_-�Mǆ�)�Pv~�ۂ��-�����xx@�r�.Qg�/y�Θ�?.9�?���\���������x�o����L9�����A�\����q���IQH��T&�g.\gu�C8�V�4OZJe���!�-`�c�d{Ȟ�2����I�wf�߉����H�"�DknD�Jk̷e�1�m(�Ŀ[o�{Q�<!w7ğUͱ�Q���Q�8O�������#��'�K}�>�kL۬y?킳Kw���è!{ �M�,�_�2�@g�����^�%W�:���ط���<:HȐ�\�����r��/"K��{��]w�W9eu� �8< O�(xZUv���x$�Ue[�:���l�-�����Kֵ�� Dc>�Ɉ�5�٧O��+x_�/��.(y����Z�KR}R�a�Z,�����lFYD���->@^Q/�1:�,�+B[	hO9�e\�w��{9;��z�͛_�)��$	�ڞ�f��&D�tDC;��D�.��%�$�Z,�M�(`���X;��q6���s���ۀ!����ڈ��zPU�R�H�=�߸j3l�)�2��ʋl���վ��m�@�� �2���5XO}Z}�j�����
6����*�\������*��~z���X�^��S�s���6;��[(Z�t_;2F��`L	@�S����|m��!��s�[B��޺Uv#����Q���*�Z�,n����*�8=X��t�p���+�e�Z3��?wc[�k� �������ʰ=��߀�9r&/W��{~��A#γ*��K�)X}��'���qxw����E Nìh��/+w�=�,���Z���^�N��U_�	�� �_)�+�/�Ⱦw�P�^ �*cil��ł��������BL�����W�c{5��5 3��0Kŝ�9�����!��<MO6���kZ����%a�1/�yi�9��%��w��n�9���7�|p�k��,o��[yiGIϘ'����'#Y��+�BK� ����Kڭ]��t�؋d紈C��rH���*�<A�-�����k��(�
줲�2[r�I�Li������Ȝy�q�Q{S	��ra�S'vë����p,7"o��tZ�X�tIx����(���\Fe�+�xZ�v�d,�>T�͎�d!����4:,���q�1�)Mg��c�g%(�6���&���p)��4��hA�	}v>�J��f���i�)����̵!R�#E$� 	��Y����ԂEtj��;�h
)>���	$���TF�ͼ�Ƿ�&"0���0�\\/��,٪}=��+,�-�Ņ�G: �ðU���gdv*�!�S��߃��?��ל̪����h�;,D����ɝ�Ģ��� �
��qV�|Y}/P])�� []�&�y��U��c�WB*N���pB�,$���(�yb�gUQ���)��	��E1G��E�\��

GG���9jr?V2
m>�K�)WM�z^�q^�e����I��ޤЅc�,w�,�6������pr?��ؽ�ڂj���������oE����D���"�.��N�Qixti��-$}�a�V�����C?B��gFL�Vr�ϯ�x��#`�5=W׎�g�\L*���zh����` H���mϤreU%�Qu����r�_J�X�=]���
�5P�:���z����C���ٗm=0�߂+��Z���l�o>�'I�^�1�φ�:���R�=�t�Q9bN�'�e�����Ul���)?,��"�m�m����z%��5ή{f.r��A�!�O�x઩�}�0,���1gz��8��19�U��UjF��I�D���E�V�OئfDO��E�V�7}��S�-���)��/�Q���^���1ɻHo�ArA�j9QG[�c?�˳{�i�lc]{��S�(��fB�����hC�? PZ�6�)-~�`��n������8�������-Y[3�&�E{�;�a)��[X���������iͭ!z4d~����h�Ny��ɢZE��]uP���ꝃ;�l�.�]�cY������#��|�����"������݄�,�!���䙝A\N/���u̾�2>y�F��ID��Lo�'�n^h�L��T�"��^c����G~�\�R����X
;����Ŷfg��~g9�@i����n�o�w���B��&��,����׮�WFx�����S�����k����Ȅ2���b���wo|�X����T#�hdds�� L�G�	^�tl����ΥC�1%��vޙ�ח٤��6w�����L$R� Q����r���σ�����0<��0wa�7	yb(�o6%~�y��Ѱ]`Rcn/#�J�EY�o*��x��C�gE��(�yV���V,w��ۄ����&$���đg���V�>�݀��T�P�2G���5Y��uJ�OSW9 ��e�����r�f(J(�y;�����Lt��$�	�09�K�	���/�!''"�	���$g�xj����!��$�@��{!��h����ϧȦ�!��E���L��m��+RH���,�d���~���Xz<��&5���ﱉe�����"m��t��rU��7��;��<;_Y��Z7Q�b���ZuV	���>�Xt��B3�1��� s=�AJ���s2h�hl$���_��$<P[r���Z{�+�),��Fގ뇍\m-.pĈ ��S4���W��1YGȦ��%
��u���a���f[D-�$"ݒ~O�G._z�x8�H���׃ȧ�fj0[����U0["��U�K�)q�����D�������p=�!���_��1l�bӹ�fgʛ�{}$���Yሥ����^�Ôb��l�$��;b)x�]<��N"y���H�3��9I!��=?�>RR`(g> ӡu 13O=u�����#Jό�>���K<��=�ϡ~y�j$�����C�|�"���3C���Z��}�H "/�K�6{Rk|��f<	���*�<��)�&@xV^(@|���ѱX���Ҩ�>�~Y��(6�����;|ů�<)Y���M�_���|����`c���hA�($JYcf���Ͷul�&�\lȟ��L_��!_���dp*y��}aR ��4���'N/cf�䙰��嚜 p�N0��b�hc?W'�^N5N��-xC��9�	}o���G�H�J5�M������'�:9������2Y��4^���7��)�KpM ����pJ�X�r%�����@53*�̿���]*�}S�~ �7��E�lIm����ׇ���է\RƼ����5ج>y�}V�ܞ�K�3�s��qctA��Æ�z���m����������o��դ���Y�H���K�7��1�S�d�Yֲ����o�XY��(�bf�[gý�K�Tf����W��<��p6Al �ߍ�U0�?�� 2S��T���t	�To�l����d0Q�q�Ye$Q��
�;�j�D��A/���TM��s���%�Ѳ"K�O��z ����J��Sm�Ύ�]��hx�yR��y�Ys����k.�8�f�������z�x�]XDrz���(�g-�|�9�<�:�d �~���q��.���6�r�>F�3)�z���a�Q�5GH���M�}��Ad���6J��]v͋����u?yrZ3� na���,�/K<�����
�0u�Zj��P�}�y�Z2�ɩ�4�:ɇڷq�x�>�-�s�A)- yF�NS��]�𙲪��ǹ�#�4oP�˃��[�i�[�*ę�'�z� ��=�J0��;	�8
��2��� �ZԫcD?1�yfhs�U���<���ݸ].ƈPZ/#ު���!�옛�k���<���~tAK�2�豊x�=G�*���kጓ����4����䯉`�-�vd�HaKh�p�Ôݴ�ZO�c�R~����T�!ހ�+}w2�G�П'���9#��u�X�<���\�4�	�D�D��^'b�#
Е�~ޝS��Joq��X�e���Hb��! ����vpi���!��%%arRk��� �r��j/ǩ�䤸�����Ɠ�n�/3Z�I�9���-B��Ti�)h�NL�`��G��Q/,��t�Z�7���_�>����Q�҃6��\
��`"�3ۘ:iA�@�ք�LOT�_� 5J�9>;�9=�a/2ϗZZH��|�1�En	�V���q����@�C��wl���z��#:'W���u�u`�v~�ݎ��[�M���Z�"�0��(k����a�$[�&�'��UF�T�[ڦ#r�Q���wA�)�j�a��uB~�G�����2�(�]�d��1=>��c_Z���I�K�Wv��zyc����L�i"��6Vj�iv�H�F��d�(8�>L������/Jr�Y;���*A�����O�1��+�7Sۢ(�����{	Un�x~��><�N$A̘��QShq"�a�L��C3��r�V����o�z(5C��ޘsi�O���$�y:K�"˘����-4g�^�U�����)d%(����2�ZB��㹼�g$����S�@I�A�i�.~o���X�hѕH>�j�{�#J�p���;��OkiOow=V'�����"�'��U*4V0[��y������V��Ϗ9n�u�s)U/���𤣃�}�Ⱦ���ݚ؂6Svv�6�!�`���s��i��5%G��vq�Ԍ7�-�4޿`1�v(���2s4�M�����2�Ի��SaN!
��%c�g��=�?#��4��xD�u�2@^���kG����|���:���T��?�ꐌ�#v��* ���r���,�D%�d��)�{@�9߮�gd=�*����c��T0�/e�>�q������Y؆Tt,�]�1F�]�(�&����1q!���M#�*
\aMf ⥸�WB��`d����]HK��H�:�g�X�3�Iɽ����m�S��o$T=����G� 9��2�t�Y1e6"/M�Ag�'���k���{#��9y����nع�:׋�3C�ˊ�i��_�}���l^����?~ʔ�0V�v6���F�x��_Zp����AhQ���W����)N��jS�u؅���X;����"G�ΆRq��'���B���-"�}�_ _�E�A]��ҕ�sL�����,[?��X�Kx,T��w��Vh���1|T�҇;����Ѓ�`+�� ������ʟ��:���5�>B|CjD-�q*�$�)90��v"g=x
��k�m�� ��rE���\bJp�B�|�%���	?�0?Ⳗ
&RL�N{��N8�%k��k~D*_ic�s�i���?��B��p+�I�
�:���z�p����hU@��:: �y�o�%%�TS���I�t��!昣>z���w>�{�3�>���T<���l�����|E���Hߣ�%�f�:x�v�H��/:��8ԺI�9T����$�Z_#QtC(�� JQ	1Ϻ�q��[��J���kP��$^L�s�8����xr��@V�$�ۑG\���y�pz��%� #����)0�x�H�|F��h�="9���(�7���1s�PI��$P�Y�'DF�ӥړg���?��Y��@�N���c6���vwM�!���H�/�� [����k�ؘ1�6kE����(cXн�<���
��Jx鲪���گ�v���+����k}]���ܣ��7�E�N��nd \�M������m�%V�q�[s�^�.�UBA{� 8�M-[�;o��+��뢌����f��<�q��d̺�����P|�+���Zێ���$��D9%�A(&`���>�#흚�;�r����m��?E���pHUx_��~n��m��=�ia��3�	���TĦ�;�%a��C���d-$!X��Bn2S8��=�!T�}�����^�	���I�_E�r�N�9��f�/�[d��h�F�jf�b��o�]��_�h��xe1�<4��ٕW�bBr��+�6Ny�!�8{mQ��ƕ� �Ob"��7�������iLо�
�wwQ����H���rKz��d�	��B#u7U���K��;oDߤd
���=�$%~�j�0��".��̖�����4��0�4y�La
C 9��Jn�Pb�rN���7�sy��~q�x�4J�\S�ȖPYsRP_�.v�i9ײ]Ʒ�]Jl�-{{�m��	m�d�������vM����{�'�w�r\��jXC�\���'�ϔ��!鿁�vU�t?uW Z��xe�A8��!u]� i��W �g�{�������e����HZA�,�M����g�g_C�#9t���̖{��A���������a�T���1�A3�O�6ƹpJ{�����Z���1Ti��7��8�]ô�O�%Rp��i1�"���OT��yV��G��I����2��]��9�)�{��M+w�������O��Y5��f���}�K!b���t`9� ��8K���ڳ%j��8�i":�:�Z�H�& `V�ږ�.���=_?團��С$��aW�+�;�5�m�_��A6�%��8��ݝ�G3�\|��6F::NS[��o�[%<�c���ߩ�Q���?����Rnخ�9�3{�,Q> �<b����ꦪ��� !ھ�zf(V2���:����v�<���6������|v��vsq#[�[�"t+���JԬ_ot���1�,�Q���⟍�7�3�8AdW83�u��񛏕�V�S��](k��`�LU��ϧըD`[ty-(pB,劉-s`hf���������ڞ\�[/�ۚ倰:����O�����}�F�d)�=ˇ�Slo(�Ѽ7>�v���	�δ�)�(�K9W�R����y4W%�:"JMЋ��2��`��Rm����%�����9�jY��%��Ყ�/�B$:`e�V��q=`Ws�h���o�F����v=�P,ѷ8MW��5cЄ�-(�� �U��Sd�J�=�.�zf)��|[�jJ�UÃ,̊f���=��r�>�������[V���AiAh��Z�!U	�̵_0�Zu�-�6�	Z�G?ҵ���-:��$��0eJ���#��u�Ԃ�G�����	=@zЕ�+xC>/bGx1���N�h��*�6�ݣ|BO;q��N�w���xM�d�%(���媉���I�}-�?T�*2U����C��a[8;�y�<���o[��U�
�E��P��hm���IV}���##��&�q�~-� Ϲ�s�ezQx�f4���HV\��~�R ���KT�e8��oT*T��	|���8��.^�A�ۊ`����G���:�K�!�d��3�#�=�,Y���ź���x�Fp9�G�J��"wpdR6J��c�_�լu�
��~�K\����N����.E��s��+��q�v�Y�վ��e�p�=4�ѣ�5j�|�a8�L8m�ơ����2>�y8�^� 
�qضr�?[��{.�CͿ55k�*\�ޑS�ݟ<��z��!��-�y����Z���+18���!�IԘ�d@! <`������\�n��:���,uVq�����_4����F�$���F��Ԁs�[�⫨������جG�Qigz$s$�<o�u�{�2�u����?%��(S���(&��J-O��Gj�b�P�;�7�π4��3I�suJ�������_1�MY`9����<����z1�5�Ƚ<�8v�ʷ��9��������w]����3��`JM���1u�]�C3�/î�0!��|k>�F�'TL]�6]wE`�2B>t|z�i8R �"#7F����;I`h����6�p8ө�;�c�# ���4����63:�3�T�ו}:i��m���G�>���X'X���"뎅���c����{T�HR���!n��P`L�秩1�L��$����/d�7?�P8a����<�Pd>UAY�mR��㍙N��~	��H5g�����iY����������mY���-Ľ-�ߊr)u);�+ɠ���c�r�U�p7A*Ph���ֻ������B�o��[�Q������R���1�6�0J2@ۆ
y{z�x����fY�A�
i�1ü���Y��zaP��CG����O��C����\'�l�m�h�R�q�U�Ͱ�:>H2�Mr@�D.I���.��0i��9J�7�@��,
���;�c}>�1�|6��L�\a��
��<��%%�򲛁����g�j�ͺ��g/ښG��HF�|v��Ë��$��<�������F_6:����	=�qY�g G����\������h�<���}�X��o�`2�ᇴ?��@��YL&J]��E|Q��l���Ւ��!��sN����po��fo�) jJ��0�(�p�M�)�	=`��'�j@������]�d��Y�~��3��r#m	է�a��Q���g�x��~���&��y��C���o�OO��XȽ=��LQ��E�4��R�|�]����^i<���i�`R�d$'ݷ7�{&Ӭ5��z�_Z~��TG �{�FE�� z��Q�O(����#��Յ���9�B/p�$T�4z��&�EP�,�0X_��fpv+d��@Q�h,�QIrȵ}��fb�J�vV��E{��:�)�s$O�ј�Z)WIP��6�(f��¸���c[�KE���~��z��I~b��3#���`+��n�t;���nM���be(�Nd5�w�ul�t� _z�n�Tm�ҫ���!U��6���������r��M�{5x 8!n���#'75��tm~$�AjǙ[�����8���2�C1�8P*����U�Ii��f�L�lY�PO/G�n)E��b��r��η�{#R�,�u�OߣXIZ��Jk����`�G��>�1�b���L�z����<��ѥ>��׭X���D_US0��	^>9�hDG������G�ᗤ�(a	ޓ��8���>P�@U���������F�
���q�r:l��_!�"�圷���.�I\�{cnf��_����A�A�N'`ŠD�h�+��X��1Y���wP<�$jzs�cy\�ˣ���I-��If�b��C�L��m4S����.������]�4�wc車4<�Lt�&�$)��'M�GЩ;�kJ���A[��.:LI͌��=��m���6���-�I��N���;��d�J��9�H��I��_�̘�Ȳ�f���np����}F
�Y�Pnt�]&��!}�v�tb�G������q"��k���G/��Y��845|"��	2��n=��?��\{��m�0�}	�C�L���";Z��($�!�jg
�C�h���������?�]�;8��U�(��cW��5s���{�������\j�u]ܗ�/��w����	9�k\� �/�;��VV��f]]��O�&�\����%���7�������Ћ5X���r�YX���K���a�W�nb$��oR���S�Yd��E���מ�+E�5���2�Q��C�3��9�l��:�·έ�Vut�;��rn�J�P{V��������H��@��؜�|,?��/;�ow<�E����/���*�������Fے��u�v\�����FYg��?��!Vcԭg�T5�2������5��uNOr�j��?��2*HRQk>z} �����\=ނ� ���m����W�V��*fʍ��T'���ײk������w���"�ڦ��~H�ŵ���@����6Q��!���}C���[D��}�$뾅�����4 (�z�Ӧy��~9��	�;�E�z���Ӳ�"�(���>�B�v��Ap(Q?��y������4� ������C~�\>f�Jw��naڋ����e��ЬNY:�I���lk���e �
�ة��*K9$��;.�Y����I�KA�P�S�b��TQ�|���ݺ���2M�s�o��_��;'1� K��M�G�ٗ�4�9�k}i��A`�".�"����L)�K�Ҭ�m]_ oz�6�X�"��_�$X������� t"����uy �O?
���M���,�X ��9ٿ�'���P�N�BӨ�r ����@�K���*>[�qڽ�V
�6����/�I���I��k���Ҹ@8���d5��6p�rN��ʨ��!�B#a淯��	�YQ���G����\O��Ga�=<�A����UQ}���N����81W�(�FI�t�ms�����ִ��xT��:=�^����Е�}� Z���lb+�q�g/6Hcʠ�AӰMzj�O�: �Hw��S��_��H�~����}�[-�@R�u �S�y�/#sq(�O���s�6`�|70�D?y��p]b-����|NR�׸�oY�E�Ϫ�|`�
|���+���� ��c�v>q
�B}Ƒj���\P%���:��J��M�\�0k�B/ҡ�MN;��1��N��g;3\�pu�����?�~�NE8.��i&r�����_�����|�)�=��~�J�u������v�N�� �b��0f����*��w��C��Ɣ��Ư��-l�l�R0\�K���Y;��{��:�;�Պ憚��>���n�?~W��%�k����Fe�bC0��{�4�y���UW�+�Ph�f���:N�,b�+���^[�B���=��,*`������Jn�P8���m�y�@�>�P���Y��_�n�K�m"!eB�X��y_���p�>�[��a.�q�fz�ָZ~~���:�";�^I�������m1���[4F*���Sa4o���^�s�P�EC�Y���mh���x5A1�����4�cu�_�~A��T�Z�Ri��7��\Cy��X�WDH�RJW<G�5�G~|��1m�C;Y��O ����&�)��?(J�K�\��U��ųA+0q���P�l�do7�������륣�tW31�G@�T��G��������"��g���!�
����|��Y4	}��+��7$$�b���5c%v��9�}Ss��&��Ab��μ���*lv��3�&:�˗2������+:h� A���:��*����|Sib��km$�I�\�OƟ=@즳c�52�o�JR�!#l�n�n�^豖���۾O�j/*��d�l��<dH����������8:X���Vwc$�E���fG��7>H?_ΐl��{:�M:èw�*=T����)�s\�޸!�*&�$Ե�,QQ0��&^���{��B2d��l\n�+����5��0���{�Q�G�G�ҝ�QE�@3���C�����Y�Fn���8��6p$g�N�S"����:L����bp)�;�3��R�fC=�H�q?>�:�ρ������{t}��Μ�������8i�M�pۣ���:�{��`vrE��<�z�����tm]�V�)�ל	p:-P�Ƙs��ub5�u�=�M���;�kw�L<�^o;*���p0�`������4�w@����f�U��i�����=�L��p���������Hk7A�pJ�7����ƇX^8���g#c����Yf�x��N����.�~�ԣW=Z_�W����ܽ2Y��i��J��+�ռR��+m��b�cT�^�_�[,sb�[�o�iw���S\5S/�~gb�uH���3��*��<�q◘�C'�!(�,��CH]�mi�N��|���+�����4t@�Ey�2'1�?���(�Ѓ!J|AY��{TnN���̮�^�E8|*3��?�g1��
B̗0���LВ$�4��W��N��赘��w�L��ޙ�$��)[��g1|��M/J+�gAK��V���ҿW�LW��5vP����C�����##����A�E�!�e<��ˊ��Q����5����d������N���K�ġ����7�K�̝�=�s,��3%�d�(��o$�L�_�i�WΚ��A80�G�	B�$$Zw�8^	}����/U��+�i������"���E����,��^ϸަ�-C�|�A�'���Պ��mbo����t+��t�t&�?4�/9�+ӭ�T�����{��D�Cm ��R9��H�3���\�]�6�x�|���u�\x��w�������X��2��f�\�k1�R�7�vZt�M��{"��w79�i���'ٜ��N���CN���飪F�.��\Q�﻾<��|�'�g�=RT�|{N49��\��ݡ=�}��'�̅Ͼ6�2�5�9cR��,u�Np+!��q�RW����p�tY&�-����I�դ�1�}�^�# ���&���I}l�	�ٵ!�l�1k����m@�����)'����o����Ǎ�|�`.3�F�����-�QZ���O˿�/��%���	�����)k�uk�r�jc����t�.T(D#u� U�D�Ѝ�C�l��>h����^	�*��_��e�� O��4~fl�c��L��şp�g�§�H=�a-�v(u��{�֜;5q:&j=���:�A��*�9p��V|�T~������.���f�l��u��Bm�Eܭ`�m}e6�pV���l�AX��)�ש@�3��"�K��}Ƕ�7�Z��K���L�[U�� ���&����w��q��WM;h�W)kz1 [�V��s
�-i�Y��Y�����𐝚�5�"sS��!�p���
lm����*�b�b�� �t{#q����_�f�s)���?�2�OA$�Y��#���y�˕ؗ$�M�_�%m=�ݬ�E�r�Zc��4;�49�
i�u��߭������6�q��id�M��J6ə0�N���Ź�or}�"|�a���?m݀�A���Ù1��6[��>����B#ؐ���q�Z���3�'4�Tj�n䙔L����f��#��1)�>�ت$��lt�_���Ga��3��f�!�ix��l�3��R���Y\�,��V�:�n��������\����x�N,V��&E��U�ALSg��؅�$����T"��3���u�SXoPo��n���u�A^LZ�M �;^Axw9E�.E�uj:������+.�6w`�P̏=<��7��W.9J���:�8�;Ѡ-����(��^�����*�Rv(�h�)��ނ��q�2Lc�@#TKs��V��eF�4z,Q9��&��B?(�~�ͭk�J��z+X&̓_K�"J�X�e����hR4f|\���l)����Ry��ܵ������J�p
{��2�?7�o����/�'�Mu�����Bd�Ӌ�7v�T�z��V�[H���r�����WAm6�Ć��G瞕���7p�pô|����3V�����y�%\n���Ur��
4��fV9��{P� �m?:��x��c��ua����Z�$�>V���Z��O��
W��ut���rZ����a#��/Y����b$/(�K�����7�ސ�i����X���d\*w�!}ڐ��xw���R�W��&���p�4%��3F��AvNCnܮ��$��BI<�R����54��U����[l5����yG���"��WX�}��nO>��)$w�Ӧ!��7�����m�܇�����xf�&��L�+��~��^Q9���\��zF!d4EE��������Gy�}k�,]�T�y�g}[]2�44)Mi��ӈ-�JH�3%�.��'q�6W���MFg����&2��[�E"֔�1g��+B��}+#j>B�h�.3s^���I�ϰg��k�֠��NL ���E8��2X꺖�^����f�)��9�����=,���Ck��ɏ�<�9�+�:)��7 1YI���-���Uor0ī��/�Q�a{��3�tRR�E
ȕ,�̜w!e����G&�R���	f�g��u�:+�xȴ�`���&0y3kѥ���F�A4������� �1�--lBXz���	�S���~"��}�1X���O��*}���Ű!U������	O�J���;���O�FUM�?��z���ԁ��B�X�8��r�=G��b��`K"ߑ�l�t��'��q�
�R(%ON3xs����e\�󷢗b2��f:<w���=��S����T7S�ZPֳ���W��e�A�߭CD͏�%���_�Q����S-B�!q6]ʬ!N���=尃��e@���o4����ٷ���^�fT�#E+"��t�����_Y�I�`0���k4c��Q�]<˄4g'3�F���q{�B���z�'�N���\�2FF�۟���.2:��/��v�F{o#�4q�β�N�E+M��U�3ʑ��Ik�\_u8g���cW�@�]��]=
J�T^�F[�~�u��`gw�B���WX�ա��y����m&�Z��2��X/�L�5� 7�����Z����Tt�ג]��ꚱ�W=�Vg֜kx~)��?E7k�/�L��ց� ��`^������f�_w�+U9��2�%͜�p�-v;�������tǡ�&��tn��P����[`}zo�f�ks����nq����S;e��l�hn �g��F��&�u�g�d�m��~���#���(���#�j�$��$��+��z��x���C���cWZ��d� -�g��b�V!B���i��CE���@K��?���m@G|q��9�n�0�P����>����r��z���KI��7Q�O�#h1\�Pڴ�I���~�Q�	R�4�x��]�촮��'�}*�D����e�cv7Tp��3�\(���P�ϲ��W��;�t֍ºu7bIlP���;J���b�����GR�d��uQ9X7BB����7��E [bd�ޟ#�ki�bCK3A�?	�7Y���&JR�aIڏ�
�^�
:��EB6b�ȐiO��s�Pp�db���u���������V�����xbD�dS�UA�<�{ޘ�/�a�ؽ]�[���x�)����H���
��:T�̗iRP# 엄2�غ����w����/1�X(��%S�:��.G�P ڒ� �r9fyQ����˸`60�I�0�=L���Ѩ��8�J�ߦ$F��Z���Y$��D�t�S��U{����n��!��8g�����17����$K��n�$Tg��G�����Qͳ�U�	Y�C9�E� ���|r/Mx��]�m�$d�u��^ۘ% a��[���O�`�ܕ;��;�9CWaŚō�l��;�;��"0�,}Z���Yw�s.�O�x�ʹ*��7sJ�kN<MH���:��r�(�x�2f�{@HhF�`��8�d]{.:�lZ���DR�Q�x�I){f��h{K�@"Đ~ ]��> �'���cuB�<���Fo	ʝem^��'D�Dt��"��1q�'� O�0�}n��&Gtpr�W��f.���J���q���5-��Л=�px��~����Vm�/���B5���ã�u� _j�o�����t�S^M5�p� �#D���`���R�2&�X�1����T�$�����"$����S��ʿO�}ۼ	�ȋ]5w��/ף�Nu���s��޳!m�]�v��^#'EC�nX����v�c�$j�����G�4[��L�@R�������1�ɈvLyS���V/g'I��c*n��Ar��¨U/�g06�Nnmj�U�~��������Yb�u���ɩ:���yiAbW����R'�R`R��`��a>=�u;"@ck>ni^��e��V�8�"��O/=��W�e�0�Jg G���<��s��ᒂ�Ѿ�3����51�`4O���]��ݶ��0nh��kK��Gg��YY8��7N?��w��lh�D8[9� n�;3�}���CۈϏ��Ѣ�eHU�Z 8�����V�����P$
X�>a���L��i��0����5���^w)��d;`����4�T�n|:��O�B������H��Q{���<�WC�x@P=��9�H���Y!Ib�A���Tԉ0��n+��{"x2���~3�y�^oDF^���JA|h�R�!�D�'��c��u"a������BՖ�dVF�y�5�*�{E��(�h�~w��|`+� �y��B}_�e��v� �cq3�{kD����>�۹�Ʋ�q	Y��}�;IG��L�M*on:ה!}�f$b�
���	}0p�
�h�_����ݰ±�"�,j+��D�I�O66�z�$��D��pV,?!��q�M�<PD�8F�ƕ4<JRWzy>�il����|��e�:��rL��z����u����M�N�M�m�����u-wҍԊ�M��`�Ȳ���dL;hqK��t)�h�K�?X��K�>L�o�ݱ.
�3Vj
8CO����{"������ߜ�V�9��g�O�/��VH<z&���XDdJ��S�gekO���L��3ke�����L;�ʋ4ˇ/z���nS��+����U���	[���&Rz&Xm7.$n����Za��͓yN����R/M�K���K�lJ���S�����ڢַS3y�}���-�	 �%A���߸�ɐ���E��/�*�jSO+t�t�����rqڋy͜������^��]yVdS��\A-���5����,Nݥ�3������u�ؘK?T�C%�د�-�����
���4}��0Rȵ����PIZ�5�p.PX#kG�Y�O�B��;
�P[#E�����6�8���b����!��Pqq`���ޫ}�KHsIQNhg}b0�5S�q*�4^f\[�Z���/��Xi�@R�p���x�7k�� �;(D�c8���#��u��o[y�R��`�➪f>�G�������"e��H���@�Ǧ$�G��ʛ��he���]T����g�8�E����{}�'q��zG`T���m";J8���Yv��Z�=�s��&�c�Gf��6k�6�=kx�H��t|���[I��_��[����`����7�,
�C��?'%9�?~Y��lUv�D����t�Q3�%�M��*J�+r2��������
�c��٠�i1��v�V�<�LQ�ުFK�"i���z_�+�"׷�(AR��g��nz����59C��O�T��X��}<�V����
��;�� F���"Z��lR�H��d��o��	-WKQk*�g\1��o�9��$����tdn^�q����ġ,v�~G��m��	�񮶅u��q��d�bb� 7��|��E�5��O�c�!C�I�����yw�g�T�m�������I�C� �ޥ�0�l�]35���O��o�}���7����4�=��d����h3!-��xo�����qJ">����&z�`4�X��T�����9�Q|�Nr�< iָu�k�C���~0ǜ3��b>��!�V�O�bۿ+�
�@�~��ie�U	�m�х�/ڊF�b��ə�}^SsZ$�.QU����:��,O#��eT�,rl�]ｋ�(څ���|@���nE/a:�~�.��=8�E&r��2�<b�r��#���e|�)�h0��S�]f���MZJ�0(d6C��'�� �k�Ҋi�q��4��y��4v�$/���1>������+Һ$�Dw�B����U��ʡ�8:%Rw7�/�
�'���P���/���5�ä�a��z�O"��#a��E8��x_
�n�Q����`�@�b���$z� +�x
�� G~U�<9,\GÿQfAC�jl��*�p���6�U�Mb�-�i���$��+VS�1xgO��nc%���,������ėK���a(9A)�O��;I��2���'��ȪOiu��t�J����6�;t��S,/Gv����KfFK���?gt�$]����;J��X_2�u�5�2��&�C|1al��A�36]B��V*\��%F��Hq]1�,��Q�"¿�����u����t�:h?��v���lcIk���&�R��_J���	���I�fU�+�ѣa������ތ.<�@��k1��@<���)��f�;󐭰B���o+a34�1ku�(@�����9�l�%eF��!�|��������kX��Z����!�[r'1Zh.�����=�	��@sR"1���H_I{m)�7���}|�oЈ��53�%=c�F�W��-��=�	������<o��S�fn%%/����(��� ��]�H��,^S�m<��������O�1������,1{ߵ2G��ϥ�hC.L,e�"�S7P@Qf�/�Iq��eL<���4&�r�+'��@B����%1���q~\��b�6V��A��-k��a�VS�
�u�N��kp�ɭ- M��v��2v�MI�3�	t���A!��Ύ��XrB⋥���AC Q���0V�M����FB��N��} ��ASj�Ѣ@d�#��'��q����_��U�t��6��g�&�C����y�Ry5_`vO�aΡ�,��o��b���[΋Z�e�NN�Z+RpZJ��	�3�čڤߧ�A���j��6qM�J���g<���U�酝��j#0���>���9?0Ǥ�@�a��ݍXߊ�~�-˲��ﶝ�gH������Y'`��#��ӎʡ	��D��7���)�~�QHLH�� y�	Sl���G�lM�����������4�e�m�V��<����I[!����S�-��'bwM��9�Ag��2��=j�,�u&�qKYe�vH�(-s�$���6�!Z;�`-4ĵ$���#"i.y&�
ibw�9~8���4M\\�#�)�k6Fe�Kb�qQ�j��&"�}��V~e )~�ӕ�=Hx\�ݼS\�T8�G�i~O��b�\�,x��)��*"9����3��l�������OC��(�����T6�7���Ri��#��̔l��|e�>��Q)7^a��
��FZhM5��Tb�z^��ms�.!y�Nf���U];�Ͻ1-'�v��
�<`Z�-�2�����M���I�0{U[�?e�^�!� E|̉�]���XO����=~!�QGQ�~���	�V/���4�c�Fk����N,TN�g�
�[�3�;�jJ�sƨ������j�2K������ϰx@C;$��W�#؅,�K���5`>�/����ڎ��tjȄY�a�}��x2^$�d�wе��i�h�_sܩ��+�g�uA�5��JH^'Wi�5��O/�h�Q���E%Uy�Ԣ*6���J�c����z�F{�F�����O,=S���* �L�^��o�"���*���ˮ�Ed;����O3�)�*7ҥ����'D5*4�����_����zU�ӄ���#9��m ��
�5=ž�0�+H�"�V��(���JP���W�)?�63���~3Em�Q3�
�'�.�A���[��+$��j����U��qyJ]+�y��1h0�؛{0;�M�En �  b��:7p�s�)V^��Db��n��:��_R���G�Q��K5����<_��w;qN����`��/6���Ӓ�| |��f��c�x�e�m�6��j/����VR�����lS-��@}���p������[7|��oиE\�D!4/@�SԮNQ�.���{	!�:�Ԩ�$G0�fv��4��=����\UE��oZ���,G2t��ȶ���e����9Ԡ��Lx����%��d�*/~aI�]���2����;�a�x��E��G�W7GB˕�醨���(|��a���%���oڣ�R#��8 S�o'\�w���9�ƫ�|}���/�EG.d�X�&�	�e����dh]?t�~�tJw=7��Sv#%��zN��|��l_@<ip.��Z0+�R3���#J���l�:W����C̃�8Q\���