��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E��S��;z��Q��8S��fʹ:9�F
L�~Tbr�)	E�+�@|'|�;m�
�K����D��T�J�Y9��n��nw�,����2]�X����y�\V@�L�F�� PG&�O�.vCu$���N����]��\$�Sg�� ٤�/�v�g��âAq����(�~�o�YU�gဧ��m-`��3$1�UC�Ő3�2�k�8؊�����Bc�1t��f�1<I�P���JyQs��B;2!^)��}�4�)�*9�/A�Nُ���F��� o�7�SRl�
�8����,��8Ҝ�/�v�;�}ԭp��e$��w���J�v:FU
�~K�L�[����uڨ4�ܓ�y
�N�3�������Տ�qUql5fUpoD��������p��b�h���Q�&�x�r7�q��O�6r��8�����/�}�]�B����#���R��'�*���Z��:�E}˴�R��I�WRD[�_Wp.eC\�[�N��C���i�z�o�҈�ܷЏdS�B�h$\��9�=����j�n�����W@��כ��g�0`
L�u10=)N��,�I���9T��8��i�!Y%��i['CaG:�����>لf���B޶�ώk�L����ɫ���r[������pשC*�h)y�i>B��5}�%^J{�E�-��G�f�<��d"x}��H�Z�M�&�k(��YlUQY�?�D��YNZ\�����^���E~%R�և�a�0G����2�\�$9��ȹk*Z�9mLf�O"����N�����l��1�ɹ�C��VD�FDI78j�:��X�Єz%��?�p��\���W�#;4|�ل°3��dؓh-�-����@x�-��Do�O .�?t80,��J�8u>�%�f���bLS���U(?���(�Y�f��bj��0Z�\4�E{ î|v%Yi��I��.y�a@|�4�1�,����A��I�xo@�̞n�Ա����襫�,���-"�a�J�u�M�W:+2#:5�]=]Bk����=c�Pe���'w��3_ LAŧ:QB:Qd�Od2�ƴ��H�!$��N*̐Ù���s�Z�C�.��Z�NS0�:��L6u�1C��y�=>�i���oH �;��&5G�8�SM�ݔ9)�z~4U®%�I�v�\�'��b��jj�\�#�c��:&���4�/�]���.=T[�OrN��ڏ�[���U��m"���X��\���a�	6��<ޣ/Y�_ɶp�iÖ�cb��;��]���	��	X�z�-�H4��hKܭSK�����7�LK�:i�i���3z���S�M(��f0����yu����l,�������[R��l����S��6Qjm�:95��< �M.��<��q�~�ӌ�]K�rͮ5,���i���By��U)W4�� N>c�(���@���wrv�45�Q���A��������N껟�����(|���W�7rKE�p�w�q�Ӟ�g<�1ێ=�x#&�@a߇��Y�y�j!����>�z�wV���6~���ݯ�a������h���,��7~h��{�j����텣1�>g??��UO����طlA1�Vf���������"/l�m�=�ܼ�s�SK�w�\�����\�%1�7 D\���ԓm=��[�ޅL�u��憵j�}4�Qfn:��=;o�7d'QÞՐ�U�ܩ:��7H��ws�@?���4�yd�AōQ� F���*Z�Ie�-�����Np̏!~1J��G&�g#Кb|�;k�W�r�����~fN_}>l�4�?��pK��jpXmⷙíC��6b`@c�p�	��1-��4T�iq,�&m��&�#�	��ֵ?Ar���k6tɰ�Z�em�O,�R�n����c�B��*aQ[�#�C�#K��GSqte[dd��a�~��N�tߋQ�Ũ � (�nr��h�3���_a��������Б�����@���<�"ރ>�{F:�W��p�A���ީ�E�jy���x��T.i������>R���p��&"��R�ΐ���@��2�]{��0'�';�����p�Kz��dх9/ n��A�mM��8|;�y�)�Sz��_,��T����x���w���B|�X%���`X��ci�4Z�a7,�%\[�s3�V�)r�'� �q�Q{���-��f�L	����ܛ��=�5��K���e�YUJɞ
�'>5 m�J����v�F�~B7�:�m[��&	�УP'Ќ<�|ʹ!����ӎ�-����"�S.�܄��ә�v�We�5�\1s��M�Օ��H��*E����+�3�ڰ~[�����0M�Ql�\eS�<����z�E-`1s!�n����Ew�~�x�u��ޑ�t��ߵ+�)y�!�PM�،���#�d:��Uּ��&z[��d�h�`������_c����&3���Y, �_3�;�r�Օ8�)S_zt�@�>��	:� F��j��or0|��M'�%�Z`�?��"��� A�ȏ�F�c���i0�J8N�#2c�M��*s?�JȎƉ?)��ԟ�����P��������;�i*O�����%6���͂�ÁŁ�pN&m����j�fo�M��1�}+�	��&������E�uwa��������=�f�vTǛ]6 ��o5%�z��W�mnv����u�m�َ�Ju̯�$�^Dm�[��0����,���w(0�>"iMx�C'�5)ظ��l<�9�UT�s�Y��կ|�t���w���];ܹS(�Ӓ��J���+e���V�1���(}�%+W0w[�n��1a�e1�x��=�2��T� �<���n��rm/����}���'�h���԰�h��V��ށ��;���7O�!w��z����4ͩ]*�����bEi`mbQ��Ok��QI�?��A�E�d�+<�<�����e��H�B�P��?��5�S�bJ,�+69�co W�6~�<&)B}�0ø�x�}��Ú����/Z��p�� �Z!��a{���e�:9N}E�>0�z�N���Sk:t��vw�����d���-U&��9t��4f��C��}�!�L�;h��VZ� H����a�Ÿt7V�Qn� ��]JO��qX_��~�����<Ϧ���u]�ۺ�ʹ��*T�r��3�Oy�Kf|�� 9T7�a1�!����5$�;Ͷ�s �i;D"��C��V_�k�ߺ8t�M��RK�=~ƪ�9�̐���I�>T~*��@O�I�9�,�	cG\t���
a/Q�]4�)i��>r?{bU@�[%]�!�"�?��@�����-�yI�2��;�q,�(�Fߨ����F����i$\�s���/a\a�$R��]5��P*&�ƀ%:��L�������{�}��oxҙ�\r|	YT����#	�iLE8O�N�3�?#4�$T>!5?n(���K���D� �إ��t/cf���u�o�>��w���co��Ǥ�&�F��zQ鮵�!�G�$�	�^�4��Ay����>t�b���Ў���h/7h�������|�t�@����~W\�.dddJ^�P߃�y����W�e�I���˗a/e��`�m<e�,������m��I�f���3J?�4��d��C|�]��`ML[?���&o9Xl�8�X4PÏ"�m8�Z�y�7c��	�(X�3*�X�L���e'����x��&�Oʂ4	B_�ЙN����~���R�Dv�VK��� ��n*H� �`0ǘ��&K��=��q����5�2O�dY�{c�+�B���ͩ�P�Ɛ5T2�jX�;�<�=�w�J��k6|��O��p\�>�2�	:�r\��\�|�+o��->�>\8G,g?�#�����'���ēY��[x�. �KZ߁�-lotkJV^ �X���0e縦+�aB=z�5�Y�Cm�l�$ O������<�}���A��b�!��J���"�~qq?��ȌH���qcUiL6���SJszZb>l��G����1T�l��{���(/����y����t�g� z�y K׿����9�#U�U<��5+@7�q�v�[��_�m�������Ӿ"��A���٧s.�kl���|�S���`��:�������V�j��H�{9�(�Om{w�B��jF�D-J�o�z���3Cb���t�)�"o��G���T-�~5�i-M~��obC���)p��]��	����%ך�b�f�4�L�*t	���k�ҿP�d@�ގ+r��@���׮��~�k妘������9��I+���_�G jNF@A	��p�)Z�?�
�h�T`ew��HwR[_�����I��ej�^ҕʹ���ϱ��?{Ң��ݛ��`��
�1���r�M0еb���	���K��z-B0�˵oR���E��b��ȱ�*��'���i���� �����=�>��.���
��Y�g�����ϼ_����٫ʱ J$q{֤bn�;{�ϗ�F_?� n*ǃ�ʌ@�3����d��[�f�����ul�B��+�=�w%�[GA���v9�\5�S�Ryn���7D��a�2��h{���lI\t�Ë�7�^��q,��kM�R*S��JS=N��� ��> Y�L����aOyN�
J���q��:ٴU��Y/������j>��ƾ���<�����C�⬴�����m	�3�[ba�����0X����JI`��2�U�ّY G �%w\|�܌iE�9T�/��o�c�G����_T	�"ل$�h��D��5Q�WCK�H�����Kl��g4+u����g����0q�5�FL �M3����í���B�����{j�	�+!�N�Z� �<�D7o|J��9�|��d�����˂�Pn��<m��/V��s�l�C���H%�y��V��nF�@�v-?�f��\�" FXd<�~Js)V���2�ߺ�p�2l��$�Eµ�"p*�:h�8%�� �Ҩ��:�^2����V�&n���*O](,A��Ǔ��e]�U�9	�cKQ2�ߥ���`Q�R�0,7���gvo���oc.���S ��H7��>i���rC�*$��p�Z>V���C��߈�R�bGq�����wj$pD�V\�sS�
�y`Qޠ͢KJp�u^�g#����_���NΘ���>�Ȋ�3(��
8c�)d�&�OG��2�IG��������*��`o�	��ߒL��ީp�|�����Z�
E��X�r�����[䛔��傟�6�YV�N��/]�ѱ0꾘��d+jQ\��	k�)�w|Wr&Q�������j����x:p���W��;���,��w@��_E��K{���ִ=d�w-%Р��X�?�����Ә�4�
�Y�&�df����g�M��a�Q\�%�L�jܵ�%}{�V�����pK�
����q��4��0���nK��N�MvyJZPD�18�E)o��u�c+��<��)�
��S	���	]�'�d�a깰=<.��1�1MF����Xb���A�qi`��Uo��G�m�)�B#�����(�8�����e����p�L�MDHZ.|M�C���Z���/�����gY�{ӛ�D��:�1�'�����8G��@�2կ���(4,��ifDMB��k�T5I'wD���d�A-l�!���?��t��Y龋�I5�bm_?�0����;wb�|�C���p��qX�5� s]���x���0X!n�5�3}TJ((�S�c�&�t�����^܈�B�P�}�T�ຎ&�s�M�l������.�V���bt�C���_����K/�1�\y�$oSr)�As��"=:�}L��,�\�T�炸�\�7���xo�����oE���(��z�@
Fd/Ē��fV�/��W
V��"��M@��C��֔9d��9���5Uu�0�fZ�R�f�0"|���@�cf�ә*JĄi	F���+��$�����ǰ��8�e��Q�o�a��0-G8���$cDu��y@[d�%h���%li"�%�H#�|
%id
�B^O9NQ�7G���xJ�8�v������Ƴ�ج�c�bBxYπC	D�.��kJXx���������]!u@�R�\�8E�`3�g�qH�_:Cw�3��	����BF���!	�p�6z�в���j�|5&�$WI�7'�a�sD��;g��R�� ��[�$ }e�1��򞁁`b���C�}��yn�t�9?R{���>��z>�72j#�&�wkN���H�9��T��G. ���E6���|ϱˤ$\e���3��<�|Cq�/��"��I���:g8��<8t�BU��L}l,tb�_���a���K�K��7 ӝ&�S0v�)�t�����z Y7,�����z�BP�&��i�Õ8�b�C��+�6@y�g|��?y���\��]��-JA�r���A@�!�<-�H�!=F�WW�%��N���3	����J�����ÕV�0��O�mĩ_�d4�M@�6�t���E䰅F�;�dgԉpbˑQ?J�eصT>��u�VM��vo���v�P�������y�*x���=L3,O,�.�2�B"�k'X�r��������.'��.&o��/]?>��!,��
N�}���	�6_�X`��*��-<��M�-�#���O�9�Bw��1$+���1����F��_�3�΢Ue�K5����DW�MhH;�pI��@�r��$G��pܗ?�W�{�̮�A[�=�U���9Li�
�e�W�I8^0��l��ߐ8}�zA����=Z�l��-tR'K	����<�����P/ջp���q�U��{��'�[��z0*\%���<�|l6Y�nQ��I-v�/4X}�� iY"Mn��-��Կr#~�I��uȍLd�7�)�7��\'ӟ��3�γWVЕ��bIK+�d"9,�P�1:�oOQ)�Q?0=]bT����8��0_;�,�v	x�>�A�~�y��9��n��B1&��]��^(��t���]~^�+�T���8��1���'�T?oޢ?�y��ig@�}n4��}�6��3��U�Fg+�j�3pa]�u ��uo�!�,�.)���n�����x�*�N�L&���e�O�Xk�Te��� ��wY5+,��fC	l�_?8(�
��t���O`�l~c91j+��8��G��ps�F������VKC�-�'6�&�]N�`�3�qOH���b�B �}���x�6r~�HE,���߰)�����Ʊ] ���we�Gmڴ����vWާʷ�C3l����tX��.�U��X
�Hu��H�F3[z�W���.�@�j�c�����22�𓃦S����^ՑC�͝܆чTŏB�����ј-8	|�(k�^pR�j��2�K��g�{Ls��3,X�Z�n���z���-�N�f��_�A�i��X��!�A�x���XԿEB����:n���I��.�{%�c~@��kҋ�/��%o�.���+����$g|Ӹ��G�8t���lȹ�
jr@,�Z,"/R��K+��������0;s�8QG/��\�{,�5�,��X�|�@��IR������:�\"�G�A�u�t7��D�б�]	x��c{��fÂe��xa�'Ϝ���~�-$���7��wۏjN������+��J6�ۤ4j�6(�{�~��L����� ���!.7�lh�T�TJ×�cz�y��o	�Ƹ��2[�7��,���ڕ_G�Ԙu�%�u-<�3�;A��:/�eF�d�Z�w6�[3ޔpF~|b6[yK��DU�xť�P
S�����B���&:niVX:�ڋ�Έk�Î���E�.�4r�H]��Ǘg��ӛP%�K�Lפ9)�z����>�Dp�2��69aɲ�(����]��dw�YoҞđs�'K�q����娽�vu8�W�'Pr낿ߨ&>Nv�Cs3�7{2��C�"H�b��a���tTQ���()�0���+Z��c����cN�J�ܢW�=���)Ç���p�[�v5����.{�"I�t��7U,���LŻ��'ɳ��,ʐ���,3A�m���&�@d�5��ޡ��VB/�������9�B�f�/���z5
��g��"۳.�᷁2m�X>M�Ɋ!y#|Äҍ[���E&yu>�C��7#>/\d�L :���H�C������3��!=p��R�z'4���vT��K�3JD+s��zἛ͟�y��ux,U�bߊ���%�g���o��h���Do�wR��"|��c�O%�3���츇͑ҋ���a5Ո�2rYk��̦�9�i�Fg���e�RѶ8�9�ñ�z�?����1������x�(n�4aޡU� 	����B��m���^8[�w��|�'�l�R��x��d"8Ίe^	dlGn�X��n�حP�;�7'�ؗ�D�V|ٚ�}����M���_S�����R�b=$l�f�~��MVȯp�nP �����������E�Q�����L��Z�T:ȡ{:���?�|U�u��U�.�b���kׇ�I�N~���j�&e�"�' ����F
�`�y0W�T�I/g�Ƿ���~�	`#��D}�Ӻd$�(�~���g��6X��^��:D��\�dN�CfZ"�¤�|?S�����;��HV4}�%[v�јX	˨#��/�iR��d��t�)��}:3�|� O�v���m0Q>����s�Z3E,��jm���(|�9�����I���#]O=`C��*OA|�h�EW|.���6=۱���/�@x��,=Kz�"�?<j}�|��n�%l|0����S�mj`�#O��S>i���,∐��FJoՌ5{p���?��0Tt��Jk脭\3_��\Ɠw^���6��)���O!ʈ������$���t��n,άu��G��_�Z� ����$��{��d��h֧�ST����/������A.1�/�3#?z�˩�K�47�uC�Q�� ���i����*���>�3�����No��]�0��eF� ��\;F�+	n6�h��'�	u�d)k8 �_�B�A�#q�9��y6�W�}^�7\X��q�2���4s ���a^g-�ZI�Q��.)N�Ȟ5J��2�/S��8߀�K��{��S���A���뱹h��p���{'�>��9���Ϭ���g!z��N1�v y�b8��9Q��Sv>q�(�'Ī�}$0�$HѺ�b�c�D��5����N3�I����*�2�LO�P~�~�E�to�I�y�6���W�O0"�{���v��k?QvG:9���b��#jpgn�뎪Xа.�y*��1�)����dbp��h����7��qks��){"�S# c���B!DS"T9Y{p�K�0c�~�3^��΁��_ż.g�KP����舭*�㴱�շѶĐ�Ptpc�Sܰ;\)ޢ=xqX���:��i�b.v��A堲Z�9>���ĀR�-����#��r��ɣ����G�i)O	P�Β��(bof ����Yf�r��P}��߫�ٵK�K*�rA'�� ~B��2|��������+��+�����
D7٘$߲�!]=�6^�\ز:V�����Lb����lѨ�ܚ�x�Hݻg�)������E��A��;�,㜹����|K���>6�|9(���d&������{`�_�1 �+�I+��%�$$��c^�V!�(�6��gt����H�`�}��:��L�����#w�QL}v�]�6x�`�Bޝ:ӏ=9i�����m�f�s��y
����ć2B�P�cZ3�x����ݨ pU���V!��X�J�r�X�����,xg\��f!�UX��c�ŭ,�nI��j�0��� �ڠ���jG{��~��H�ѫb�q�v��F�P>��id��[�^�NFC�d��+<��bL}R��ź�p�ǆ3�����';k��.�3�m����ɒ��#��/�y^`%9��3݅Y�	��i �iŪM���5�]�p0���e�glM�1*�^v�L&�g�f8��͸�ߋ��&��b�0$���îTp7�AedrL�\l,P�T���=O,�.��m�[��?.�HfR_�V����@�������)x����$f��L��X�Ǌ��N�1���X~ ��i,����j�ѫ�1���N��&�ͣ,s���a{�^n�#��ðIVjI@4�O���$L`�"��ʞڳG��b�Ԅ�F9.k��;g�k/D�棠��mX��r ��xP��)���G��#ɾMb.\R��{�bIJ�4u��M�V��5*�jFNF�|��k��_^6�C��y\Wf�Q2=)b�û)	�����*9t��9���tR0��+|-#_�<���	a^���/S��`Ů.���hC ��t$�G�d=�3�=��
���0K�&��8~B�\F(�����}^*[0��X��$�h�$�3��v��1�J.�p�f���,�"�V��e�%*K%8�!Պ.]=��ct�l�k_-�T��B[��9�F��%>��~�N�ΑKw�קY4>�4)� 
�Y��pf�{��pWڸ&�A�t�CΫ�>O����H���Os�ؗMۖ)"&@(�3���e��,M��yo�ݫiU�r�����2Y����qp{K��:]�h�4�Ps�DE�ٓ	����2mKy�9	i�3�p��E��� ��*7jŕ+�����E�{M�Gw`j
��!מe��6�p���.@^��yOZ��&��aL��!��5�^�c�|�i��e�������o��PA�a�
u������ -`Al-pe�0P�����(���80����^]yZ}q�m��#�G�k�6\u}�g4�8���zP`�}?�@��n�w���P�L�9����殛+9+�M�$���g�-�Q�.��z}����E�%��Z���hLO�$�yf�^�\bE������FOS+D})��e������3�'c4���f'���P��5�M:�%D�����&Qw&DBaPߪ}����K��n���5�p��e+�q/ݤ�� �E�@�.��ME|���������vh���@GX��y�Цؑ�[��鉨O�@�z�]h�r��#��7�����ɇ5�D�?N�9 �&���V�nN9�[w�D^!R�0F(�t[�OU���)ٽ������ጦ��!��U"����c"�uV�F0q���Ŗ��v�1Ş��e��.>NP�$�sl̫/S��|m��}�����w�3?ǭ��d6ڴٜ�Ip�Ud�<|���*kR�E6�iŝ���ʳ�a��}h�8��3�;'�z圽���X8�������[d4�{`�塋 �I#6��ʨh7Fa�L�%Jr"��X}u�(�(�XS0ͳ� ye�H�#5M��˰Oh�n�ڳWf6�M��/�U�c`-����o&���'��xt@����žV����J�����i��G�|k��W�0�9���^���o]费��p�&�1J�ї��r&�r�\���1}����D��_��]-i{�[I�t@��y�<�����p#h�yQ8j�[�I�e��Vx��W�m6h BAUL=GD��N�\Qȓ;@n��c��J�W[�N�Gʸ�]p�z�.�z�'��7��\<BJ*�q����R^b��*��,�V9�&�T��b�yry��_�ӱ}�m�$��鄑P8W,V��bĎ����A��(�������<��LmL�S�3,�_p�ci�5 ��Q�d��+�V ��R3�Qy9�́�^�d9#��S�bf>8����Z
���
���~��.����V��!$Np�w�d+u��[��
]�\Z�e��i�|�i�3sۚ������ �c�2�u�������K퉎De,Cʒd���#@�]�j�KD��M�rw3i�mal34�Kؓ��#E-���4��8���j��H{��ػ�G���u�l��X+c���AGX? A��n�O\i�[�����J����{ei�:8�d�?}C����ys_��@\�����5��f��y%x���e��.84���(i
�?�q@��`��4�k2�igqd��V�5���^�"^�z
V���c;���q�I_�����5��X��Z�5fw���Զ�_�C��蹽}�7d�;�E��Egh����C3��CI���;�����u+�0ޓ��G��c�z���:w��,�a���fdFP�� /v~ S�#u���� @j��qӺ�(Q4?��������t���˂$�˴�=a3��g��|.*
���=�2sAV�ß3�����X4�+~v��@�P��������ɎƊ7+�[}�{ٱe5-2z����sVGm�!���Ͷ�hƉ�٭�(��C�JQ��#,�E��=�b�ҥ��x_�?��j� N7���o�bT�Yd�1�,����kq�$\Zv'���{���9��x���!�����SP6]�SX��2��X�
g�'��������q�o4��/�	�!��I5i@6lU'��eV5%��cη�ĳ��N� ԹʙaNڨO�)���\�WK�q�A_|�g9��~��;I�t�(������Z��«���\ܩq?��^��OGCm�
$�fL7S�`�&`wE��b��&D瑙�c&��&�e_��D�/�l�s-�.B[;��0�+���Y�f�F�O\9�u�2�ȿ���XBC_H?��0j� �kQm�0�|�lb�7;�x�36���@s����D a��T�m&�'��2ʞcq��|�➩q|���ĥ�ƛ�+�b%��quZA�	y�}���m����WZ�D�C���L�W8�J-O,����->�芐����D�xKX�}�z8��[4�9S�"
�U�C�R:0���A"�J���F�T̵%�[���R�_�ĝ�J����3�=M�i!���/�Z8�u,��m�@I[��K����C��ה����q��u
��PR���e�� ^U���80?�o���H> �k�2�o��c|�h�oq������2�=�Vi:��C]���B7.�CO��K�|G~�Z��R�mC�ROH��̝]MvKiDb���I�k4��1T���&�]&���h��F�u}9�Z�G������w(^u$���d����u`!l9���sD�SF�p��o䑵%y�uA����R�Ts��Mxli3����9����@�S��ڃ��+�3F\Ysd_e�j���?��D:�;��q,1�©��a���諄�O�I[Χ��϶��P�p$8�A��KF��ߦ����V���9h�E���K��#OiG��Gg�����n��/��M�zVj*`?���G&}L�-�Gʑ�)�M3_Q-%Tm|A�{6,�/��r��� .�b%6�2������F ��/�1�7�0�b�~^�j����8��S�?�W�M�O�J�L�9*�ח�þ�~�Y��B������]+m_X�Ø@���	��c?ʚ��3MI�A9�~�k��˻!(ܴЦ)���o-I��u2۠�u?4F<� �L�y��*�d��A*rW ~��������E���b�ve�;�f�J-��`�C�ן	O�n�Ӿ���il��Q�����ޭ�����N�U{�o8%Bz߾E�	�ǃ����$�=���e��*�0����#�Y�W ���&�1��%(�f� 6��sإ��(��ʩw�iԊ�8���0?�>���u�8Ѣ�_m�:+��ߐc�pBh�]�a��M�w�3}Ϯ���ܔ{�w�^��%�`���F�[Z��yrX|��E�/�nz���Z�'��a������)>����S�h��0���V�12,�T\��渝�lՃAa�ֵ> _B��WTD�(�VD�y�X�\�I&L���k���0F�W=�6|�*@���v����~u�+ 7���Ѕu��/��:��hr����I1���ܚZ�O�\������T��6�MӤ��x�2|�%���l�<}p����A�`�F4r|�W���h���;���a���ϥC�h�?
�U�'���҅u������_��T��ƨ﹂7�(�?+x��h��^a0@�	+����Jh��,�F���#��p셱���Z�tdp*槢.���Xj�Z<#R�*���~v�b���dN��n�Ⱦ��;�!u�tGn��?8��N�\�����#����֗	Sp�~�&�d���4�����qQӀ$�j���$|��x��.����S�������A\`ϵ�|;��Kx��G��JX����Z6H	&L�;���(�
�K��kX������)����u[H[�}�&�zT�g~��Re����āq�g��i�h�>�=j{=���1{�q���W�Z�9�h��iM�߰�7u,��;��N�0?I����Dc���&�������WWv�f����_ptXyt�`���"�M�ЫĽ�z�Β}
�+`�Aɀ.=Y��wr&�JWȫ��t�n!_��(��2��+����|�E���`�uU����~K��۲���'3�7Ţ.��u��Fv��닷V�S�U]T�QN>��Nt
����-"\$^�WS�è�B�0ұ�w���o0W���$A�DrWA����\��u�T�<�M*�l���O�:��\�ߩ �TI�ɇ�c���J����I�>h�&)�!gwbAo�Dk���Xm\�gbg3=o�[�}�qNN6�6�x:(��櫧�q	��w�WP����!��q�I�*���PE���B�,��CSF�Q� ��]u�&ĥ�A]o��?K�/p*	h=�e@l-V��(�Y�1~kƼ@7_�Rw"��%L%4.-j�=�h�n�Ec|�U/�Be�bI`�0��!�/�/�%3s֐��ߎŸ́�%^a�*{Vy�|�\/��_Bc�y�D�R a�M�y�������8?�!�uw����v�MQU�o�s��̛���<�3�|u�̽�$j9�zy	O�Q�)k�)~�oj#���â��f�T�x�!�YM�u���A1��R|�dq�O�f�F`[�n�����f	�I�L>ͣ'�%Nʸ��I���������_I���&4��ȝ#�W]��"�IӠ&�*�� �π����>9��|΁_�֏J���G8j��2[�u�CP-��t�B�K�|��C�v���+���t �3�mGb��#�Y�:��*	��+��ҡ�l&=���� �\�����K���C_ap��t9}J�dF�
�V��j��Ji�c�O� >m-c����K0~�ŕ�B}��
�"9�C\�!3��4����o�TН��"&	X���Q� Lוd�O��$*�-L�v��EpZ]�eri
p��:�|Ȃȥ�Su�XU|��L��
�tY79WYzK�,���S8�w)�R�_�Z��� a��sk�b�լ������q`y�St��V@ q�W���T��+���#�@EFqrW����1��?�K�G���qL��2�&�l��)`�(�&Z���% Ee���1�1��i�k��"��Z���V��q��s+���;�ZdsZC�R�k:.qrS��dB��Bj+��+Ѯ ��azִ�Z�x� �ϸf2sbX�ǷJ��*u%_Z&��<S��7P'�G�����{�M�s�8:�L}��-H��u+Ld� �4]��/�Fk�2���IZ��'���$?l�c��G��3e��s��lC��ed�9s��F�u�pzB����S�B!<�,S�եٓ��M,�M;�1e�;�vv;.9�@�#V�)�F�f�E��Yjy�M6Q�.�J���gi��L0ξ���q��G?#�{*sP���&b�h���p��,gSd��Ŏ�K+Z�vI��oBx �CD���N4��Ô#bh�r�H��ѩ�M[����/�z��3�l"J+𖵯�GΞ_����C{������YX�ܴ;���d�yJ�d{N+QR0+VoN���ۋ�����#u?���v]A¤su���\��J93���t�{�*}���Ʀj���/+�����������:��Z��(���p�19J�%A�ſV�t�~k<���썉�o�_%�a���٬��t� γr<��a����,h�G[��$
���:ǔ"u���-1�C���޹\�*u)%�fz1��\~ @*�G��v�w��� (�g+�'�ڃ��l�r�/�?>���>_���&d����>
��T�)vo��3��-��Ӫ��ے�vA��	�G8�X �:�مf�E�@����[���J3�v:��6=�ɪkp,zG
�MD��'�W�s����k�*ʒ܆�Ds���3���), ����@�Z��ǀ���������g��Stob�����{ֿ���[i��D�s^�Pޕ��P��~�Cg�z����������1$Q7��Q��R|p�K���������8��+�4�16�
-���v���~�s)ח/1���� �E^u��X�"�Q]^H���Dh����Z��`�	�}�)�UH�5}����c��G��K5��l`�P����DU���|o��d9jh9���~ �
�=��T��
�1�b	��Oȵ��UP-g ;Z|�c���9�⨊���[pq�{��&�{i�7�Н�˧�&;�y��T�kzh��@��>_0��[�af��L֜�$�Α����<��pMu���Iwc����p�'�c�����r��F�J6S �ş�����)x��e.�Ux-e�O���QK�Ŋ��P�/8m�`:a�@&��}O�14���bI귐�Eg[���W��N�/�۪��,�$Ɛ/�!��#��jسw}��ݳ?A�NM/G�x�[|2X���Z��'�	t4�ķEғp���|��H�}�\��[�ڲ��%��MEE���� ��F�/-��H{6�4rҲ�L�`��@�^�fUOFoe��xqC¾�Ƹ5���i5�(ݦ����m;���
�d zvfg�U�9!:I��[�"z�_a���E�R���X�`����/�;�2e�o��I�H�r�=���Qµ��7�,�}�>���s�����=.�]��<~���]$X�7��:�Q�"Ҕ���ҧ�(m���\Y��&O<Lϣy'T��Z��(GaD��$�������M�-m�e���^����+��l����-�b�wso�w�Ʒ5��@q�7$�\'J������4&�i��������JKI,7,Z�
���W��ϰ�lX!�&~9{��ѝSY,>��P�M�e|J�����������F<\�KC��D�ث�����
����5�r�-0��#�������#xi_J�rp1�EsZ,��zX�F��lA����G��I�''8-�a�΃���\����k��kv�j��or��N��ۚ�t\ۇ0"	S�*��OY� W(��rv�gB���a)��� ��h�;0�f��)�E�r�
�.��}Z*.a/
ߒ����z���h��v�"<����*.�Qg[-4��A�����l֊*�	נ�#���@:��yY�@�C�F�ì �6���>������L��s6�e�C��4
����zæৢ�I�|��0�{j�Ap�&���Y�h�v�g�������������[���h̩!'Oë_�p��k���������_��:s�����$@*��0F��蓌����i��"W��m�ZX LE��Jׂ�����V���5օfҎl V߂���%�﭅H�Ͻ��B�N����e���U
��GBYiC�bq}��$�O��u�����*J�D�SV4�"܎ϙ2�[T�Gh>�t�o�"�,�c�
���-'#1j�#y锭��2����W*<�OL'd=]�n�*5<e#HJl'P[�D��v�P��x�m��2��;m}��|v�����z�T��GLpU��3S�U׉g/
L镅�w7�����P~ѣ^e1-��Sg]��x�Xi�Y�d�" �Iz\;�e�V��ʄo���fP�H�􏻪V�H����g����}{=��5���ԟH>۲ۉ��:{.��ER�@b�'��sa;�7�2҂j%,M���5�Ei	Sк�5sj�,e8��G.O��;Z��o��dJ��Ř/�"B� ��J�A����b���U�������V#A��6�1����騞�HV�)L��V����cj/�Գu/" Dg���Z�\��2Ϲk��j�\D���>�#�oS�g�EyK{y������#C~ҿo�;�@]��~��9�8'`�J
�cd��[?[2�;�9��>�7���Չ�{4uܳ?�a3��TI�).�x"�\���B\����v��\��N�g�X/�GU0K��D\�!�}L�}�V))��"�yl�b�_VR=�i�1އ�F���~�iQr�K�I��������9hn淽bk��t�Q��U50��� ��:�Y�E�Q)�a�d����]}�"�G{�B^pG!_���X�+G٬���^01�=(�Y=��o�O4r�ٛ���B���!I���Bu�n5��W�M[А��!�"p�Վ�M�A ���a<e��B��8�UC)��
��W4X�)�+��!��@����y����bP7�H�0v�Z�\�P�� ������X�mW�Zn���`(}|f$*Ro:��?��Qj]B$Y����U�'h����*T� p�
Vpq5"���p98�
,!�H�eH��>�Y�؈X��@������c���K�; �e�I��{�8��ß�$3�j�؋��Ҵ^����7r�Ccw����!�H��Ǻ��e� ��3I5��S��4[�,��h��\��/`\{Kz����CՇ�ѥ��3�i�V���Q�n5�'d����g�F+�)�V�A�1�����&T�OR���օ�Y����p�F�+/&@dz��C%�D��0'_�1,tHq�G����P��9��{V���}JJ8W�� �_VI@�"(�)ź
|��0َ��V�D��#���B�")HG����u"�<�����(@g��Q���<������(������N�0���砧o��ov)S)O6�`k��X&Q�c�R-��r�� MK1gu+70���~eE4�zA�������Q���p��F@�0�{��NN��,tA~���@�,57·3��K[��_��}���DP{1���
&�m��_��w� y)��X������a2�dv�3�`מ�]y.+2�QJ�M�BW�^��.����]%�M|�MŊ�p�kS�~�B�a�|�fn�r�m��a� �^��{��-(Gvl7�̘��*��^<�	�~Aj 6���H��پ8��ծ���k!��YM/���K�ϟ`K�Ž�Ȓ'W;UwR�r:���|�Pv���=SM!��K�95{5|n����#��V�'�>���|���e������ku�"��\kԑ@�E����.u�ȧ\X��j�&�2rJ�e{5#��6��c��E3��
m�m� Ob�DQ�il��h#�1 �UwRE��>�ۊ���=�nwƢ^��o������q����� � V%a�ڔr����r��̄�h���P%~�!����N̈́�-X�š���I��$O5_Ug4����� n�Ǵ]0�:2�	X��l�؄��_�I�[�1��>��殖��P�\�an~��oJn�_?�M��?���1�)��Ƭ@�5�ie��WF�8�JX8k��B�t�]-��խ� wf�����AGi���3�Y��R� �eX�!�w �J��4ˆ��bE��n�gXtvO��Z9J�m�����Ҧӷݧ"�N��Ler�$"��s�	λz�z����Ѷ��Z��]8B:	&^U��-h��<Ā���J.�h�m<�2�e���	����:�`��-T� UƢ�쟱Z���d��r4�b�Їҗ�C���'� }�A�0�牭m����f��qLt�����[�xD��i�<�'Z`��Edch%e�.�ShH"��e5��%$��`q
"�O\�3���:��1��ۺ�?k��㿚hW�*A[� ��fW0�Z�t/Â�Z54o��n���Y%�C{j�e�ou��O��ˋ��9{���n�N�	� �G���0�����Y���4�%�xR�/�G"(]8�rf�j��[�<냝� �zB�N���#`�	7mʾhh$5�4�7ױs����o한ہGwF�}&c0@6V�ٴ��X�
���"�v%���7�"�$c4�ɢ��B����m&�HeP�or��Q
�$N%��;dn�$�S����I��#v�Z��ky"m�|۪Enf���ԭ`#��&^�~ߥe���~<ȴ1��P pJ�τ��ÆJ�h}7�s&-�AoH38�	� ���B��8�j��oIT��z�oO�A�iВ� �g���HYl;l(������S� ����j9�/c��\(N�+y@+��P(���[1d��o$���=�۱uT3�XUz�ώS�r���CϿ:!�X�6�ݲ?�e��7� ���؍�5�^�=pǏ��SПv�ؼB�I�~k�G��4�<#jD��'%��͊M���yr�ͅ������r�|/�:��Q�M��1��l�,lC#���t��\��;��"� dw,��@1x$/��~q��mB0�=*�v{��M<�i����P�7�V;�D*����a�|�[j}���0��|�B�\�F�-���,��$U���.0�Ǒ)
Mz��ʇ5����.�e�9g|�`A�%ݯ��R�Ìogu}^�Y-��nr��DY�W;���pљ�����2e��K��H=mN)�]>Ũ��b�4x��!��S�C&�C27�;] ܕR���o��&]q��$SZ�jլ�ͭ(��d�n��~�QI�4���2t��P�l����`�?�~���A�fu����mr�ƣ��*���}���f&��b�C�+b>�u3�E=]��w�ywuE�p���xeV7t�|ɜ�D�6�JAH�y~���n��VN�n�'�� ���|�C��G�.䵣:���/=�t�}:])�̅�R��6[��L+��GUIy��(�_��l�6�3&⪀?�H4f�`d-x�K����1�_�A+�)����J�f���U~���qj�j�PZ����(��̀Lt��];�?u�@��{b]�-u�����(^
�M�jǨ��b��b�A�. <"��W�H����,z�����%ڞ芖�k1U�{����^)��gM�hN�6K�H��lȤ�Ae��!�! NCM�L"�KV�V�����1>#�6�yTڂ�G��%s��@$,b,�zֈ��A�X���ݳ'��l�`��l��>�J�+�����jKϥ{^�V�A���� ��E��ۨD�g�]�3�����P�k����_�\��Kswt'O�yz���ԛ�[1��O��]B�E�Y�21�C��fq�L{��T$l��K,�b�ݠ5��/�>?���)_�ڼ�]�"�b[sV�a��&BV|��ؚ��DC������['�����G��z�8kŭ�aQcT\D?�V|a�����m�v �v�\�6]�;��������L�t
��[o��K��V���b��1x ���޶�9�ԉ������ժ&��c�m��y^\|��I����D�􀥿_�E���,�P�$K��B�v%.a�/vEB��d>���:j��XZ��=H�	��@L���C����`\��`�9u,Pk%T���B��`��w*6�opoŒs�ν���A���C���b|k^��y[�W].�m��"�O�b�7�����7��#<3QC�[7�K��ưΗx�Wt�j��#rCߋhm���=���9a�~p�.0:<?���E�C������������ [��{	�&��oY�d������}b`��Ҥ�˖&��Eܒӱ�}�ޞ �O���!]R��l�0��8�p����数���&0�{b��=A�МA��3�ců{��� �`���'��$��!�e�\�MK�G���v��g%���
�Ȟe�o�H�U�4KYc�uЕ�{	�z ��s�ڶr"�a�����Fm���Q�a���>1)��:.��<a)st_�����q�s�{�t:��� ���tOd@~�Ǝe9����������z2�@��8�~?�\���R��}���ߺ�|Ж������2@"B	�����ݴf�����U;�)���ͯ���`�2�����4�A*��ٙ�u�*�=*�{P]�)�"��R��	����q$�5*�����ok 6+O$�gH�M��J���R��⯿��L_��`w�eha��v�?��&#Ҙ�I�����7�7ti�ŗJO�dNh��`�OX��j�Goc��/D���o�}�SViNS�.���+�;[���e��)��f�/�2��ߑ�P�lE��
�=�3��bf��������[e�@ϛ(���y�{�vl����s�l�t��z%��)�V7;"R;��焕�|�@@Q����K�yQ��e����'�D6����	"��Z��Ф�r��2���آ!�s�C_k{���D>߫�Z�]�y��2v��fNP�12z9��y슉Dx%�u&��穝�3^��eΐ��W�Zz�b�+ h�����jp�`��
:����{�肰���舟dqy���װ��<x��O��?a{�������Oi:����g����KҞz8����'d�M�Q�>]�����a3f��9�#�*SnE�T-����'�^U|�3�E�'?(����}�����IN"b��h#��TNT�͎�WyfӴ�n�֚�%�����n}o����1(��\��t��X��w1�A�W��S���EO�=q�D#�l)/f�ƈ���"f]46��\�}$��'��J�6@��hs���0��E״81q���}�|����v���	��.����X��iL �����ud
�?��O�Z�فm�p`g�� �ۉX�Ms��)�i��$t���na��M\��h9�J��o��G����~�ῷL����{�!9˰ ��X\P�r���.a�|u�Vi��,3�[�\zyI,�hB�?uPO�\���!PdW_
��Pn9D@�.������-�Rg���Ϟ�	�0 �ù*[5~��󗰙�/��߮�_:'�����Ϊ�=f������$�|0���扄�uW�z�9
lێI�Ȇ��ss��;�����-BTi\�P���б�{�d�؅�#z��(X�!��%�͟0��� C���U�o��/k���k��/��� ��a��\o�S����a���w\�� �����G�"����C�wEA2�*oR314C!At)�R���.�4�&5�60;�,�_����wµ!\����^�VŞ"U��xɟlZ�y��
C0���v�b_:y��� d��"G�P�Q�|�Y91�!B�3�c����h$�b��&�L�Vû�~����"���j�ψn5�`��f8g��Lp9x?��㒗�8�������S��3�]�]�����G-���������:���-�̗�0-��C�i�/��X�咣i �`�O4z��.���7��۱���)7&dЁ��Q��ˁy�If`Aj�f��$��(�7��ݢi<GG�fqA��B0������[����h�
�23.UOX�.�4ڄ���n{��[W��S.ҤMq17��o64.������U=1���gas���{�!�1iV�HM��w�a1�%ט{.{R8�p�	\���-�|���'�A�SQ�~��O�r ��0�L�	���Q����0?���R�%�����" [��ڣ>���]~���-��L��
�d�^6���=7_��qxb�}I&[rVD�UA���g�2�Q�Z=:����Q���5}�m|��0��,^�䌍˓��3I���&���~���3��q�������ʛ&���(Z}1�����^-n�Q
O���&���U2�	�g#Wdp�8�SAD�щJ����"�e��^|z<~�>�1�\�M�\|l�_�L���Q��e>D���GZ}]�a{��V�*4{���}�sl74�����hk����2ڶ��(<�6�M��H����xoF�[�7�����%����9x$�8���ֆ��#.�(��}����M��98�ꚱA��>���?���}1���G��&`m]�z��Qt9�a��9�!�L�e�I�  hvo�AQ˦e͠K��T�'�_�����/:Ԫ�LQi���ˆ������o�B&¯+�6��N���AtƠ_R�䥫�*u��.�I�P�^�m��g�Cb�<J�J:�h������Ro"2�%�<,�(�_)�z��t�|��������pL�"c��Բ:qk�r� �>�Z�o��z��ˮ�Bp�R��a1k��������\�bhĳ�w�m���R���;�8�^�YVʅ-n�~�ћH\Ue6�⧦�{� *Q��_	��?�<�`�������'s\ا��y��e�T�n�Zhe����%���XKk�=wl(W���W��=�6u�����Bk��>3�&��!�NP�Z'#f�L�i�m�*33!Cz�(��46�P�yN��M7���3#��b�'Cu1��_\:��;<����@��� XK��L�I91�k�a��F�%����|��p���b%U� �U0�/螚ƾ�.�4�9߭��_����?z�Y��m�R)�^xu1�L -ݢ3�OHK�7�ܙ��Rs\d`V\��f7�-�w��Ԧ�ik��_k�ʾ�:wy*���2t�ū�T� �P[��@�������e��9�ц.]6��������J�P�ѣ��;1S���Æ���a�I�c�a����8�}�Ғ��k�Ub]~c�8Gj���T�i`���\�'�mS��_�!@�8'{H����	��U7!��/��b�lZ�U�!�T"~ H�|����mD��T��3�ͅ��`�?�@Ew;i%��a�v�����N/x!��o(��E�y�m�wy|�'=�x� - �����[Nb�Kn���v8���eׇjl�����a��E���mC.#�3[�4�	� �	�kV5�oEI��k	��y���ӭR�/+������5Y�b�
}al?���f��e�d!H-�,%q�	S�S������7(����z4 #�;0��{
��R�a��R�*�)P�x\/~����7Y8��O>�m��A���^��6��H�aS�p�Q$FF�d�?���)�B�'N�t|�����<�9�Um͝����k_��j�ҧjVW���h����۔�7��+��uFBk��rP�����1d�����K�ooi����Z������QSУ$��DK��"��,�T2;hO:�~��7J%2�s� ��2LuaAj�w���$�	zg�s��,��wgPY2q/r9��	�_��T�MI�')�M\� J�����`�x�����<i�E7V ��rIq�x�̈�#���-�0w�~)�kL1n�I�^&�YY3��Y��E��8:��{w��yҍ�6EW�x"\�;��>5ү�g�Q�O������"���Au7���F����Y��P�$�#�?�`��Ҳ��(6 �qUt��2^��&Gn�I�,�R�Mp������1����s�g�A(AT���\Xl�3���f���a�حL��[�_IkD�><���>]��{���}�b�@W�)��j. #��&H��1�u�'!�@�^r���e?��p����UZ���)5p��PJ����ef�Ixl��YU�,�'paj�b�0���{EM�ViI�anQ�hl��7"����& ���u�af*�y
M���#���d|����Y��2��O�Z�@w�'j�e�A'��iB�?o��0�C�Dkp-�GA�Ǜ�4w^1f�_� �Q��S�ۗ�����T�\��/�ᖖ`�	Y�U� -���5�d����*�!v9�-���"�C�5sf)\H]����_�3;��:ĥQ�Kza���ýҙl̜��Zg(�0R�Op�7�vv/��=n��I����8����˾���7t�Z7t�-����&�]��֋r�F�T�>����W�0����ڳq��Xj�i0����>ֹP8g���F��v����`��+�� �_���Ptm�%�E�ҁ���n=ij�F��k���������5�74�2V�}P�-���X��}4�& �UOd`'�Ԑ��2�h稷*(S�"[��Τ��Xfjlh�4Q<-F�}l��3y�i�L��.I�Ԧl�>%�Ov�WL�f�+�|/���|%��DD2%�cܔN�int�U	���9��	O�a�A�B��=�.�蘆o��'��%`�k|�Zp�l� s��39(�ĥc�
_�D�(��֒�U���������N �D�2�PH���	��43�[�>�ݲ4�*�qv�z�����	!�K�#��i�6��=q�r`�so�{�ڏ
���K;���x��� �����Si3�ۤds�H����͢�]{�q�Gy7���8�=��:��H�e��<I�78u5O�+�Z�΢)9�E��(�����]0����`Ua�cT9�#y�r�A�a&���'���!�!��0�i��j?�ߦ�?Gew���(�5��<��Į�!_�3{s_e*
0�bJ�k:��eu���T\bO:��Q@�*u	��C����K-Gr,&�֣�lF:�}�q�P�,#f
y�.E8r��`[Ȯ:`�Y�Z�z�P�"��6`YU����ԙQ)/.F��������[��D�>���^�k�Ii�;t�g���=��S�O�`������ t�5�&�EǮH%�J���]�&K��q��w9�NQ�dǩ;	��bN�V����0�n��uWD�ʓ��H�� 9S��'���(����4|]uJ�.�E�(�	��:�ʇO�Ƅ��XNz4���[OJI�]a\���X+�L��W:�h~3NT�&?}�/܏m�!Ҝ��!�>��ٮ.{�nN�)��.����΁���f�e�����T�k�4�� �ςǶi>ו��mQ�n�۱�T<ֲ��cg{v�M�gѓ�"�y�������ik6!��=	3쁤� E���p�;���&�2U�� �T����P�0��"�˃��Vx$/0���C!�礼�ޞ7����דrm|�5�p��#�6*����ߍjVu�%��ܥ��՟��j�%��¸�02H�0&Y���e����}��\5��[t���
g��U�p߁�ܤ�f{1�@S��Up6�1d����[�^pZ��{]�.&H'Sǳ�7�o���n)0B�;i�2�.�qI��GV�x`w���g���i���^[lzT���/�|������9Y�<�Nר>q�8�f�KʩU���$���!�H���*|A�X���R��߹B�U�n���A0?�3/}���oto%���v���˦V6r=N�V��!�_���	�a�%[1�;,M|*��{�IT������|Dp����
Sy⃪L�W����+����gH���XW?���_�C˩�p:��O��>˄ �,��X�{�I���V�v7}��qy��J�?W���t�J�����*�4,U]��K�ߺ�~u��fKo����~�!�˸3%�v6M5�׫� Jټ�d��@�_��s�#9~w�RϠZԭ!^>�x��^K �Q�MS���Wn���"�^��r6�'��fi�^��-}3�t���X�TT�t��c��$��8��a0B����i�Ȯ�C6՘՝q8k�3~q�k��8w��'�b1����	P~�n,��.���x��/�k(�ڒE3<�97ڈ����Kz�fN���jK�s�.f!5��x	��/5N.��Y_[s�h�}=��G_b͛�4���b%2lNﻼ������e��PA��:�G����:x�=���X�}�j��V�l��с�����*.:%J�'�:�TF���)���ND��P�����,�;�	�-T�D�ն�����_[R�6)XS�.\�4+v@t!7VCZ��v^�p��Y�~*���H�����y]�ak�Ql1�IDu��(��'>ٶ�*ϳU���k�;�=��@� �/>u{�G �1��vfU��!�6�Q�S�p�Wd��m6�9�?����*��=��8��=XUk		݂��@�L_'�s�_�\�*pmL�,k�1]�B�(?��m*!����F��c,���5�Ķ��?{`r����.c��H�	��b|���M����Z�j�	� #�A�S�^.� ��>�D�m����"���rޡQ�\�� ����Eȯ�C��4�v�Y��?hm{Qf�mk#])oʲ|:$��󼧣���x��J�)�e	�[Wsg�G��:b����:p�[`��{X�$햴rҞ�h崕Tt}Ґo���Oo�����`�t���~�H�%��\���y��A��76�A j�׺ ��Zy!�nf볔�-bg�38�ک�9��xi,��0�Zq/���!�a���!XN@�w�ۓ�]R��ڻ��עì�F�
�'����kR����� �ä�F�"�tl�O��,-�*�
���Ǚ�Q��L�@46�������Ř֎x��B9��W�֯��U���g7r�!�\��R����#d#��5�i�M�3�����r<s�������
s}^*8�	MUh���^@�����؋t�,���5�?��+ Q+��@�ͣ;�<�ծ;�+��Lﱴ9�2�4P;#,\o���p��ǩDE�0V��k=sd�4��D)h�1�yHl��4�5Ξ%��K��p� ���"������6��MǷ�_O$�w��<fk���d��x�ف��P�@-ju|��jڗ
Ya[y����A���U-'��k�'��]�$����Kg�:���|�.���;�8���:��}��T���/qR!���U��c�� �@����.(��yN����蠶�h1ړ� ܶ�H]� �t޽�R}�p���yf�x�C�y�����&!�'����n��i	�@�|r�������Q�����J�w�+����k$7�E�YƢ 9W3��H�G��O@T��L��%0���h^��)�Ro���#���g��㟯P]���u��=
��ق�H]]��6�=�O�@���k���i�7u����H��ܙ�7v�Y��0z��=�w��z�<�"S��o�1e��񁥲뚖
�%4~,o��~LFQ���j'ul�����&o>-�,� �SGHs�-�n�l{2GB>����A�,Z��:���|~Ip��e���R��|��i�Ss����?z�Ȳ��'���)������R�1��k:���oQܢ�T�)�Y ��Z�H�����`=G����e�=C�>��wW�F�yZ�:SuFuhg�����D?Bq�o8c4��4�k)���E�2㵚��LD�S�0j���L�O�X�"��U���T�Raf�gCgT�� ���IhZ>���0d)�J�f�i�d@�Ԑ�skF8�/��_Էƞ��Zw˸Q˟o��f_���&?q�r�OP�ه>믉�I`��z��EAl���m������r��}� ��)�ȱ@,U�8@�ER�P	��'���"������˥5{�˖:Jf��Iy�w!��4���B��je�.����iMǱc9�[Ƹ8ׂ��X��Ogr��2��Uܢ]<�RO�n�]Kn��G�����������!�<6�{��L��h�L�,=3ÂG������R��9��0��{�$#�W#���`��l<9���KW
E�X��d����|Pe�v��ڡI�i���컔���[$B<Pw;���wG�<w/�|��@.^����.���M�w�t�����by0+���N�I�@�Ѕc���мj����J���������u�Ƹ����I��W���x�ƴ����&�)��3��~��,Qc��AC� 31*���k�K����8�%����g����1�!��M
�M+�}[҈��F��0�I$���Q6>��),�6��w��^Y�G�t����f̐�� �p���� W����-�u�@��Z������z\c�ˇo��Y���mS� �ss�v�6�H��=Y���G�V�O�bݲh|1ܑ#.v�EL�
�^�P�E���:z�c�rrlX:���ƅ���n��0�x��!+C���L�4�݆""0wU�`�_��5�(�~��A�u��f��*%]��Yv���{�����8�l)���]�a:ž��d���=H�h���;��	�Nh�`jy��e�b��S������0�B38�@S~�n��+;��
I2�����utD�ȑe�_PC�)�I����I^ʏ|tu:(2{��:f'y%�he�4�*�t��I�M�Ş��s�Аʏ��hq��6�9��qq���xڸ��t�# �6��Rǈ�fp]�E��<�s(!��3Q^5	�}���k�.)7/���%�%DHf��Y�4��K|B8����~A7k&��lf]z`��[QAb=�η$u�<z��(ݦT����
FVx�1t�wV�xH��Y��l��b�_S�~�Q^)�^�����f3!�m^Q��#C#�JY"/��zFo�DC�T�ח~����hI���h4��H��Zι�z��̓�~��_��rjkB���4l�gmEé���LR^�.F����Xjp(��rW�؅S>d��&w���_��B"��Ҡ`�G̓ƺmE�Ƒ��}�"�8��z��=ӆ�R��L�[���p~x2q@� �K�@�y9��HʣS�	l#��V��<���K�������_}�3����8��	��e�%U��&R�;�%AP,^�'˙�y٨Ixǃ6���a�QS�o���Ȯ_b}���SUey���W�&L��z��UT z»X��P�8඿rlI���e��C#���m��G�V���!2�4MR�T�����^���I��M�7ݢs�T워GW$��"r.�A�����㟨��ٿ�^�)�O9G���W��2E�'DF[��p��?!%@����nN�0�ͬ���������t��-����= h�G��6�>��n�����*�4=9����ר�?$Zt2v}O��+]��[�O��ʥ��Z�v�_F9XH�]<�3��\������)�&S�zb5c{\b�Ìl(���-�����OLx��v��r^ե3�(�3�X{�mA7T��n�Q��8�H�B@�9�[��z9�M�n�Je���'1vB�w~�'����(�̔�vZ�Y:$&��f�(I�� �g3LE�w$���S���4HIZ������o�:����3]b?bS�m���r>�3 ��j�39�6;`	t{r�]CF�Hk��-g�e*��\��'p�)'��a�3� ݵ�gא+��a�P�nJ��c�}d��3�4�Le��3}]�a���:Ԯ�PD��SJ ��P���q��[L�MVt�gB�-F�ug��|�ԹkHk�U��N��~��>��74���R���3�I��1�'��>^���(�mg�|���k���O=����t/���;�g��t�)������a� '���ۭ�T~�>ց󦨦>$!�� _�?�N�G��?��\H�5!��+���]^�H�dw3MA��y %qҿ���ܯ���n,_�ik(џs~�+�=\$_�NpՕȼx�ܘ�tw�A>V��٬�`�ph����p�="�<��ֳJ?�>2��V�_B�����Pq�7�/up߱�g��A�>���ܒtOP c�#\���9L��#�T�Z���:��dRĲEa�r�w_�f�m^�_�f[��&.��K���� ����=2�����&dǅ��1*�N��B��sy ,�ȝ`��W�A:��mQ�U��o+D�����<���lKde�*��M,;@������@B����楜~Q;|���b�0�#Uf� F���B��vp&�p���d�qO�w}/0�+[SlHE�d8�q�9,s�+b!�a˘�Z{9kŨ��N;�q>Q�E�{y�h��:�я�@\Ľ,�<��ݘ�f��i�;��ƻ
�~��'⤄�H��u��[c��[ep�����\��ye��yOړ�O��ήGs��,�\e�Oy���d�����R �xyE�{�=n��*<6-�
�tGD��Q<QRU���+���g�O�R�"�ca��1rp�?���u�!\��2��w�� 'ߌ"4�H�#��q5߃�[��<!��#�[	��9��պ5ц2��qO�R��;v���>�^�^ _<�	��in��Sv���Z����?$��e�v�Ga%d�B�l>�X��;Ro�����:-Z���0�*�x
K�Rn�g��=
N)�J�M��E;�Q����#��D(Hn���~�ӨW[�v �͒��3PcM>�:�L���=I�gg�"O��F�<�iU�d h���H����$�ݣ�X�U�01�gS���̀�g���/D�}P1�̏z0�꤭���.-*�W��wn$<I�|V�6ԑ����	�13�3�v8�{�'�U��E _d����ӊ�~��i����V~/����@��L8�7�h�����zg������g�:R�����L#|�D+X��N��И��]:3�{�\��~�%:�;glAk�g~��Z ��e��)[`L�[0��Ʒj,�,�L��PG<�5fs��$��n-��h���i3��C�Oj{��;��Vqx�TTl<k  ���sU���L܃���&�[��$���6I����H�O:t�.�M9pT�AŠ��e��5N�s�~�� �����ʬ��;�Sz��s�;/��/��2A�t`㨙 Oq��'���G+�G"��S�
d��ı�`�[��ԑ�v�l��*�z9u�:�e����A��3"�h�_3���\�UVq;vib<݃�a�-ڗ!�9�j�摡 A�"����铣��|>�q�v�g����@���j����Wb���d����,����Gյ�cF6�cCn\��ǂ�%�>�-%��O�#�PrWG�|��K���A�a��Ӂ���Ë�w6P\_�w�<nK6�
�[.٨�١0�:
�U�j2ɔk��]����	j}�I�C5�O�}������.�	1���
�DDD�h��ե{����C.K�=yŻ���3l�>ਢk��Y�����B��'�����A�zr9=QT(؃~%+8X�m[?�3xk�~��^�E���k�K������lu�����P2nM1�����w��;�#�>�Ob��)�C��(��rU�R��	i��zF��|�E�y�x��e��;��&g��=���3~�?|]��������ܾ�-q��щk4��1P�v�\�*�A���G�_E+�\�����Du,�@�F@�A�%bL0�4MJ�%m�-�N>]q��c.ܧ�s�ᬚ�~�*� 氉� �S���q$����S���H�ƅ�Yf���e/K�t�8�M��<�'��������|����A�Q�D�[�$�|���C�)�#ZX��j9�l�[��U�8�<'Aŋ���Iﺙ������@W��ݓ���Z�iy\�{�5<�N���	 �T ο��� ��J7� nT�K�M����o���2k�Н�H���!Z�/:�f� L�>��9����CP��@Ŏ�*ؗ��/o�������k�G|;n�O�����އ"R&:|�����������M��l(�P�t�_���^y�\� �:|��2�t���"�����A����]\���Y��Y��{���<�C�T�ϕ��G%yʊi�E��WE^Q���j��ѡi��&u�9���)�)�u3\Ag�)y��g�`"���8�qsTF�NLIr�O�q�E�"V�,K�W���cj�J�5�c�{T$	�������P���Kˆ]��l��W�{�ϐ7O�NY���9u���xv�"Z��Δ���FU�us��ow��,���ɦRL��lf l.^��o5ph���'?yG�%�Ջ7�%�֥]�P��R�Ps1i�U1�PY�K�m�h���A�����m��$�k��^r��qB)��gU�+��#�jEf�ԙn�0��hV3�O���N��'���.����sˮ�+������1���|F+����m[i�iz�r˼/=M�X"hd/�^>�Ԙq�)$��(phm���<��RD���g��nq��ҡ��e
$Z�%��<fG�?ש���xe�����|�D������Or��G���D���Q{���5�\��gb��7�0V��_vvzx�9|����K�G��O��>��q�=H��bg--� rp�Âܼ-�/1��n^ۣ�J*"���]t#ύz��e���S-J�r�/���U���sw��i*�q��
W3�`�d�$ٯ��ԕ_|*'�3]��xd/R����
T�U����PM�nJ�4�m�
���������5��X�Y�<�e5`���t��E�^Y��cE���	�]���U0;����X�V����)�55���	",��o�lQ��qdFh���fꛡ�7�1��`�2�U�������Ts�XYW����c����b�B.X�C]��h
[����I{�y��l?��-}愃|�n+�q��y��\}��.���]ɹ�]�(C+s�t�L���z�
|�W����x�	����i\�Bh���OM�.��\�`�n?�p�l�����ǫ.'l��u0+�v�������FI=� �Zuj�G��h��z�KN�T��]C��p���|���\
�\b`�L)��������R���I�?��G&�FP�(��D|�5���]x��0�,��o�R�܂�?�9���v�>GA*ڵKm��>a�}�;�@�,L򧙽�*֚�9����b�S-���&�?�h%eFx��@l��sOS��S��-�7r/^�/+�Q�*�]_E��3m����r@���!���1�C9�_y�	+����� C
�o�h���݊tb]#r�#�9ע��q�S��+�Y�:�Aj�2?��Ģ>aS�`�q�M�q������o��m��];�_�Xr������2>8�����EU�a┷��x�#�����l���P>Pҡ�N�3����#��tl�wf]���)����m��	���L�5�i��n�{�����g,P%fI+:%�9t���J��
�_����� 6	9�x(������2e��I��6V3��?����`��8��.���Z3�9��b�Ez���%)T���l�Q��I�� U4M���:�g��<�fњ�ºi��/R�� 2�t��z�{�6�E���BAӶ���`���9���Zw�j����*6�7Ytc�G�oe\�Oj���r'�~{Æ��M�nΧ�? +G��?:f�i�b}�E����(<dtPZ~/ۥ��=��U�p$�'��@�_J��nͤ'78Z0~����ǃf���Q(�ֽ���>�ae�=CEJ�=����	R�e\����8�۵Ȅ�T%f3��pDI�����8�#,���~ \.�xvi���{�k�&�,��Zw�᧎@�+�@G�}Y{�/X��]�'gVta�b�=fO�v�z�Y�-Ӥ��|5Ѯ>C*@F:J߻��GW�:�����'��zA��搇�İa��7��Գ��������n�׫i��L v	�?o��%[�.�N�p^MUAב}-c(2�������z/Z����}F��r0�u�����a�"B��� ��L��7��$�����f�D"�r�]O�C�s�u�Ś����os29������ޭ�Ѿ��x��uBmt{�M��ByQ��,������Ɵ�J�e�Fl�m|��O�潛�P��ٙ��mG{�s�|�m�ڞ�a%p��P�����?*��8lU�ˋ ��s�G(p<���1��Q�=e/������~�X<��nQ�?Kl���M�.�v��A�y�&�;\�Ίa&�����1�&.�#K{e�h�ߞ:p���񔔸�D�L�V�'ʸW���8�ֳ��LS��
�Bu��J��@��9Y�s�zM�T��ٜ�� OH����H}��{o�fW"ӈy�H"��^r[F>t�n�=�Ͽ3�צ�o9Sd�Z6�U*���Yx~����ڤ���H��"�����4.�V�6,*�;Mf�"{V�{�$柙$ث_N�ϰ���Öp�|��ҝ��!�N���`䘩B�;$޿!�X�}ϩ՗{���ا��O&U�yc���=|�z�$/��jL�A���ٞ�$h_���ԫxf?o�g��J��}�?i�ۅ�i�̥/��6�3��aw�h��rє�h�;Qo���hԊ	���wN[jUzI����
�w]����can2Z������������*|��|r�D/N�}�`�'��:��͚Z���L��z�Ƕg�3���egP�`��'�Y�fm�h��e7�����/�@�u5��>�(���sxRK�X�e;�|Z�/�2ez0s���z�C�e�#�K1IF�4��W���ә�oT�͔~�2d�m�r����j�Ani�N���gk�J^�P�A���Ç�W���E�rUE���Qŀa��JWd��q�pj9~�v7��Y�$�9|R^i{XP�L���ʷ�q����?���0�H)n�%@.�	��p�w/� V$c��A:����uR�uM�z�e��:	�>=�m)�Ǥ��ϓ�K����i�7�
c
�3*f�"�db����
��ԭ�zԊڜ����z)�"%�b���X??�v��kt\��f��!xy~��?�	�@�7��F��i�}�h���P���6f;k�pZ��O����;_\^J��Fc%���;&�U8�"�-��poO�\������g�u���*���$[������j&�{ݗ)ր�:�%Ӵc�����b@7��*�X��ȅQ�m��`L��ZO���#E#�
�[Һ7�EZ��]��ױ�s"��)�r_�������*֍��/�ʯ� t9s$-|��k����2g��5v�ұ݊���{�n|�jͪ�H��fxVY�"�,��z0�&+�m:}�̽��]�������� �����F��
�-Cz�|���o��B0������'b�?����@�n"d�Z�l}��v �J��52�j�l���d��a�9TiЁ
AHA!
��s��'���w�ل�%g�c�a�����S��|5[�~��X.{�Ru�G;a��/^�����5Sl-��M�zUz.�����5=^��+.Խ��wu7�ep�^{Daԛ���T��W�o�ݻ"�[$�_��c��h��8�-�D����^�Ҡ�]���S��-���U=��-w̮�����<
����%�o�X���t��p��,�)ŧ��z-��� �P�V[�݃>Rg�/2�
I�:��;�4�3�B�a�H
lGfd�'No�?��TQw^x;�L�����W0�u%���^`WB�J���
��	"*K)���"	�^䘂`@p��Q�%<�˜܇8ͷ��-NW�#�s�N���g��Je=�-�b����ֵ)�	�R��, j�{¿	{3��c"ž��	�߈=�_[j��_�?�,H���cz�]ܳ�g�<hn��R�Ão?��w]����'Zۥ����0G��!V��[(�,m�c�0LU��H��]���� f8J�������%c�g�R8O�h$���~{��^�b��c�`�LV{*�C����� L�m����X}�1�qo�����s� D�r�WWx���]ǷcWx����l�z����&��"�������=O�`	%�惇�hG��z��A���xc�LgF�ʂ��.��R1�|PvőNz.QڍGn�����1��hi� ���O�e�S@�+��>\��I:�۽?Qizs�sr��8��`W@�3���B�Ҽ� �;� J�5Kȁ�����3T}��Rm����߼^߬/^SɃ����pZ$'�k|Ϸ��ҁ��M�ƥӛ�60��A�^6���~�A���l�^����n�(��./�,�-����>7�?Q�|A��)Al��h(���"t5��B��G d��B����WwH���y�/Τ�D�� �$��8��[4t��7K����m0�ƫ��N #5�%Vk�C��ov.�ֻ���i��㯁��L݀4���U=�C���5gq��P���"���^0�v��z�F�kA� K�zk��Ug�l�j����Fh����-�*f�����W��ȉoyL�l%�<N��K��$���X5=�NMnǽj�Ja����_�h� 1��q���+'1E��d�m`��pĩ\��%�@1;<�1��Y�����GOSS=CB�A"C�x���Z�����5 d����C7C�0���/�_�E����37��C���B݌�D,A���t���Gq耤�O�
48>#C��kM=x�	:pԂ�A2�z��y�3�0���A9�N��DS/4��=S4���܏z�~tz-͵O�wpY?V����h]��������|���?�-"��K�q�Z����&�A�%�b2�ݎ��"������
A�C#��fPtѳ����ԥ�ɦ3#U�3#�B����'��Ԡlw*Nhs%v���3C�)�N8�g�=��
��H��t��k��s�L
0����4�9���TB@ ���h(��ːс����?xހܭ��^��3=�41	����w��2b^�N�Jڙ(�i�
�G�Z!���K3u�Y�V��Mܽ
�l?�l��KB4�y�O���J�<�{KN�d�)x!���^���ԏ#%���'C~�I���%���af'Rl_iy�-�v�lsbG�@C��g��e�T�5�fR���AD����B&-d� Ɔt�[�;��|pV�1J��\��B�����tǤ����)�,��I��G̎v2e��`
�5��M摎/���^i-�����߾�d8D�[��y�"��!�Y�B��{�OZ��c~��"� fD�M���C;A�]!�H�����K�jX��Y7,��'�X��Ŭ�Fk��V�O˗c��X'����/�8��X&x���В�S	��D�s
4���%�k"�ڙ�Ւ�'��W\���-�'��Ap�n+rh돁H.�⺂�kNI��m�r�	ߪRu��qЋ�A+4tgt&s9 9�͚�{���O�o˰�����g�AO@YSsf5��O����ޢ+��Z�H�Zu����B�J�#���X��ө�89w���R��G�7���%���d�������޸�O�7��J�bd��$��CJ/��$c��G��[���	>���Wgv#��Z�Q';���e��"M�yCs�""���Zɀ���tZ,���7��N��F�G�untm,-B0׉���T��Ԛ�NBqŏ4@��Nս�qkh'���9��	�_q}�K3��>�XOG�3�'��1NVC�M��e�m�t�g0�h-����R���Z,GӼ��Q�M)MM9���c0�q����+�cC���X���mE������t�f�0�C�&���{7���	c�c�3q���$�,�z�>�r��Dy��
bv�:Z��iȀpJN*rd���p�b�l;)�F���M}�Fy>��R	7O����a:����H9߄�m�(�v9��"��a�cy2yՒR�=	��xR?A�
�W��zY�~.�jy�\��-6���;���h�r���r �X,~Ёi��G"�6ꊿ�W-
,�����Z��e�\���k��Q���f'��n��C�<iޠ�I��*
���.�6�9gSf�wW�~��{�)�=�e�wP���ty��w(�eB��P���Z��g-���'�Ԛ�5vQ�q����NG�oU��qZocz
��_� k��X��|�YP�����`�m9tG�g���~}��Zv��~��\�t