��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�����ręʔF�����^ǹ�*l)�tf.�<i�(t��@>S�7�Kۺ~�۪�����x|����^G�M��^���G�#t'�V��w�YP��J[���+�J[�K�4���UQ<E�ET�u�:GʛK*߷vt��ܪ���$���wՊ�`C���`����Lt�kY�:��b��O��vX�0�O�[8�ң�l/��J�d���*�#>I�|�PR5�z�+���Q��"/�޵9�������	���hX/15Em��N7�S�����v]�&����f@�_�!�8�􊠖�'>Φ��U�_�>Xq/}ř{r�>���R���e�δ�����t�`)�D�e�f�o���x2�&�i��띞�E;}^�l!IA?"
M���G�LN�ߩ����(��`��a,��d_6X��#c�����dI{�:��I���GA��1!o֧:o!~a�?���D��L�*�Fmei��h�e'cf�GN�a8\,8�r����"KuZe�&�l�M��HЃ��>̖��>���{���E��WqY��[���K����u�u�A����`sY>��� ؆k���0�ۉ��Ӻ
���~=�m��v+����b#k'�S�:P}��hx��4�سp�ߛ		@kv�~��ݗ�lݓ4r�uZ���;#}!�k��wQ��QN���x�T(���R�Ve6"ix$<��U������#&��)�j&���`ebE��Lr�	e�dB({ޕ��<�O����W�"n��h���1}[���ojU0-��w��Qr�B��-9���*��{����;�D �及�߹��6�ͩ�_) �˽
���|�񡀺y�$����n�n�?�<�$�	mw9��)}*R���LО�^R�R�>��l$����/d��)���`B��Q��E[�9�:�(+���;�SG��3L�-v�b�h�̀";�nWf�04����ZGQ��/n0"X��^~Q|�F�r��l|�Of���59��4vr5E(S�7�1�e�")0�*,Ў�(��+p�:=C�r1��Px��_F7�l~Zݝb��k�S�T�'�J��B	��}���A*�qOT�Y���D�B� bքop;���`�'�+�L+�O��M�r�Ϧ�NJd�	?z*V;J�>�7�c�ռ�QcY2��l�E��圝������ӧ�n�Y��0�M_�Wu�*w��}��<��P��"Rr���4Ɯ�B����|5l�H���K��V���1l�n)��{�;����O�<��~{�\�n��g twvN���zN�<0c���<N���&�e���kO��"|W��h��j�i?��h~*�-,4;��$d�[�(�{��
kHP��b[��LR���5~��ӳ�Q��we���VX��w	/� �a���.W��A�<𳶩/����������`k�f{�us�5�q�	�
Ճu�,�{����f���3���/��`)�:&D��^8�&h7���B�����o�	l�MGXY�D��as椟)�*�	H'\\]�_�>xk�����屠A?kC	��<eC$ ���J`̆�oC�"qP�mlP�W��d'D񨏠����v����x��f�I������]��9[ڼ����>�TH�~�̘�;�18�E?q�cXG�t[Ǫ���]7X𓸆tM���һ\�& Ƿ�U���d��׸�4���}.~�����a����9��/��9�i�ҺE�ݐge���NIb�yo�w��ҳ0�~С�������h�=��i�V .ܓp��-��Yh�A�����3��z`��s�*�d1�}�,ݯ��4�>���`k���r��O�KU[H ��n6�<�ve�e/�^�q���i��Z�U�1�ɖK>p$u��DQ��{��B��u|�k:���{�0b��7?�k�	@ ��$�[@���&�� E��	�����[�J�RO��q'�w����Nh�;8Ğ���%k��(����o�L̒d|���:���C�>z��Pc�>( N���A�e�#z���<�3BU�Eؼ9$ᱬH=�$�~������ʺ���Gʫ���*y��)��I��q0o5v�=e��Z.q[*ZԆ��3d�޶���0L/�g" u��ZȲ�;HJ@��Ѓ�F�b�^�#8�tk"=r>%8��-�>d�\H�k1lb]�(д4�LR4�9�g;:�~���-Î���K$��$�%���;�;��#S����9�	K߄�R��B��?��ƺ��p�?R����X	^R
��D�I�1̂��PLO~�
+�%��c������K�v�����h�zWm�NW^����yF �$�$�4���'�XI	�]��a���&���Qx*����z�MG�U�-w���b���E?ln�[��:��z�!��nPr����r�.�'H/� ���#�Lp4���#���/++*��mc� ��+���Y�GGk΋��u�(EϿ�U)ϳ��e�gA�G�Ҷt���������i�K^��Жv�?�$����;��VO�X�x���?!#��u�~�r�3���(�%�a��M��b��?�*-�\���@��]���> '����S���k�ָT�9�柤�w�e�I%�j S�"yq,s넶l	��1ru�H'�g��h�O�Z)�}U�1�����2%0�~%���g'��.����ǒ�v$h������d`�yԈF�_%$8�}�;.A�"T|�(�\Pz���*�bCH+�D�*�G�¡�d�b�p��FU6�	]�_4����4Q..[�+�ac�ի��
?-�ޡ&q�O�����1�/��Q3�$["6JB:�9� �5Ȅ�Qٿ���ix���ߏ�a�����(̬yx�l	��@O�K��ep!z�*l���Q��"d[����C��q����z��*�д��RΗ&jG�Nw���/��qZj��=]e���^Z.E�b3c	L/,b�Z �����;����%�O���wX�9L^2r�����6ys据�Jz�''e�o����S�XpQ��,q��R��L��k�i&$�`�׭����ԅK��ϫ��b<�A�|��>}�ڄ*T	�d��κ5���H�w6Fh��BL��L&#U�z0���h�����+)�?6t2��<�xI]�`�I~����ɟ�l,է��3�^�:oɋȄj�=?C�E��6���L��)>�d�G��bs��D&~2QS�T���c�Wi��spV��3��tw�3�[ʹ��4>^,�y�0�a'V\I�͗����"_"�W-4�}I�z�ybm���M߹��c|�n�:��y��P'u�N.��6B�.'��w�4��~�?Օp����@1��ք;���ؚ�����`���r�؄A� k@�C� ꇈ�b��n�_�G�'{	c�v1�W��wF%�%T�եS0����%OU�*/6`�����I��$�TM���RCR%�M>��-�!#O��:�k	p%�:�)4����GG���w��7�nf�Q��&n��E�*1lw|¤MU$M#4�Fow����
NFq~w;=7F�]�殹hU0J�?���� qk}%��:N�c�t�θ��.g�i��D��HVᘒ�xz��.�֯6�m��e�F�i��?�0�)��p`3&�p|7�#N紱��a�������&\5�������~��v�̇I�Q����N�� ��=?��K���� ����Y^��~@�J�}��QH8�lP@*��y�Dzxū��`�L�S�țO����`�]�eNVI�7�l	���# q,��t/K�K\�0D)$}\�UC%^d=�����{9����t�Fr����;�<��Ĵ���%�����M%���p��Rg)*��J��#- E�W�h���N>��+'��m&v���>�8��\��!0���T�U3�J�c��^$���O�.91M
�O�=��֊-���6�a�TL��#�w��}U�0"7Q*e�g~�m�DaR��3�5��˃o���iIt���JL���De����g��V��`�TzN�Qs�!���AX�JX�Z��a	��5&"�����|�_��?�{$����W��p.�f�]�z<M@�E⩀��~eH�}�M�5L�ڻ��Q�[���S��a����j蜄��(��}pK�c�0�Q5�+3\��배t$�qjg��FL"A�����V͂`����x�q<@��ݴ��%� �M��%<�D���r߫DR�fo��lkJ�ä;]�������f�B��~N�?,wh���$�ٳb��8.@�|,��sE1E�
��.�t/�|�`Q�Ϫkz��}/F]S�ʺIX�5��a�>� i��s���י^qK�K7bz�e���a���՚�|��l�� 8_ьϯ�G��P3�n��S[3q�^�^�u`���9�EO�؜4��{H�}� 2�� ���h|]����V����
���z��Cx.�=]��
��6a�%��t9u�B���ME;m����}^`u7�v��*�u�	.�v�$Ev9
��{���w����ղP����4�p���ΌFj�dQ��ef�c�׊V_��mh�&�h����ψ� @����̍tu�̨�|�3
�گGQE�B��������IfU���/f��#I�I�b���>�'�Q��T>,o�컐X�����2������C�ɘ���������,g��{�A�b�z~Dk���$�t���Ҏ��A��Q��xi�#�հ���xa��8�8�<i�Է2S�-���HX�x!��4��(x��[ޘ����D�v�*��l_vC^�(8A&bu�gooYWW���c���Akt¨)j[��k�����_=�k2	��:��]~�o�	�'>O�9P��˚u)'\\em�07�'�y�sz�����T�,`�������/�ߢI��}_�.*� ��3[�8�_����I��p92:����<���El@�B�=
�	a���3a��$/�|"nԿ2��T�p��z���=Q�+��H������hn�w�owwU�� BE�oM��u�w��fy��P��N��-�ʊ̜����f����2ۗ!���x*��f���]X3��x�y� p(�]��P����Y�0���E���H �8��3���d^��s�u���w�dH(��Ǉ�p� ��l^�g/X6@@�&�����j�dk
g��.H�*��� +f���w�����$�d��5W��*�<�o$.0_�[m�H���J�)�Iܶm�_a}`c���E�,�[�z��r"�ƚu�2EgK�:� ��A�Y�O;b���\h+��J���Ǹn]���1�o?j�(j�z���<�)�(�{�B^��I�=�XTG����ύ�LG (�h;��z�\����ur~9�Ȱ���Z� 4���m��=9)p�*�m]���j9xC�h��­@�,���vU'����>Mf���@ɵ? i�
�o9Z]@Đ�q�S/B�tZ��,�X�����pF�ą߂R��[��K�8�Nq��3��*)� ,q�RZuf5��~v+F�R� ���Xx1?�g�ҵfXz<��qi��Ml���G�����m۟~·	7�:`��1��Vs�Y���_\���6Y�ǁ�xG�d���\�[>ǚ�Qwl��hiL6���j�+��1�-��fx��F���**�u`Yدe��R3����m8�K����S[�}ycӃN�R����P�m�iZ���w����Wȗ�� �[�j�Ro PqL�{.m�l��r��A)�{�p�9P'�}�t�u����֛��E�$jO�����n�9&��B'��hT���c*�m6�(�9���2D���P�ͧu�yr��%�[�n�È�uu�t}@�/Qu��_3�;����a;V8<�ˑJlEÝqvk�b��H�T>����K��"p���
�y\�SN4N��(D�t��!��kM"ط2Iɖ�2�/D�3���5�+�H�D����:g
4Ԇ%n,��"B��ؐ�[6��*;��n����*_�E�,�1W$|��N�1nU��`��_���O���<���Q�~NT�p:�$���X{n��A�QՏQfT�W��g\Q��f��)#/pilXB���̂����4)�ᑈve�v�>��&&

'15Vd����g�Ɵ�v's�`������	D�7��"� #�@���*��@�16@2�ɟ�tЎc��E�;Ji�N��OO⯠�1�7i��.���[=�Z��'j�GJ�"�����Qub�����������]���Jg��R���;��ȵwǠP����|U;L�D�Z$�:�;�!{�	�<|�S.��_V���j!�Z�.i|�E��!�fN�lN��I�4n5��,�`2��n�U�!��*7f��ƽ>�mw�B ��fQ�Goa�9S*V@o�|����d�7múU��c��Ϥk�+�nͣ���S�摄�gO�}�5x��N��|��q�WR[���){]� e�!k��z(��	]*z�8q%c]P'O�7j^B�8U1~k����̡��$O��+��^��3�����%Q5��=��S�]!)��Ś5�$�gA���z��.�?�r�(O�����	F�2��V ��i�����'"�����fD�; Ɲi��CCYB�k�4gr�8�����#���N%����\���$�+"���nW�i��t��Q����� c��xˆ�Ci#_C�'W!��K������a��P���&��#�[�-�+��|����X a�����īmf�$�YS�K�