��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	���ʂH�__�>g�{fԛ��
`�[A��Q��/43r�� �K4��<��{u*�b������� �^��F�?)�ˮy5�H���<Y�"u��Cg��/z'��������(�pr��aI�b%l�!�[ߣI�`k�{�-m�T�`����d�uf�g%gӹ����TX;���9zeOǁ���	��X���<7x��+	�Q�����?���$��vr���H$`k*�^n]��)���4�N�}<D����2~�\��U�Z�Y����HG �7E��$H�뽛�8�T��܋�B���V%@$QՕ���G�l��l�k�]�f�M�5�M�p�����8Y4)�lK"��"\�ۘb�[��"iǮ���\!
��K=ɗ��S��0�^��p��q�i�f3u�.�t4��[����%ٽsR*e�i'�y����
r���0�7d�|�w��UC]b��{�rt�0@�~��5�^_H���6����_X��9*���5��`i�`��;���c�҂��id���t$�FHCl<���Q.�P�$����Wܗ��y h�+`W�Ȕ��y��!8�l���EH=�l�_s��7(�R���;}^� ��A���I�&��?�x��WR�X%%�K�
�F𣘓�(>nf&o4��֒%����k�JSv��f�tb�.�@u��l�J(5��y%��w�R���YS?��tY��Ƨ�ֵ�S`� �����)�fd֮P�]���E�Z�Ɵ���Y��u>D��U���}#RwT�"&�/d�?�pV}u��[�qF�����p�u��l'�2'h.��\TG���8<���Ε���H��#&<���L/�	���-��}���Ł@�#������ڗ��r��<[��J�u
u�-?$e)V��X!Qg`\3�T�ί��`�U�ӾEu_��.��@A�1�֎�z���~��Q�k�xq��l�Xf�ݖ�>�P����.-ui%����iN,Y��A*��b�IuK�T젌��v�����x����y8Z���H�%0�~��F=r��h�WԄK�H���鵍�p�$�����I�-��}�c{��M�K��=<�G����m�%�86:(��ˡ��F{�\�֌M�p���
+�����އ�=���Hw��7��L����ۏm�V��*�D��0���p�����6B#W�\-��h�Z�"L����t�
N�^��Otnxfՙ����4p5�P� u�%(Rl��P<���O"�nβn��b�eCz{(<9od�L���S��{�B&�M8�6"0�cӌ�� ��lrɈ,�"KT\�(o��ܜ�K�wO�6�	�P�"R"��b����a����s��cj�j7�je*�tsvj\)����x,�g�����,�7��7z�����a��$���p��~�`�Y�3�����N��L�Ól4qXg�=a�!�t$7�p���Wĩd������;f���S��������Jٔ�/��M�Js9y*#_*^�>jʷ�ʣl��S���d���������[2xz�<`���O��D$+`�Ȩ�C�M�| A��C�%�q 9��/՚�gI��4G�θف���+,"�f��Xc��Yw���1���K��!� I+�g��wi�$Who;�"J*���N�	�*w+�~�s�;Y�k��&�Ak������%1(	�u��]�Y�fgː*��݈i(��(��:��G��$p�6�8$I�wyM�fu�Sp�\g텦�G������|@5/p��şuw�K��(��:��|V������9��y�T��:S(��D"Y¬_�p?�K5�]�U��˶�*��@�8�i��wc�$�h���Z]�����Sd��}�AtU��B�����wy����IG�t%���\#z��;Q�U�=��8�"��u���R������7[�����Y���"p��P����Q�7��+��R�3
�~#�pg'�!%��X�R���8P��H�5�w �C�Y��xga�4 �@���.�T�cJb^_T9:� ��p�_���y�ݓ���]�c���;v<��'f�Rl)�
21�e:�P�|�k�"��QO���jCl��/l���z;��G��&I8
(]n����*n���ۍ ���)Oo��?ƴI
�`v>��6 Q��0�:d0�ɷ�B�����e��U�5��7;05��]2��<�/�K$����
�L`�=<�?5���X�	��A���K��|cd�l���wBȓd�
�IpNPV�E�~�M�[TZtܧg���>���xT��> �]} \���DF����OڥKed/x]O�̂c$Xp�~<�pQ%=��%�|�;)3�p�<�u��-�{��`��YN�UC��J���Q�?i,M<2�˞���;R ���B���t��g��q��b�Q7�������9�y	CdA�5��U��Fg^���ŭ
LR�BL�����y�y��$B=\���_8v�K־���?��4�{|0OB�SF��ܫ�[c���2sN�.L`�"i��$�6�=���g�:d:a~���D�k�4ub��x��i"z�}QQ��j��nǍɦ<цq�X���pi�:"2����Yb��D�7�u' ������S#��8S^�~��%@ ��([�
��P���<&�Rj�c��/����?�O2�fom℧H�X�����O�kS�S��������ř�ĸ1��/�T�Q��3=x=_����=�]Ltvd�Q��W XL7�3F�' ��W?�b���"��Z�g�]9 vt{��SH�EX�=�#w7h"��ͻ�ϑ���m���t��K� �ʎ3u��'��9aY��\�Ch��{�[��f��{��
��
�\���qf����Ho�!+�+�Q�� L6�,iAl��s�%�R�J:<��П)��X�G y���㮻�~��r�$��-EbJ��w��G;X{��G�t�q�è~�G��ҧ fL��ku�g�$T����7�[�^���n���@�x�>@����吋��}�C'�rs���Y\�C��[IIX��+�[3���H����M����g��r3SH	·�6�!�(�����]�%P�q*b�j�1�M�pH��|g�L�/��/��a�ɟ�q�%Qc��ً����Y�_��9��wEow��Qd�:ɂ�euGg�(���^Wŀ���(�� 4Y��.,+,�g�8���l�y��]q}��8Y���	�h��S2�Ae�ڎ�U
Z���c����%F��=��A��ޅ��u|���B��8�N0F���Kn��r��y�O8��~��0�[`�/oZ���>��4�+ʇv��Vv=�G>��&�^�I��8dʹ0��tC���R�0*�s��^B�Nr�����/^t�:���cXXI�rL�*���s0� �
�	V("q�h)�T��a+�m{D�K��ʰP-.]9�:e��gBL��g��C��"��t���$_ ��Y��$���&�p��ʇ�d.���<ˤ��}(�7�_z����V����U\��5�H�/�I�"M�[�K2�'.Za�m�M,.k���2��c����P�����\��R��M�� ��ʚɚ(_�2�Ǚ|;f�.�vb���_���i����E�D-3��O]�� I��r�!c��,�W��kLE�W�Y��[�SƆ���Mc�����y�XKJ@�:����K�u%�KB�P�P�+��Lz��)�O���|���FĐ>�YY "q>׸i��1��7����8�x3@*���=JA���V�%��H̡E�p'������;�l����i|!>�Ӕql  ���-v��;�-�q��=�C��7��r�RB�BR�v>���8�G�, �� "Y��b}������1�E��8�?Qb�^�fS�y����L����/��G�P�V��%��>	%�yN=��6�z��#���w{,Σ~>7���Uы[_*�_�j�ךwT��h[R##j^�S�3G�1ށh8W�r� L= �a�wZS�Z �b+t֢��?ڡ	�^��+"3 ����9�����Pzo�|Q���p*�,_�s��)�*��(�E�L")fI�瞇qj�{�7�RR����]�w�L���!��)"p��:�&I����M S/�^��~Xf<��'���s�O�M(�;�z�V�+-�p���c^�yРP���5?afKC��WoX��1.�h�SFᜏ�p�a�π=x&�8�
���-����5�Z�����ɬ#],:F��l��
ָD#�O�
�����p�qR �	6� rPq�=��r�?��<N� �}\��!�=��Ǭ�EVX�̼��ח-އ��G?u0�M�Bb�׎���� �����A�9JڿQ��,�����=�lk?зk�ǩ�eO�*�?^�����,��O�[��I�+,�O�X��T~��r�?�y��Xg:���b]	��Km�N#��:,��kkG�N˼~b�FisJdb+?��Ƴc���e��!��ؾu(��JVewT�y ����Dp�p��CP�W>���ق�@]�T�-����[.�<q�����󦁅ahlA9�[�}؂a��9s�}ckV8��~��DV�j��AY�D���O������p���W@�)�Co���]��A!��/��/�|7��)1�^B���A�~��0��	����*�Uk��:`�(���Ps�E֘̊�オC?Ѥ�:вߴfI�{K�����q��2����q�~"�dŔ�m���BnM!/����E���_���W�o��=�:����eep��* 	�����m�Pb�ڟu��A��e �� �	9O��+5kQ&�b�uG�C		�;q/@�ē,H�BKl�=ʄ,/2!{F�*�dPf�F�G�4*�T�2��P����-�v?�¸�	}��ګ�I�;Z��+/'(/fP������4M<����:��B�TMlߓ����iEک��p&j��밧7�N,�>�ZO�q��a�J���*A���;�b�iu� ��4`�g��Ò+���b��,,����T���i�3Vx���-%@� ���E�?yCR�y����-a�O�%�şS-Û�@Phs1���Wފ�	�+��T�a��bBQ,���Hٓ�^i6u>��������2���*��桏��nF`���$5���^(]���e���q����ڑK�fx�YU�s�����%�6�s��D�B(f�sb�R��~�Y������YQx�#ό���฾��y#EW�R�W���N�D� �`�.&�cOi'{�&��}P��;��k֏�f�-�IuϬqj��o�Mٗ�|7�����O�wȌ9Fe�	)~���\8XBI�{��+���V7��Cº����y�	�"p�U��������d�.�	�|B���F��wF�g��U��������-�r7Ru���� v�;΋6��#?;���U�mKXj`A��sk�q�$�i&�s����}p���;�>��-�m�z�R�X�[�~�����P�7�P�b��8�f�M��p:7�`6��� ��I�RA���kY#��{���c���7j_��X��tƗ����b�����64���i�Ʈ�;I�^Mw?���A	�Ak�e�/���Ҟ������mÂ�@q����9��d�_�U��@�\�4J��u��" �ߴ�B�/y�����W�0m������N�c@���̶l�  �I��Fw;L�hbff8v��O)ݕ��n�����u�i��~���U-�
i����M,:����tQ?4���v<S$�ϷO��W��Y��ּ(�Xj*������,�3�^���1�8�v�8�J�v��-�E^�I��u7�p�;�n,���[B˳������1-ͦ"T &H����ן��w��D
H.Ǯ��j��匴<�<)#�G��y������A��Tҁ!*��Zu�}_�2�";�o��)ίެ	�x�,�.h�C�&����KM-��	N�	fl�	��}k��=P���������I/�2_���D*������*nk�u���Ǣ� �jbUڊl�(5���t�]�!���.�lU���]1���شO��х��amU��rU�ģ��\�x��%���ն�uz�Z��)�����n:�AK�$҉S�{��T3����;��6�;>�����B���}�P_u�hJ5E� bJD�����^���+_�Ե�es�����v��7~X��F�L���H�8Ռ�O�Z/����DYD���I�c�ԉg
��!6��3ĲKiR�����+���K�iJ����D�*���!xQF2k��C�����~�="$���IQ:,[X{(|Ҏ7w��{yh�] u�5��	˔Ӛk�c�t,z�~kTվ�TkL�V�o)o��Fh�^ �*�S_�$!���_\e��y���UZIaqƈ&&d|/�$1{�i�yN�e�i��F�>���� ��]�;G�b�=��E�����aҽ�0��C8#�R������mRا$�MM�?��������^���Յ��W���t�y9��7y	������^E�
�f�x�TZ�t�P�����Fʘp��������Xhs�j�� �g5�y3�E��FFw�;���Y��y+���@����r<���u)�Wݸ[MM�jX,���x��JH�R�	�������x�S�n3ϕ�Ƶ�VgI�?Pk6���r�-b�h�C����|8�O�8�D"�����;�rX4	T������`��_�� =W��ã\
f�ʩ�WӠB�Y���jx�����<7.��c��E�|Q��]��h�e����ʃT�w����^�_�����fz6��-�êm<����OO ���<�x�����D@�Vq��k���v4��E1u�o��5D�����_P���܊{��l�4���T���'ֽ�ȅ!��y86�>ߩ"C�-�k�z�[[��Vy������,�xl�dQ!� ��7�s'��3\�|M���C+�{[I�H�P_�����#$�#0aT�%GN����=�$� {0�l�������:�AW'��{"ܢ��^kJ����Gj��E��|�a=����z�Q'���`�Jn1\oxي!��:U&R w�v-�g-˷�h�	B���8C�&�3�U�Z�#�v\��v?ځ����������`�����Z둇�J&���Zj����!����}�S�G.Y���aW�1�/*��X�V��Wͺ������o0�l�f�<M�G�
u���魜�dh��)ҏ�U�� 
EP���9B��p�n2i����h%�y��"=g+� ������[������R���8R��3��,�e(�2Ǡ��p�A�q�Xi�y����/�f���"��2�_&:$V���q�T��\�LH���k��v/�Nz�E槦�um���m������6��r��,����q���$d��-KHk�2kYs�m_5yI �nq�)w<��1F'^�	E%���7��r�
4���;�,l΃�!�q�3��N��-�$2�t�X����`���049߭��o+�%���s8&v�a��Ԉ�"�̡�nG
ON.]m�(�M"|� %<O`-�4n�P�����u���g�ZL���C��ڂ0��.3L_��`�u����B��I���&2��W���7��U�G���!b)SS*W]pn�����Ym7�$����By��<�%ʃ��ɋ-�'&�� >3�������ed�$<����.\1��ϒQ�����[ż������}ΐW�(�nPop����b�m~]#1�;�&nq��/3M-1���/�kc~��5{:;�s�F��	�9WVѫm\12���/�0���<`�B�Gjj�[3�3���>� �^p� @3���X~�q��8�;�1F�ͺn1��}��XS�\�'���,�F1G�����y�R�<yY�t�����(�ܧ"������D)�
�snaHjz]B'K�7�[���	Ԭ��SiBh�Bl�����?��ԛ�Y}ߨ�Ց�9�Cce��wʌU�.����o;���?H�y�-|�]��2�$.Bd�2��Y��)+���ó�j=��5<��$���]Ēvy�?m0fm`��4*�z�������}�s�^k��ݡ$�5w栗�+1�0��i>�:F4��_�\d����5�++������i-�����zw�o��bs.����4�<Ih�!���OlK�QU��O8��e9�z�� _ڀ.H��m�}=��Jo�L�wŝ���,��m�~Bb�F摋�lGE�������a
�e�R�4�4>d<�%3E̿@%̷`%�^�o�g�ʽ2B�Vc�
�<�D�e&�+�ώ�&�Q3T	˥�Ƀ�T�E����#g6}Έ8�2��O�=̾R��[?Ĳ��&������|Ql6����nu�Mr�83,xa��A�F�%|C�:&���h����	Aމ�+L��;H��T+�(%�z`q9�h��Ԯ�p[�-^�"�I�&o�A@͒^J�TP����^#짔�U��,ݢ!߫�������Ei��Nl���S����L9�(L��?Uu���v/j�w�_��[Z�v���)�@́�RK
�dn4t?F��EU@Y�8�|��T���$��d�=V؇J����h�X���{)x/��rw�����|7\]R�;xv����	s0��zLL���]���}h�ņmK�Gbz���Z�R��M��U7Ņ�C3���?"�G���VZD��aȮ���}�Y��	�w�B�EC�U������� ��wj��7�W��jk�	�t"��:��S��ʌ�Ә�%�D[0�FS�&���ѽ\���Γv��m���{\�j�8� �+2(}��t��!�X���a"�ۋVe����ɉ����� |��i'\���^�b������&rM���c�A�@�����:���C��Q6_�$���6��<e�ƙ1`2Dw*�������n�}�5�K@��@�8�Į���E�Ė��V���é�	���1���3e�x?���ʔ��D�u�*N��]B�{�̍Cz1�ţ����[qPz� cuo�	��w�K?���|�bײ�7�/I��|}� �k�xs�����}���/h��G�2��:�/Ǝ$膈���|���ɱ<���Ϝ���>'�b7K?�R�*3�{���!��6��V���,�u����Hd7��L���ڽ��9іx;I�a(yr��4��}2�o��'�����|�J؇�ё,��?5A�=)|N_�:�CCQQ��Hi�X��ݲ6n���g��%=T�)%�#o���T���>�fz�$_9w����G�;���`"�f\�k�4u� ��rC�_��k�V�e��}���v�
�
!![���A�頵C�h�'����=a��@c�����n���xEw����H����ڕAӒ
�}˄���{:�t5\�c��G�n>Z�`����n����.�[:r������m,�9m���U�Ǌ�X�5������Q�JG��1r^���z�g 	r��v#��is�������R�P?���~����9��� �:ڴ	��?���9�7B��#&�C�I�'m�U7��&�BV� ����AÔddv\-�.W�l�A�n�{#ۧj�?7_�%@S��U6�i�?F�����v!����Z��@ӌԪ�ݫ,:����@s����B|b�	���7�kxl�l"BD����䥂*4d(!�Ȟ�M:��.��fkt6f �0V�3������E~!ah G��BE���M?�$����|�b%
�٫�DU*���k:1��k0�r��^3�zY���ѱͻ���o�/JP�(�c�� �8�{ +�C�:�z���q�x����U]Z���W'#(z��;P/��A��0^`׬B�YQ���:r-(�O�����^�	ZL�AJQg��t.�	S��q�	�͐�)-��>��T�g��!
�@{a?*$	I����}�կ�`������,���A���0��%��>�(�P6�^��i,�*��[� ��I�N���	���@\�
ub���[wp~ں��|P��� 8w;,����cqH�������B�CmYAb�c��S+��1�]�^ͨY�2�$%� �C2�>`ڐ���JZ�m �u�{�y<�ia�⬞��<���h��t��>d������=����x�����6_o_��\�q��`�3ͧ+ak�$���H�CJ��'�Dq[(��r"qB�T|�`xbR���#�b+h�6�A
k�Bf�Ai����Mj[8s�'� c;?c�R�a Jմ��j����0�-��^v��m���G�[�	n6],^5�w4���R�=�(Uu�=�����ۮ˕�?0�M @w��k�bc�D�F�-�{;{�]a\�`x�~��J�4	b�#~j׸,� n�k�5�aRR�/�\��`/Zϟ�wdݠ'���L]Bn!j���Rot���KS�B�o4��J����Nh�a�vw�D�����)π�V˽9܄���7`E�i��c/�T�����<d0�,?!j���������I��	�UMm���=���`��)�гZl��z55��6��Ύ�')���g-\�پ�]�h3�L��������!x8�6�D���V�8G:�e���s���`��%փ�3�"�a��s+�,��;�tԔb	'��\9|�n�����)>�}��C���_���{��-�z*xS�g~���6M�|�Ly4r{_Cުɫ]�-���'i�'��kɓ��&�X��_BRr]L��*x�am�.
|�%��,O'�c%��lv�+�� ��%f�� J �XY6\�tV>��3����&3!�;�r�qj��^�`�k��O(/w])Z'~nKy@��m��Ej�d����%�npy���tk�1ߠFfL�����hd9���n��k|���N?K����)x��:�E%ج|5�z��c ֜����@���q�jT�j���C���oݞlUo���kq/�wۿF�&QV���r3��k
M=�WՌ��V�YӒ?o�B8ת�*��,�Ns(�Hn0,�P^�`_r��s����&,z����nu�n���� ����"�rw]��5��q�;i�i�!�^ji!Q&'��*M�_I���4I�-�[�Vb+
�g����k�W�I�]n��In#/��Q�d<�;�ַ�rȤ\0#�ċ*�uc��@U}غ�	GP������A�Q��|��q�����z���a�7 ��"%�`���K��Ͼ 7D邜!����A��sAh�޴Y���'y���.݉ŝV�װ��٥�Pv�jl���>n�+A�H����]P���lX����%�嫀��%��7m�R���-�]��%f�j�f:V
!dLl��	5����w�{�	��l��8���?��2'�����͠8��7�rJG�= �o��ꨔkL�3fo�葹�Ȑx���2��Z�:3�w�&���\*7�B̱��U������9����|2�{i����V,���Zu�Wy=�޵0� �������	_Ji$Fe�m2oǤ�$`���d3`	�e���?@�<�T�K��=�����=�(�p5)j�������]����n��|�H��w���C��|VT��.w
��Xbu
�I`����/�/��ݷ~0�Qk$��Gǧg�ȱ�����Y���iIy��Jcb}A6���1H�w][aK�1����*z�XSF�����
ӯZ�%W���U���\��`�飯������eٶ���l)t}.��z�ǚ�vV����M}UL�j !+[0���U�4�D��,��K>wtf5@`��J�o���i?/��3n�����fIA�U*ǅx��dE�^�[�~e�o@��R�Q��N�Pw0�鬌�~�b�ۂ�v�YB��S��M���Iњl�0i���=
6�w~_f�X@p����N7�����y�,^��d��z�n��1�h�f���{,Dfe��j<�#��V蘿/�W�#���#��J�/J���2����RMxRk+#h��k/��U@O�!Tĝ��*;���Ph%n&X����;@0�p? ���y��tz�	S�?v� vr��`�<�'�ּɂ����=�բL������U�϶.	��Ηߋ������h�r��3��+�(�bz��C�"�\�/�qM�$����S���4���0`S�,�Hߵ�Z7��u��T�ރ�p��_����f��
�fC���+t���������A��k�3��LR��L����fI	*��d���uK�4熣/�>~��p�2��kԐ|��=���`n3!#pk\��R�	�:�9g��6NȄKC<Ą�ZJy�!�pol���P��ZY�H(U�,���;E��/s΍o��K���+k�bRxJ_.k��D9�W��1���Ց� ���Z�D7����W����u��R0��6-6�9B�z�o��%��CE����z�\Ya��O���T�@����yV��hR;�"vΨ
хr�B�	���;�����*	��b�FE�0��o=I��5h��2�䅇����Z،f��;%��ZM��/&:���˧���6K>�J�YD�,�����=���S��p(P���9� �rb���T�V�0�Sm�Hu��I���A�t>�=lN����e����K�Q�٘ؿy�2��,⿨x HQ�a!�>1%?�m��Z�F�Zͺ�����;!Pۨ��慜���묚`��Tꈯ�ޞ����`��s�?G��ɾ�Co����~���E����f�
/J�yB��b��a�N�w~�w��|c�c��{�#g9�@�!�=Q��b.���^�^���)����R��)sR�:�yKh�T���O^�"T��6��w��p2�tB���ls/;D��Ĳ���~e|��ʧ�~���8�C���$3��P�g:��9��J��r�s���=b�N�m��b�0r*f_�,�2�'�~`ty��������,oJ:�kγ�k2m0�\H�7Hr���z¾���P�6��9��σ2��;�8R�o�+�y����F:#��l�����r��~��&"C�۟(O.~!��6��ԧ�l�h|u�l)-�ڐ���Z
�h	]�G��(�)5l��3�m�%����0��ؐ���2�Nl�R�͵#[��y0�x��4`�e������jVЉ��%��ܯ����P&m�90�Ý'uL���o�����]��9=WO禩{���#vX�:��s[�1���[Sf! ���q��D��ty���¸��
-$a�P�-�ߴ}�͌�0oxΥS�l��5���G��Nާ�xA�qYvsN�;+J�\f>l�!i�bd�@��a��L�>'���焒)��O[�Z#'k�����Y��{ �Ô�5�����[�&�����*�������"�#��b�ֶ}� �n^��2i�d,(aP��9󼑸�Z��wTW#gk[����#~�q�q4cJ|0�h�7����R�ݽ�G>�8�m�K��ݚ��E6pF�&ߎ�N��ΥD���9�=R�b'�s�&6=
�H�|�%P�'77��Hs:��?>�^~{(s����G�Fg-M��'�����a������'{B��$�gJ�N���G?g�^  �i<��[���Š�*��>e� �!���/�R���Ri��󛎦g�֫}d9ZbC�
1�b{dt>ž�y�_�u�W�m�EE��]���ݓ���i�L�w���#�Dt�J�[*�>������"���/��1Y�4-[eqB��*j����X�O$Y���9y�~��Sr�H���������%J�����*��09v�RَW���S�ffO��ah^i���^�h�4P'���\x½���=Us���Vtݬ�d�t�<��
���89�����츫�q@e�A�^s���O�c�J���� �k�?��uWxg��
\�Բ�'ws�{�����GH�0�#��_S����g�l�Ȩ�"��T�H����,cp�!�d+��mTF���&�:��ߎݨ��^q�yf�A�*�n����/�(:�ı��� $�LefG��ɍGf"pI_#���\>�FF����\��z�BɃc�	t�A&b{��c]��Y�,��)����(L���e=m���[��*�,-`3a��%ޣx���6����A��Bk��*G����I���q}�5�C�c�����
9�v���Z7�Ot�N�!;���)�,�Q��y��PgJP9b������,��>����@���BF�h��~��QN{�O��*��*t��M'Ϋ-�ܿ	�f.�w����ڝC"�s���~���ω� �^�����8@K�)'w@�"�+|:ع28�F��h�������O-��."���q���MP��i�S!������yp5�*����c�ޓ
����z�L,	��(EH�#눬E�n��I�#cQ���s�4FTP�w��׷G%�p^�7_�k��Z�~��ܛ���o��&��s�ۼ�4	1�|��h\��%�z׭�X[���Ӕͼ, �ƙ��Ļ��xF�P4�b��� M�Y���S<��~,/  �fkZ�*f \U��˩�) F���Z�|\q%�F7;
߸a���<Qϑvd�#O/�|�2�5��C��Y �XN�`L;#w��W�[ֵ�' m�y/��$�GW��s�0�	0��FN'��8��T 叩�C�����B@����j��|۽�-�n���s�����0[�gj(Z���
��Drz	�%��*n��i����&�|8ucP��JV�o4?�A��^Fܟ5�]�Ԟ��D�_v�yx���2��Co%b�탑D��Zr�����Cn-2R]¼^��vxz��B.��1'�7�k0Y�S>����N�M��en��������wPP���܏_�ټ��"7�|)xN;=g�IAO�vuI/�%��~�Z���=�B\5�*�����㹬�C�fj��>���@OП>� ��BA�s}�R�,�y0��G��hNiF�[!���%qN(��V������]���(����7^�o{͘a�kt�� �F4v 9u.66��rS<jy������*[��S�D�!��C4�z� ������-)���g�v��U�
�u5A��������$��;uh�Sİc�D*�UW�����x�T�1q*+��1����,�"�m��3�U��B�{�:Tӳ��JҒzvĪ�&�X$���g���T����YZ�z$24v�.R�G����B�(����⼘#$�[]t��/L��נ葘�Kө����`V��QgsQ����dU�x�+�A$#��S\Y��D�J��Z@z\n�F�S���nF3.4R��ۍ"�R�]t�23�J���i��^>�Z��A����2�6e6��$�9J��g�'��=c�����X��Ga5�Ń���G�A)�Qp�s�A�y[W���1����|5$l1^�aR[����Z!@<4����-�_Y�����A�G�9��E��yN�8Xo'�H�b���L�h!ݭ����>c��z÷�)�]뒌��{u>�Ʃ���*Y��ɂ]�����`,�ϒ�-6�j@8g� >��
;F��Dm���v���aKP��/R|��)��l��t��T�ڬ�B��]�n���a�_0u�a'�[{�#��'�7q��Y*�����Qa��c
�>����!Mȩ%�,��!/0��t�w,\(yU���9%"\��߷��i��s}���?�]��O"����z�pE72)6S���\�)/Fk͎�xJTk� k�`�O�ǐPY{̞*|���D�,��Mf�j>�#Z̯�܊ꀊ��P؆�~�dL ㈢������P�u��sS����VZ�S=���3���\nV�{�Y3[H)25ߥ��F����e�=6�b�~a��lO��y�Cx�g���d[$�w�����C�]�` 4�E1�5,���g��`��X�:`�-ٱ��E�� ���`� ��.-v����Kd�����in�ǰ 4؛���|m�c��g�v�.�a%�_��|�Nl2��$��*~7���?��
�X9&��F�����#c3𾤞^x���%f��'5�@�ִ�AZ����)�����]#��`V�@�): EW�8����z��?�[?����:���x���xŝA���-仇੫靠��]y�z�b�r#��y��E����#�鿷�mՌ�59��%6��4#T��y��ݟYb?�}�B{uL�{�
8��j�b�;�z1 S$#יR��XXXzY����֩�n�<
B�M�[��h?��-?�<s��	�8mce��퐃	��Se�^C��h0oRqï�;�cg�N��'GF�J��s�4:�9�'s5�ֵ���H\�V'��_�A�A~׏+��3��R���J�b���m�ԡ��	E��1S
)-�ZLeN��4��<�j�5�
�V}��3��x���Y&��S�qL����kz���zZB�ho��ln˥<��zM�`�B��Xԃ������;�:P��̛-ң�s�&<&:x�{2��غʶj���S+[�ݿd���\�� �0�`���l+0��!^Id�6`��n�j٥�Q@7\}>Δ�"%z�KI�Ӂ> ���!�񸸯����ģ��Nuf�ꤛ�D>,��6R�K���J��Ԯ&q��ypx�ᯟ���HJ�����GN�`��jt��Kaig^�6�> �"�{M�+P>�M����y�W�-uL[Q���Ŋf-$�^��0>�H���"<�����IԕQ3t�����Jߐ���J���`pc*n� �Q8zҜ���|�ҫ(��*�^�@	atn�<�K�����1�/һ �]��hݭ���MW�;����;3�,P}=:#��Q�IT��mk����	�`u��F�P%r���5��4�V;R����C�9ʿH?��,�5[f_��iX�q�MW��=��'ev��E�5x�w�]���(�P|�z�:��CP��2�S9\��/���/eN�!/w�AQ\��e�wE.�C�Tw�5��D�K�-)��p�}j�Zen����'ò�%�f��[T�s�� `B� ׷��ȹ����(��{�R��m��P���#e�3�p,�;���Dî*by�0A�7%�.�'���\OB����Q�-)���!�$Ĺ�I!Kt���J���++(�������kƴ8��tH�n`�=J�X��7���7Ǟ,�#��⹐�0	&�VnJ�����$ݵl,��t8�����"��ζ�;�
3�<�n/qxG%
�|yk�_��}ړ��_�5zz�5��qTK�	�w����� �<g79븁��ٸ��˙ Yc��o�����w��Y)�[_m"`�B���C�j�����.������MRt�����ٖ�yGka��)B4�^M}�E����Y��K�9�/����!E���-,"Y�!�S�����E�@]I?��~�9v���M���'��?T�+F���쉙т��X��@Q�[�V�x��4)!�b?��"Ȉ��<�5�w���݋�%E)��$����$V�����7�L��r+Hc$(�Cⴻ��n���hس��6fy��7�W��4jb�2"�l$䀥�:īl�����Y��HuHȚ�^Y�?7�^�B�xJ��4��q�	܉AR�]}��J��ƣ\�j�A	�s�-�s2AMB�v�x��'}�ɩ`*�vT����
P��Vk�>D�2�gBa�>L��2��o��Ը����H����:�ϡ�U%BKi����KT�J��EN:s��}�B����=����b�� ���nc�B;7vQ�V�<��}I&���d0b��F�L V����Լ��f��g��d���6���C�C�IX1�ۧ��s!�]0������_S6�&-�H�$�3�Ͳ�y�(b�P���H2�v��>��St=�H�����R����t�*�>C���T7;?z�lKJk���@\�qp�P"e�$Y���v_�{7�>�fʱ�wu�J~��0���>Э/�5ыh{<=oi�&J9���]IG�����e� #V�
�*_o�����3E����C ��M�E%'J5�lI���C�����爓�>_u�֌��Д'�n�J>�>�/�}��!x3k��w��P�����za��Zn5;
�A���j.9�����_V�tN�(:��b".h��q>�ĔEZN4q���kR�6X�o��\����|>�!�H����Əb)�U�SQ��R�hN�e��ozFg�X����!���(���U�Y�Cu1[�������Jj/=/«��cpL�*����7���EWh��:����+��ܐ�j��������]Q~��l�*��2~��^� Q���q�Re]ݫ������+ح���a=�=b^�p������Y"�aq��X�.�\��r�J�����nп������8�/OQ%�w�;������@[g��jSz�@��K/%��W���@�#y�*�o_��g��������7Wթ�kD���N^l������H�ot$J���K�j�R��qîU80B�?��ٲ��2�; ������h�����;�:ݍ/`ϿL�`���b�����6����+'��~�-d�.���S�{52�붌W�öj��D�%0�v[�R��S�̀��L�.�Ӊj���?��s.�>��5;A����N��`�����>�+�A���:���Otw����
KH1��?����@܈����
t�����d�R4�L�to����+so������[[l��̏�6J8�p1�w��#ޥ�#�g��6Q4<�%{4���U+A\iHy���jD���n:�.X՚����DT�S9��`V(w%�-���JO{��>��@��.5ǯSLa�
�&��|L�o&I�'�4���MO�ꗅ�;?O�1B7�>F
w�΂�7
��۵�Ľ=ӗUi�j��T%��+��t���4��?�E:��萌r	`���ǫ~XEns����#��_�{Z ���A�1����Ix�*��@��VvM�^@�|���9L<^Yw \ e150�o�el��S8z[U�1��.V���)"��+��"����{.�Ǹ3R�bQx�hcZ5`\irV>�;X�#�/T�G��hte]�MA�2�]��׉v�۫8�^F�Y���ݪ�޴�I/ScYG�]hm��
3���r�%͗Y�m�I�0��ak%'���ۙk}�t�Zzp���R�	N�\ǒ&O(�IS$�׺U@���M��ܳn��P�r�cP��0"9��aԾ`)5�-h.�Q]��μU���$Y�)v٨|x�+�/��j��B�è�t�Bis� ��
���*� m8�Y���؄�(��������󽺏F)M�)����Oºr�r�9�Udc�`�6�o��7cL���P�n�.fO2t��+�~q̹��؇���Ճ+/n|���tz��1\2>Qz3g;<�A�w� ��{��"��C���a��u����P���^ �dbY3�>��O�y�͖�7�N������!7N��hA�ɡ$R5���J�L�]�kxuC�lU~`p��O�DM�F%�>7��7�M!Z|l4Z	`!h�G�� �-͆Zȵ�q0(�d�D�j�3p�e窡��p��}1�C&���
s4��������SQ"��H��h�?[����(#��j�0��Ø3%�=���W}��~����Rk��1w=��t�b�Bx��"�n8�#_i�r���159�i��!��)3��]�6Ḿ'����	���$�T�u�����N�tz�M��@;��S� Ԉ<���X�L_1I���	/7�2wIl�;O��sdL���⮹��*=�U�DB������48P�KyT1"��`l`F����]���V���6K����˩q��U"�3��f��-.N�l�ُ
���2��w�$�ج����B��Lf5�>�V�h&��� ϧ=3h��'��O`�􌥠&���� }*��5�e� ��)�jhGw-��dvlfs4��N[���(W��\�����B-G�n����$6�A=��w�~����2P��0R�b���jg�5���n�T���򺜲̷����yT��lɉ�x�nR���C4���ȅ8���Im~�aW�
�z���n�����3њ`��?�F��|aW��m:���u���Y�G-�"0��X����	~WJ�Q��<J�	�(�'A �"�k�)�6�9w�Ѐ�DK[[�Sm��9��%ct�Y��@�\���:迯��=��QGsG��g�5w�zY>q�Q=��K�^��0+��U9����zh��z_�:�:�F�����;wRG�"9�.���ݯ�����s����d�]��=˘��VJ��f0Uv*������ms����Řj�n|�� r�v�����/�	��MA�Aq����hhGN��(��;?�d>�R��iZ>�i�����/n�k`z��l|�����S7ok��.26k-r��ׁ�}a[7�7dW�*	�Zl�Ʈ���^dvCL�:e��}�u z*�q�-����ǡI����sV���
�Ķ$1������"{���b��Qj��3��č��%y��Wk�.BsC��G����]��(�ʸA�5\\<�gЗ�)���9"��x�h2
'�[!��X߽p���J��w?�A�kv��K`�۞'�i�ǥǭ��]5k��x��A���x��M�e5�+�qp���#��p��v��/�,S+?�V�+Y�@���a6p�sQ� �:a�g�{�[��vy��1Z��(���-�ӌ�X�)l3��Sy z�A0ȋ�e���~�C���B]�j��j"aجB�w:����Nx����,H���$��]�F}���|A��>�Ϭ(��kp�W��ѹ�����i6H`�����ɑ�挥�[»wMf������>0v� ��\	�{@a� ��@����%P�VLG�h�d�'sɰ_�u�`��X�=�f�;�݀ۆ �/t�Eut^D����6�Ee�T��nF�\���Q�+�/�b	�T��9�=�	26�@L�����
nAfz5
��qaB^;��e�<�i7�Yh������PJ��V#=g�G��Ħ�����������ɨ���H��5�X6?c�	+h�fRb�u@β�C��@H��f):���/�6�i+QZ��t��w:ϯ2d�K�\S3�Afw��B�R�m�%�"8�Р�I�B�}4˲+d�:n���Չ�c�2L���j��|��vq�p\�<2>��W,�)��ClNļP��"N�����{u�R��%v�=�[�!P�O��l�K��A�$c������r�,-�H-B���I��>v~K�5̺�= ц�)�9n8Gse�?S�I��vxȜBv��4���V�D`��AsqG��m�KV)�?��";آc�c�T��z끻Fot��S��͂�&�p�W;����/$��@֛8���'�X��R�%�P��a��K�	l7א��<�����g:)�����u��`����[KԤ7~�`���*���r���6���&�|�긽Gc�tJ�%�-�vf���j��n(��Q?�s[��C2g3�m�3����}�Ҩ�H��E�؊��n�I'�M�cQ1��i<�zܘ�!c:(E�]���ć *�Z>|����U�����7C��O��f����!� E�Vmf�9t>2R����~r��E��U�K�]�2���<���������#�o���l��zR�e�˭p���́%H?���M�� �=����b�e0�ʃ��qz&Dm_�ʖ��I�ӰAf>�����Փ4|�]�4U����������vH��?�����˗R�J�
�,�����4=0y7�sqo�2,I
"%bF���R�T9����>�Ϻe��#P��#^f3�&c���_���NEˣ/�$}b!�ŖDD9d(�A�����q�3��Ο9�bC��̬v)j*ј���r-�X������X����Չ����ZV�R>��� �K�S��ü%7��Q�-�ȧ}��+�=*(V!�R=*��a�z����
�M �� p��IpK�d i����o�;r�x~н����Y��s`�=�$B��Y��,Z{��~���'˨
�y����3u�p�1�_��)Fy� �њ:���fC�"�R��Ǽ�!�C�n7�j�g/���\�!UN6�9���d65��5�8e��6�i���6�+:��2�٩_��T!~��xI�8��؋akUjj���4J��o��¤����3?���H���ɫA�1�4��w��!~R��MT��������(�Q��.9�R2U�e9F_D\�FQH(#�[���x+�-S}�V���%3��K�,XګK�N[�L@^)&o2�f��
C��MAD����	6jA�	�`��;=�*����lCFo��B�OG³c㨖h
S�Hx�����o���~ruxwxɲ�I�EeG���!x*�v��&�B���>! ��'�1b��3�����?�Ք�*)ͦ�1O{Jr��u�`�S��s*>铱��)!�)&�0�u�.��g��]^�c�Z��H�y����LF�jȞc-r���R�Z�C>�{T���4^���{A��3L��>�,MJ%,̍~��B9��H�]��G�R�%ȿ��3�,|o�ZH����~�¼����M�U��۲o��>�F˦��1�n���Q����8a�-��`fS�p۫F�|��� Ö��ҋSڬ��o�EJ��~��xu�}��ѽ�����;��������0��J��o �W�SbU��H�=!����	���ꌚi�̎��O� �狢*6�qQ[H���'�O�Ng�?�D��k��kL�;�^ػ#H�#y���&�	�?��&�:�;!�L
�'p�#�.��A�ݸOi�M� X�vˠx9wQW�o�K�
�� �,C)�6w?`�R|tiԦT_y���aƎRE2���/��?���n�:\��|��I�X�--e(�ԍb��F;&p.)���=���^���{F�؉R�GI�0����R�85S����,0B��ͥ�Z0�XT�TM�J^*���F5�+w�J�r���z,�u.q!�|�����Ȭ�F9�b?��hw��Yp��;88dj�P�`�Ji��AFp�Y�;�8S����,ז�( {���[�qj>�Cu?u۬�R��;���w8�S ��g����֭�W����,�s�0!BS��w�m��Z�Ȥ�ͨ�� TH6��`�A��jJ�o&���_8м1�7�9�e�P�>�h�w�F ���!3��r9����$�ų��;�����Q�j�&�\�4�+ED��1j�
s�V-����eUh�*��!�t4��i�W���dGI�d�rf�"ڿ�X�R��e�fm�CCXG��x�=�1��>��oEu�\B=������Ca��	ؑ����|��o���G�d�v�[��p�W�xD�.��z�;�z�O/
�Q8|o�3���t�>HH� ���0�v�cp� ���L5�ʳ��g��@ O�M�f�nM+7�N��ˑ��UU��jB���?-�s1���=w���	��3��/~��rk�-�|�9Tק���6Q��l�}�V�u�~A
퉵����o;ͷ�F��-�-�+�8�YR�9%������Ms˳e�@�T�gΏIq;����vFڦ������ ��2jmOK�$��	��|\����0���]�o�pŹ���ۍ!6>LE�'��,����cƙ����jK�C�r�F��o�'��)����Ø�iFrPӈ')B�o(
�l��B�,�q���/�bF�|�xL@	<+d>�ޤP����@i�����+�+��#�2�#��Ǘ)$����38Қi���.���P,A���k�p�Ws��n�6��g�3c�\s�~�
>���bm�mF$���`
�=������@������ʱdz�7xV�W�v����Vبd�U΁��
�V�Ξ�m��Q�$�x#���V/Fo,Z�~W(����>K�N�Z35�k�;�^����렏����t���d��͍1k���2؇�����*Fď���|v�M��/So��������4��[���-��)#���(%�7�6S0������
Di�D#X1��Ŏ��{U`���<Z��?����4�P���FKytc|
Sv��dhɇ�?�;v��RV�J=��)�Dm<g6�4KOΙ��<Kq�	S߭�4���us?=<�@�{��`R{��B!�����GER,[B�O-5���82&.����ʨ���A�pS4÷4�dL����9���5���NU�4j��ȋ��cB2�������(L����v�@�Z� ]����{���e�{��7�X�\W1����� �����i�/��a��J�󋆫_���;�n�݊P���
���b��U�\�N���H���-��Й�l��좧!���b��N̛�ʠu���w��9d�Zr��ky�~������g���P�Z��7	���,��;j�tp�N&�cC��\�!���w]{��8�n���6���/��a��yI�䶡�_����*lћN���c��w�?��C��s%������*2-KWAA�n?�c�\��M�ps�_��!��P��0՘��w).�t�*����r��S�f��{�h+��dn#�/�}5����rk��<��{����JDm�K��_�@�t���?Ea|M4���Y6�W	�D�>�th̲]�Ҋ3$:�6;8��u}"��wi7��!?��o@��D��KG���/um��UZ(�J�z!��z3K	u?�?	b�P6BV�B��3���źB���:��`~+$��b����e���x��+��Qk�!/�X(㶧���/�t3���|p�`.�a<҂�?��QQQ�*)�aM����=u��"�&,L������C��%��-Zs_P��"�&\HAD�aA�
`A�\S1I㷃N�s -�?I�
�y\�e��i��	��n���k��PB��6#�K޼lQ	c&W+3Ԋlr\��Y:'���!q�����E1F)��6��t�O>�ԇ��3�p���a$N��\������@ǒ\3ϧ�W��@6��w7�1,�D�3'߸�V������bS�tO�d�Q^���&���	W���1��u�Wm��A�n������[��D���[2�yE��%{57H^�:��L�Q -p`bTR��镗�Ǝ�~w��t���D^b�M��?{]�3݃�(N{��ԇ ;�®�B�fp!+ƿ�EY�qR�������$�D&�P��"�ʙw4TI��z�A	�9�ɘ��0�H�-z�!�CٔM�����K��CѰ�5�E�K��	�z��*���T��ISp0�K�5E�/>1�)�������ftfK��`O�&¶���]gT��f~�s a�X �Od��b�APi*>�KQ�:/U�~?������8*����DH�z�9!�T�R��@�G���x��Z�8�[�ʺќƆ�c��f�T::��|H��K7^�s����?��%�𷁌%=kS��!�yS����M�WͰ�Y�M�pS�(�a��ڨ�̲�_U>2@�,�P�^d`p�NK-o�[(�s��BF*���3mg�ڙ́����h+^v� �,�X2�>Z��0�=-�0�W���� �F�Q7� 7��QT�D�����t���IWv�%ÉFa>(wܘ���1SO���"�i�{��/2p|�7|��w��G=+�eB��PB��xa�A�D�wn��w�Q�3�Ō�u4�硔	�s7v�'F=�]���y�]E��wb�` �է�#u�E��^{�0孍����l�;!W#����nD���Ix�r9�W�35_��z��,s:���YIz��&�X�������cG�.
��F��� �r�Y�qɔ��"�A�z�HU��_Z��~3�	!��8P�d��M��P�����^�4��'D�~�}������K"����/��O�1�'L�{���3��/�)�x�;�����)*�P!��u:|D~�529�1~��")�b<�6�����=b�|���ͳ�L
/��e6g�2�n��;B�[�0i�ۚ�m��xA���7]eώ�`n��+�@��C�&L@�.R��H�!�h��P_�ٝJ�@��@���p:D�Qx�^��]���s�#ySOX��J�5*LK���(��s?�6�A �ȭt �<��$�O�%Oy�%>vߍv�)��HF�VO�\zh9!ҳ�,$�h�"Tg���򍾰��ׄqq�Y~�(Yh*WK�ghCQ	F�vӓ;��./��F�W;����"�a�;�`wZ�q.�2sI|��8�b�;�oN�9��x�Lb ��[�;#X>�r���@����.�R���h�w�r^��x�Q��N��6�I�r��׋�wk��Y�)?�I*t�NNM�4����	]��:�&vf�Z�-ug��@\#D�0����h��
e�"y�o���*��к*�6��@��P>�E+�[�cԧT�����?��b�����L1��2Y��!1n�fX�_�_z{��G5Zd|��5iO��9��8O�T���<���w+�/eT�t�>��7&0��k�L,/'.��}�S��/1��j���[�6�*�V'w}��tT]�Z�ѫ�#h^;�J莲f�*6�� C:.��n�#�����;[̦�/��HK�e �&s���~��A�-qava�:N}�	Y$�������r-���X`����9)pn�O�+|6��A
7�H�ڙ]�����/�2�乏|[˝�hO��"�K T����^�U��J������^	Xu�i�y�h��[*W��92�uy6�m6�N��R�[���������(w%��2Ś��9�%��J�.��<F�^$H���e��o���}:��÷���_�����O�܇I��gi��Ԣ�twiu����T����u;V�����0���k�EgE�A��K�z�W�@�b�u�4~d�IP��$�|�7�E,̞-��(�PĂ�F�:��c�Ɂ��Њ�g�����|�F��~�����e}�;ZH�&�99��U6�+I��c�^��װ(���j�be�}U���n�\�Y]C�;�F�2v�I�'� DOT�L�T�����cי{x��p�^e�FŇ�?q�𧂞n��h�/.6��!�	ވ]��B�^3����I�W��+�r
�K�=�|��O�k���#~�.l7�PL��@�z}V�o_�E�x��ȭ�=�5$�![�� z��Tg'mi��N�u���A7��`��6Փ�Ƌk��F����({�n��{��,��Oaym�Mn��lK@h�e��t���>	'�����}{�qLNA��6���^�������^�R�V��ei��:~�Bk�!�-�������_?�N�q>����.Bt6��c�5�O=8y�N�t,�V����
�!�]㟂�	)��������d���a�4p��ื��(�7@+�^үvr{WC�Os�1��ri� �(�e��U���s�
xSZl�v>ہ�Ɠ��Q�'�]I���;`:�%���~h��ؕ��0�Y�o��������h"���^v��)����8\,]0�W$i��ԳN�������$��q�0��εBV;���seֲ�FtV-O0;a-����@ڑ�R�����R�8�s5>���4m��a��tNR�Y	u4zJ�v�����O�l�,����Y�]��jsUD��C(H��MSO�틺�Dֵd;�ƍ���r��N���;��5��E�K��wq�������l��pޑM�*�!K�C�1W}����SI3�k���=�g�z�\lC���m����r5p��I;��-��T�8�=W����g�*�>���[�@J�����.�*UF��>z�`D��	�8�~�����?����@-�,�ց�~��r�����N���$�ڑ��೗A�����Z6~5�`~�L}�Y[������I���ˏKԼ���|�;�rJI;�uL�,���զaB��dE�ϸ|þI�U����2}��U"F�TK�ќ�	Z5iVw^�V�m�4� pz9�9��9�ؕ�e�H�k�) ��bZL�$K�p��\?���,�t��ǩ7b� �ͦ66�gjm����KxW��Wh��V�u�� �������ցR[g���q�����O��V��u6�x�3/{#�Nk�p�?��2��(C�?�����P+dCh�O*xt*�-޽	_�yB�ڌ;�5��a6�_j�^�p��Z��FbP�!*���ٽTT�w��"�b�Y�*=ڈ��Sd�Ҍ2�^B�V$?,�k��`Z�&�5�pP��蒵+���|va3=ٞU�����s��@Ax{�2��/�əR���6ӌgDB���6^PEv�W����a~����@�~�k���g!nA+ԨpK��n��c�w�*��үi��p�^~g6�����g?s��;.>�r�>��Y4�`���O��t���	���g����ROѤo]y���#�'B��OI ���$����6/���f�	z�?��a����B,�lWC�"��+x�����"`&5���mi����ĕ ���	h�%�Ⳳt)�h�LC� w��he�l�l�\k��m'̛Fk�Y �\K߂��N�̘ʬ��Χ2};R�WOyB�+W����]�bＢ��YMlqa_m�7ԑh0����e�5ԢE�=���o60x���#�=�p ��/T3J0��>@�+�͂��&N���I�Z'>�W���_Bf��p���z*F�x�~ƻZ�׻3�UJr�;�.7������r[S�#�+Dx�D�=��t�c�nN*�֔�%R\��G7[��8��Nqs�h}�r��S����	��0w�Q`��#J�D�{�5&9p��=#��oȕ���>�E���i�}x)/0b8�<b^���5F�c�T=!�&��"������:��WYY��Ɲ�G�c�}�w(Y`8��(6.#7�d�5�ӪՎ)S�@ٷ�[�]���HMXv�fP�?pᤲ��E6 ���g�H��w��G�V@mx\"�b�F}�:6����~ҙ��u~\r���ن����e�[[6:H:c�� ��|4"��6���ɰ��������xxIu ���162�����X��0"�?!Z(M����qm֓w'=�"#�fh0��i�9���`�Opt�㻖�ڪA���zκ�f��������ǎ��i,<*��,v}q��ŊX�^��n��Lg�3;���� ��N��/%�/����6�jl�ف
���ۦ�+23+�g�*�օa�R
2a'��j��kr�nYݥGo��eU�$�����V�"t<�٣��z�r�ݿ�ꍙ�p
#?z�M��o�6c6(��X�"'6�$b[$�v�*��fP���Q�|l3n�7" �俠`z-�ZF�8:#��t���>��@���i���'c������ѥ���!ƒ-hv���p 	왅JmjaY3��Xc:rƋ��/���ω�ڧ�;8@�T��HT�S�<@�=U���J�%V�~�i�������B���ذ�i��l
YG��d����W"#*��6!
��y�=423J{|Z9����mqp�@��-ڭz}& �l�/rB�e-�2QE��RM�F}����D�ݢ�w�h��H����]�w>
�?|E}φ�`�%a7b~��z�6R�B�x�����AQK��������S\�DE4�4*2���}�7u���ͮ�MQ�XҦ���w�x�{*�CP�Pet�]�ll�t�`J�a�,�f�}�.2̽��ޏ:1�VJ�!K*y��F�D�+�`�L��R���s�\ �N��2����FQҒId���_���Z���#��i�jH��2�M�br�J�q�{F���N����XMK�%)A�L@y��V֐�D�c�i��Z�<� �g���oK��U:#��؛n$�O�����n9�B�pI�e	.�a�t��t�عf��J����d H�Z�'���g'��%�6ʟ�0�؅��>���jJ� �8�MI@S�/�cצ�	�����Nn@p:�&�rwp���/�E���qм+���J����9��S�^x-t�o��j�!Y�,yK����yK/N��sԖ	���::�b"	�}$`�"�]���j1�E�6N,�םS4 \�9�HV�|�~��y�׷/��t����W%��;E6Lh`@)N%\7�p5�"Qb�솅��Ε�����Sh�!�a��p"Rt������B�w�zն|2���C�V4�$z���t�Ж��G�U�p>�3B9W�t�'������h���B�ϣE��X�72��P����R������q0W�@�ܷ~�Wi"��np�r���S5qJ�1�T�Y�_���X3�Z�U1�k?2��L�K�NI�����R�Hx�e)ӕ��ϛ<ޜ��5e!��f,ɱ�$:q�3��8����>��t�!ϊ+�(MG"!�R�S��k0���W�-̶c�?#��?5"Ά��9K�q�_�w���^�̊�a��v�rO�5"o��Q��$I�ӭ�V�:Eg�j\F`�I�e���ƍ��|O�"yH�m~֪�%a�Q���J�a%�䝹��F����{��,�vԏh��A�ګq!&2b��F���XU��N���>Y��s���~M�oO��@��o	�����k|�Y���-rt�*n4>ݞ�.�����9��+}J�s$���=r��:�ۡ�*h��
L���8���<$����b��L,5�aP��*�P��������)c��	�}�CⵈSڴd�y�"�O��4pOpL{��Cb>���S�S��z(�p��.��u���U�H�'�����1>v�
�.��6����2B+�������i���:N���9OYL���C-��Go/"��czw�X��92�g�D���͐��d��ړ�%�:+����6p��H�?A�ó���sR�4Gh�Ŵ|pMO�^�re��QW��R\�A^�rWM���a�}�W��OC��!�Q��k>�K0��&���.�4���'2�C�r�ݏ�"&�jO]=(pr��~���q�#��ě�5��ٓ�Tcc�.�kw��N��3_�z�hA�
n�g;��TY$̭7>����T1o#AxJ�7"�����D�8��v,ai�Z��屶W�����lʎ��I�SQ�21�_!;'���~|T�X��2r�y�����y��g،n�[�Q��@��$\��$��.`_�F�~l��cm�bpc
O9Qy�"�zYj�o����Z�B-K� ���$���A�o���A�x}��%�9�IJg�&�`͊��oKVw����E���*���.l7���|�~.8�q��4$������gT��~�(� ]K~%���%
v_�<dx���_e!J>@�"Ji2
��#�k����C	��)z�鿮��1@"[��p�y�j��ͭ���ڝd(����MS�����myq�EA��/���	��:���!N�%��@�B}�3m��\��1T�#Z��[�"
�S���v�Y(n��������޶��i^��:���##����Dq���.����p>4�-h7�f���.S~�_�2��W,UPd�'��)r0��r�?�����3�Y]0����!|Ӌ3_�.�
� j��������u�r��	?Ϻ��OW���I�<&�ә��'������Y��;f��V��Q�vZ��=r%7���^��3�sq��Ⱥ��<�z�����62�$�?���:c@M-׼��)*f v�����+X�ؒ��}��(����Əkphll��!$(E����H\�#�ٿ��I�8�vז| ۖB��jG�NP���f�5H�֕p�uУi�̏��e��J;��no�ϐ<��������ڎ�֢��b�_����&��֏�j��3v��)��郛R�h=o3�-�ɴ,�d?��מ���2i&��9@�q��c �1�z�ä9�s� 5�9&\	[
bXW)�F7e�kH�;�?KsJ�/�հv�:�/p6S8L��TU���b!8��;�x@8�����qMnH.Tm"�#:�i�H���dgI���������Hu�H�g��e������;���x�\ԕ?�wv��.��kiќ�H0�Hi+�)�zC���qKWp�������ek�K����XWb�h�$�#��o�a[��'n���� k��zW����lC ꠥ�*G�/4GQu�$TΉ2���b�v�)�������cHG�� +b��h�?������ؘa;מ���uJ+�>~�.��QWT}��#!�MGaF݊����s�5x�Ɯ�Av�pt.�E�����T!KR�T�zpK�^a��yp	Z��ƸA�K�*�x��,"+h�Y��DF�6L>f����ň����#5��^�6҈�)\�I��V7MӦW��_�t��c��Ȥ��P�w��5�Ta��u`�E��c�q�cN��/�!j`��>��I\��Tߦ @���K�5�#%�	�/p�g�����a�V��\�#iq�:��}aǌ|J-PR��Ϭ�x�����aY�0+!z�R,z沊x#�ɧ� ��6�ݱ�4.W
W3~�Z�Vu�N�R[.%�*��<ϴ�c���xh�d*�*�w_P��}�_��hJe@��bِ�gr6���]I}���s�=�<)d��aֵ��-F��_�Pܶ8�O�ȌZ�N���F�uyl5^=P��S���A��2L^�W��Z�K�lx��PY����W'gA�m)���<>���u��e�-*�J�m�)&���+vLcB
E0�'@���0KX:�1d��%JQ�Kz��wl(w_�fZ�	�ƭ>�+#@r��5VB��sn�\�enE30�����%;� ~���-S���4��/dÎ���&��ţ��!m�>�<���4*6���� �k�Y�|<��;��r*�2D��\��B<�y�<\v	/�U9(��GT����s{��^
b��N�m��!%���h;?
��
w��W<Q�̎�/_'uUv� ��߁T[��zиg�%OsDM�N��oP��L�Q�L�qX�(j-�)\B�������?BP��`D�+xs��d�W���L���fL�Y�$������6������R\����lo��J)���"���S���Q�n����3η۸
�Qt���4u���FDś;��fg{	��B*z@�<����!�#��|+>�]�RM�?Q���ܺWҦ��A�'�D�t���|��:����;:��[�1��ƴE!�ju��0B��[+����Q_q
�	D�j|����q���$/�dN���#���5��7�*~A�7���WH}nv�K�5/#��r�}oO�$~o���k��Hȸ%)�����#��B��W<[����])'�J��u��,.z<
 ��q8�ۑ�㙺����@����{�'ry��DgW���(t4�*U~C��D!���]�E�6]���"ёͦ�,N�TH�Ա�ul�����ya��{?,������}F�B�-&����|J�*t����F�$�#�_)����98�qi��s�Jgz�ں��1�fe��Q@g)Ϡ>�8��$�xtIȻE8E�&�e�O���G�v*�+Z��@��3�
�k����j�e,i�rs���e�����u脣�_��wkKڻ�E�}%�6����:�dD�����,y�8�^�5������F��;��팛���#�+�<V�Y%��i�p�KՈ~[�Ş�=iaN�SDgSo�M$�А!����%���@�A7����2�L<��:�������3���U9_���^�[r�7�2M��%)��Dj�e��6!8[S4�W�Z�"��6В'�K���Sa)�B��d�XYS�{hW^0�v�dj*~�|�W?N�1�I�H�ZUC���,L�b'eǺ��Da�L�E3�Z�a��SE�F��� g���I�����KQ$�"�k+iY�T� ��A����O�SQ��8�chǢ#�q���:�$��Q�� !��Ƒq����M���մE�+�
z�[�����3��s��!F'ZO���7�{�z����TXj���0��	�jB��M��뼠������0完鷈)x����^(�c�nԜ����ĒH��=������k�0�d�IV�n"�4��Fc[��.��x�_Ҁ[(-�3>���_�"��9�`H@�pїm�o��`e=�$�}it֦�e][�')��"M<R���q+��V��k��]SϬ��"�ϣ6㗑��n����Hw��,�I{�g`Z�͛�<&�DFߙwO��y�������v��K̅�;m��B���'�6+�����۟o��"t&څц�=��ųe� X*�j��^�=��X�$l�>Q��&�%1�6ho82׶0/�$#D?r�k�5HК\���|��k�]>6��������P�r�����J��>�.z~mf�3�eC��#��w�� �k^o�}�G &9���hie�|��t�]9��((N��������۴X�w�T/"}^W�ݤ�b�>:сA/�;त-$>:�:&��r���`
~1�ݺ��\
8 [��&wܔ�x���@�������\�r9y��da*�?���+�v"�{DύW�'gt/oi`�,��0��$Y7�F�L��' B�����3���<`��&Dڅ�!��F�?�s��[�OL�M�EsY_�[Sc8"�����|�J`-M"�Ƙgm��[�ERK���xr�����1�+�1�;��}	�R��&�"k�"VQ-�uO�>��A�4�X(�����I��=�����etY1՚Dl.���E+����`H6l}�N�/���jQ!�J8��\o�t���yj�+#)��'��Q� ����6{,Cp'����m�F����U�Xs�)s�]@����,)�4:8Q�x�i{xaO�y�w+/�$1�)T�ڋf��,��x_(^�sD����M����>q_��M��	�/��k���1��J�N��}B��I
Y>�4����+C�����L����>����r�n�5`�}[>/�m�P�{M�K�ņ^����_R+LK�B{*� ���I�9��L�5���6����]�[�a�r%���d��"Z[�:r����M��ު�sr�JUjr�]Yc�w�X���SW��2	[8�I��H[�^���t\\����*�M��b�/?��G�E�%���������Ǩ�/i��:���̫��K�o�lw����&j���2kx.(X�,N�f�|�U���̽�},(/W�|��m3�]ݞ4^V=zڎ�%�(�8�Rðgt�CI[��'���0����li�nE6|ݶ,�]8�&���~��;ՎS�^^Ҩa����|J a���A��~~�1���9c�=5�Y�7a�ͤ��j��տ��N�j�.V�ĊM�>s�������F����V�w�I��Fh	��¶�QJ)VN�գ�M�텆�.��Kɮ�����ȍ�5m;A�u,CPNS��7��x��>V��khKb ];���X�KȬ�~�����R�~sl"+���ʜ	U�!�����������A���Wm�=�Q1퍂�����<.U�^�݌���@�~A�f�qS�
n�s��������]ǱS�W�v����6m0g�z,G.	�=��?J���/R���"nK�������)�\�M�֧�R�o��QP��gH���H�S��"�.�Ģ�s��<Nh����r!M�)5ѐ�_���)?��P��ڼ�A��ΆBcs�}��엄N5hmT����<����p�ە���s�ϳ}��k�X�:����/�⤡�|tᐟ[J���l��؞#�S���P��}�T��~�PϚ�,���K���ْ�Ic>VDV�E��@C��ÏN<���R�6�9���#j���!�6��B�d��o��(ǫ?�u�|��l�Ƈh�Rr�T�cm�՜�I�m0Z�0���o���C��@�Jc�Ѫ�m"��9:z��Kލ���c��r����r��'sN���Q��p�'S����U�5`�{�X0�[d[���&�zR�+��١��91�Qs|��o�d��?������nbЄ��47���3��%y��Ʀ�d��H-jz&U�Y�'�zc�k 
#�,��n�K���0������ I]�}�����{���\W@���-�14�!�}ejB�o�0R{cbG�'� Xd�Ek���L��'���7=EKR����
�5G1/E��J����[n�҄
@�*�Q��i1�{�� ,�Y���}��i%5R����G���_3��rg���3,l��������Q>^c#@�N��&yʧ&A��C�h~�5uP.�!�f�V�Cl'֪#IZ�F�
���<V��i,����V�G!�0��~���}��Z�����@���9D�"����Y^��d�Q��/Ep�[�m�ƹ�!�\eB%L�E��L(}Ɲ��	�ک��5����Î�PH�aH��h?��%P�����L�� �ʦ��B)�����C�K3��~\�tk^Iu������ZKh�󱬽�V{��<{�]��zC�`2Qo4q�C�]�uXR�Ѻ�%��;N �J���g4�vp�G%��l�����a��6�_}%� Y@ʑ��cwL�۽@d}J�e��c|j
9���(�E"L����J��b�W�8%�)��r�D+�}��!k�.KUW���QV�!25��� ����z�S!�7������P:<Z�6]���}A�ϔ�i�)dj�`��Pb��>8I��8�b+X9v��_IY��f�fӏ��
���	4�~����'#2��ΦQ�z4����TvN0��T�'�/}bZ��ⰲ�(]1��Xp�;���N��E��9�!z�R����ɏ�.�70U�M���MO6u�ɬ
��*#v�����Sfq�j�˖k6��
�:X?���[��3����4��{��Ol<���|Dl��t$@JMM���ր��{�/�S�.~ecX��D
XP�5��:eL;�%�`���h�&�u��B=x=��a�D=؏���A|&?��^�v��h�a�5a��Z���u|�����T[����FT����?� �ŵ�̍gР;�`�O�v/��BT�y���u������eiKv���5����Yί����Y�M���9�����������t��o��Q�݃�O=I�Im꜑ p�Q���\u���&zñ�2��Mh��a7��m�-'Tؖ:tP�g��e�����9���C��&�8��W������2�z=�M�#�Æ1
��߸%�)���u�Vc09�;Y��M �? >3}%XV]Uh��8����b���뜁�M {���V-�����XVV,�I�S�m��U
biA�j#K��nx��i&���X�l��d9;���2���6�T�j� "��2����&,�� �ihE1x!�����6��g�	-�Ϙ�}'^�و��*�LV!�&��ŃvN@��ۡn���e���Ǔ��[,�5�fH����!J�)�=S<�,��u���c4�z�:N����|�t��+�>�Y`��f2�5T�U��?H�h�����h[M��}Q!�|.ךߥߤ�䑱�\��G��ٖ20 ͂��.Z�!8g�I�}�7T7��˃��M݌�!��J���g�8 ��@3B/%�D� 6�6�0-H��Y�/�D��;��� Vq�뚒|��*�I���Ŝ�*��@8h/�qZ�j2��{&Gv:Ƅ\e����D�OV���� 3��s5t� ��S�H��JuqG�$�{m'��3�D�ţ�Ӭ�d���O���M�r���?(�[|�����u?xg+�z��N������B��^�5�����۩��R���K �|9á5��Aft �T]����8��0�T֓L����W\��A�a�}u�C���cB���BvI���*/��f�1��*��4����*���>�C�&��J8��."�g워X��,���@��E�����L�Pk�P� ��}Z��)��M����}�P����%��aL6�e-]>����:��p�����N�X�c�D����Ү�U��Q����k���:\�c�I��"y�%�p�5:�R���Zρ��wD�k�=%����#�mY��Q䛒8w����f*���̶�B.�M��������-�^j�	���h �^͕��A��=�!��a��U7`4��f2^`�͉ o!�i��p).����n�^<>W��ŕ\,�gb�I\���5�N-[�sH)7�����uj����b3����װ�ٻ�~���p�<����O��6#BڼV�%�*H%���bu��t%m<M��:���F��`� ���"�`�����>6#=i��}��M`Wrnb�-�.=Q2?�I���\(1��z���`,�� 	�׳���	XK	��h��j�љ����*")�J�k�[S7�:��<�L�0��ct��%���|�}6��Z�Q��	�!1,ݖ>��`��>�%���5cJ�H-��u��(Y[�z�Ҭ`ɓ6
�v����m"֑�Pʶ^4y<�(lBg����Q;�@k���g��`�=�NLs�pR5%�������}����m���H\�7��RM��q^?Ip��[f��2��a��u��olS�P,�Z��]�Icr�-�%��q���Y�[Eǯ>��}#���xo�:
Գ���b5c�*y�ކ)��<��x}��0,� ���T�/L����^�j�;��sg@��`�{GŖ�Z��?O��@y��c¤$VD��~��J8�kQx��/&�bx��C�s����\:N�1��G9hHH��dOZ���<��It���]�@��_�}	��K;�9�J�E_�~�-{{wB���K��v��گ��=r�__5����B����p��'oY���o�֋��%=��/����X�a�kk�t�&�Ʉ��`/��9�]�>b