��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߎ[�zZ$D�H�=���3�r�-�7�Y��B
6����I?�����k�'aQ=$ X[Mo�o�����o~��P>��]p�]�9��D���M�y�~I�ʘA��l%�T=���溟q|��iN�NL��zH\M�I���u��L
�{��D 0�w��h�g�>%����2��*u��ПmX��)����/�̑蟕�H�����6[_ �oY&�,P~�
�c��~#�	�5���6VCA�F�_/�c�o�9JW�c#�Et&�.�Zv+^l��!����NB��>��92�L�'�ߩ�Wآ'Smf�8LH琝i�iݴ�`")S���먕���N���t,*�e�^�Ҧ�
���9ӌ������O.EE����J��h���~/ 6�û�p�r2���v"��8�V�u>��#{��k$ݺ08Ls���w6�'c����O!�M��:_v��V$�����8	�&N�գ�a�8�^����[\�Y�����־,��ْ�Ҕ#��]��}?
F����@tFB���Cc �V:�����5gPi��CJ�Ҝ]�H��q]�f�n2۶�0B9�qXgPA��I,3Pj���TyK���Ww�Bu|̳ �˱%�_ަ;G�dT�	������S���Q��<��*���_�&����������\�Y�X�� ϕB����9@�<�=������cM�x�����`j����F�j��d�`�gx<�"��C�R6*�^{Ky,2LZ�g�^D�>�~���d�_)h�(�"r�~�4�娓�^@���F��II¸<x�9����[ʹ^OFS��D���ڴ��qR��P�8bG��,3�3qZݡ��j0B�>ݔ {����!�)? r
ť�\�B8�>��W�o2:���D�E�~��#��l)C�yC�S�vS�bR�.]�w����ÿ���Tq�{"5�\��.����Udj������6����?�������L������w:3|oaz#����rkr�2ؖ@����:�hK3R���_W9�i���K��}x��5���ï��+�<փ9``�d�W�[���kjS�����ټ���`4Y�t;��mGG��*�H��� #'��| �EgUp���)�gAu+S=�+nz��O��*4�4b*�|Q��Ls�2��q�n.Wl��!��Q���+f��-ƈ���{���Q�=����Vdl"���XMPoZ�5���������AK�V���'%��x*ʰ��1�Dn���-1�ĽJ�i�l���=���p��o�������&-�"ς������5G�q�	 �A�fs�D7 ��H�<L*�\7�$߆���y���A�c��������l(��fr�$�sw��7L�d��"ֻ�^��uDmQ؃L��V(H�%�l�-ыW�D_�|��*q�_�ie��DK��2��zb0����9�_��YQ�n���5���~Zgc���yO�D3Û�\��)��jR����@c�Ң�[�::O �yyx4�tY�.�^1U��R���i�~�Ƞ�������H������~��6Ъx��A��5�P��~ǀ!ϑ�n���n�/([6�r�+��zqa Y�?M�_Sf$-�6t.��{"h��	e�\�#!�c�:ZR�*k�E1%,5I���N����P��Uj�
�:x�����W0�u�3LJ����Q��)���l��"i��s�jΐ<R�X-#1�)�A3�)�L��=�;����cK��8��&��'�C�Y�+�;ܸ�*G�>���Ϊ�aٱ?�".�����~E�P�ߘU
 �\�)��zAM܇mxc�4�W�2b���ݔt67i���R�D���T	'Ș���Cl�8��EӡoaY�� 9��A6k��N�h�+O�����&���,�D�֢\�� Gz��g��eN? =�!Jm�"F>�34i�J���q,�6�+�w�a��z�A�>�h�v<Z�����VN�\�.���.w��P���!0*in$T�Eg��H 1�)̳O�:������l�x�z|�i�SaBP��W�� N6�Ք �4"-�0�n��J���ö9�# s��sl +�gv-���#�3N�9�Кq�HY6k�*��I��H+˷~I���4��8p�^r�EĪ'�Zkmq,�u�A��͊��<Wb5Ke�q��E��|x�~�pqڎx1�ϭs�+~,�οV�Ɲ�E\h&s)�DE��%�;y̡p�:ݨ�p@�T�����!�W`v�������NR;Ob�i���_O4��2c��ع��6������̌�p�b�,�����O�K�Ӧ�>�EķR�����ie�h�e���Fx�����mJ��Q����[Q�(o1�W����0����#-��O-ВC���V���09f�fBU�)�I������_�D�rRw7�G� c�n�FfNK�8"5Iz�@�d�t��M���<Xw<{ts�{w�B��P���p��PG��n�O_����_ 3t�����y2i?��['�X�Z�\���#��:/�_��H]u�w�Ɣq�ܯh�
Dߟ?�
.|�[��,I���*r��\/p�?���y׹xؼ@������84�)��"��߉����Ҥ�<
r�no7I�F�v�w]���!%�̔�i���?)4
%˅�nȦ���.L���f\��0���3��`��{J��W�@ � ��9е���AJ�����gO��v�0>F�N \�2@!�I��
��ah��m�^�wX�u�˜A�������79���$�@ixxk���ٮ:�3t��3KvZP���f��/"�
�v?(�C�.�Z%D�$�Xib���HUrBL۫�d[�N����Md*Y�7��{& #UzQ��	���$��3p�2��x�x�^Z�"�a	�G�
~��=A�C8������i�v^�΅A�
��~T��پWޙ�_2�OS��A��D��[Ugـ�9Q0ll��G9}.�j�U��,��;�r}�Y-���=�҃�1�Ccr$7hd����N���#-`��9�9/��D	0ݴ<������s������P���H�O�|\QA�k�S�t�=��_�������S�l�A`�����~C�3�Fn56'�QWʑ������Մ�ǩ֞�~M�4��{��P�����+-y�`u�7�0�� �I����5z����Ai�J�
���v�ϓ�fkj�o����ء���s4��S�^'�Ú�%׳7�<E���Q"�]�U�5J��e2��k�����_���C���h-2"�N���>ͣf0�eC-[�[<7;N�D:I�� ��ϴ�I3�p��1Ĳ�
���338V)�˲���&(�$Q�i�{9)�������6P�_����S�[&����8jlҮ���v�֊�enR����G�lC9�ð�=��7«<��iXh�ӣ�
J.�/~wp"Fo��ÁS<ex#��;����%�J@e��G^+]�x��`��M������-��0ګ�����ͩ���#ł�G���[�ݹۣ2�F)	��k:;t����x"ҳ
�i��Dw'(0^|.���]<�Og��[�s?�ﵦ}y7_n�_��u��j���ue�Ȯ}٥��ة8��͖�+��]��S�ui.�=H ��������=�~��E���L%_�c��q )ūp����Bzn(�ռ.��,��2�D� �
4t��&Չ���U5��ظ��(�Ԯݙϸ[W�����,g��9�f�ܾPyWTu�� *��Ǐ�呗Tm���J���])G^?��A2#F
�i��5�A�\�+��	N$sw��+?9��3��H�[pR��CV�2�E��������x`+o�Ky����M����(�|*+�4H��g�9���)u�:3�=��	>��Z5!�>�@��4����]_�F5��>��:G�+��`|���J\�OW�҂���_+��5g�$"a�3�Y����c˄xV�����������`�(���k&{Da��w������ϴ}٢s�+�a��%?�-n�;ӖગT��˻�l){PE���57�d5C_@@`n�u�A�e�quY6Ю۲bun>w	�?'��G���G[ܺ�I���)7��B�<W~CO�vp�>�˫��h���\�b���h�7UP����6�	��զ��<�"7Y���}[��5�e�+�����<��'��^���֬Z�V��*��: p�dm������U;(�����
<����d��_Y�O��`��nE쯩f��ɲ	r���,/G�๕($Q�@��1I��7g~�1b�(�|}���o���w�L��QW�I�o�h�3���Q�*��\�j��GB�/-LN�W?|(ҝW��骚�D�8.�M��z��Q� k7�cjA����aƞ��n��M`?{&�~H؎�ۮA�3��Tg��e�Z���w�!=55�|�gl�q ���e���$��'z~|�A����w*��D���'�z�-��s�f�n$=��(�|�H��'����^�A�^�`ܽ�x�Y��o^��ä&~��i�S��5@���z�#5���8�]��~�<��吖���o�sD�fMESA;�7wi���b(�͠�7�k���#C4���7��q���>�Ԙ��2W�vn^�e�2���P�~Ӡ��+ �7������F¾� �,ӈ� ���L�>�J�M�ً�kњx�X�8
W�xg���]|�r�'���c�RP4Pp;-�&�n	d�������yc����h,4W�oH�SaRQ�^M�;�洦����x��y��2X�t# 	�[�l;�>4Wp�O����<�)B-�N,�2�M(Z����u�9�ظ7���;���:8�#�e��>��ϯĳ�A2�&�g�X�4~�<��?FO$������`��)���\�/b��ִ�9::J��=�A$4�8|�������{���Y�� �	��DD���kI����� �U63��G}y��8n�#/
!P�b��ʽQ��-�b�!���A1��I6d��W�6��pd���W�7�B*���;Yݱ|����g}ԇ���7��T�!	R%MV�=Ó�z~K�7�@̡��
pV�O��+�ͮ�ĝߧ�_���.�6{]1N����M{�1G�����2�G>
��I�x*��(���Q1���%���"	���j�f1����C��8M.�N	T]�͕�Ɂ]�R�A�.B^�E��6�m�4�Y;�*Z����~��ތ���������P�q ��KN���kv^e���>ʢ���2�H���m�C����-?�݉06� ��J4f�p������)��.�]
���5���+)���QY/S[������׊"����]!��$�`�	�I�t�4N
��y(�զu*ԡ�]l���*�����%�AR�"S�|���h2r��`��>���e�C3�h�K�<J״��\	^7�o��{�O�������0?�V�S?�%m�ۧ;�r��keP�N��BI������E&��t�ր�?s�,0V�6#����6!h����4*��[��K��5��x�DWj.��Z^�՜e2y����a �WФ�c�c�'���$�6ao(�V��^��(���ݸ^��qok���81��Ɔ��tnĆ�I3��*=������9λ"�1ר�Ӧ-t�WZ�2B�_�M��9�p�?	�J�.��H�a0w��-[k�;%*����� �]c������K*i5D�����\�c�3��5�� ��^GM�d�ܔ 0c��h_�����ɛ!%ɥ������'���v%`�� ^u=6����)��:�Z6$ϡ��6�ϟ:�<����J��]0E4bSա��{��LF��T;��@�$�����u���\��ȃ�^%l\z��"�XV]y{���Z�;���yLJd���;a����YK٫��x��IB�C�������L��2)_�R���$��&����Qyf�2�r3d����
o��5|��Z�e��3��ͬt���W3�f�1��@����� e�GW��zj�ADXY�O��T=a2`g�A�dD(1��Au�"az� H�D���hʗ��8�;c�S���Cz����{��o�]�ifFN�/#HK/1�ݺF+v�%
�e_Yİ�S��ע���-l[xo����]譂���T��֛�k]Z����0���b�X;*L�*��BM���#��X�� ���鍅18Rbr��R�0v�.���;ꦬOЭk���;(����� !�ų�%�x}��=!`J
���'�#���Ry[��2����Cf|������C�̪��(�!�e�D�H�^�=�=޶6���SrN{�F�������V���]�+8a�q\��'|���!��%�3#�h"��0��Z"�c�@{)��9�k��1�jߋpw�
�S��cط�l�8)9�G� ٗG��y6Yu��k�a�ÎB�Mf���5>��e��^��3y��+>�_1���`nu����XY�U5�2���ә/�jJ����<dD@T2��CzC4��h-��R;��ȋ��T�o=D"p4����o�F�\k����b��ؖ����O���
M�CQ��D�e�/�A��eU��,�6�=I�m��%��L���Fe{<�9sp�:���WV㖩�_/�`#��-DS��y�0~%Ӟy�٫��䤪��W�'��6E��y�j�Om�ND�$*\��dl*�!v�q���@�p�s4�O�wђ��n��D7@�e��oI�1�$|����ڵ�� Y]��I��*HL�Y�����M�V�Q�e�u�ҷ�s��C�UA�,��?>��	^h�7pEԺ����Gy��OVr�l^C�=��[	�	�n�n��My���:�|�v�:+[��1�WFD<�3�u>��?'���gP�u��z;x?h�!
t7O<8�$=�zƀ��u(�Sc�}�*�Ɏ�KҭZ6��{�5	�9m����:��5�b���f��=��6}��h��Z�e��_g~V�R��c��g��>��P�xX0���f�P�h�M���QY��sN�����^;��W�+{ @+�V�LN����&�R\��f$:�� PdgR=>�s������UM�6L�]2ڂ8�S��<�I,P�;o�X�7�H�?V�I���"�ýժ���&-��F�Vcr)V�z�����+��<�O��`��_���G�G"V�M�*�&�U:�=�R)�qE�Ѵ_a�/�w���ɽIp'�k��.!�"�:��o�>��<C�L�n�m�xnU��'u�$� ����O�9��\0����ϡz���+�_c��Y0ʧlx)��RXCJK�	���a���A	m��~#�d��P��ۭ�6׬dg���]�S�۟�U�����u5���o��������g��bZ���݉�o/�\�~�s	������Ǽ#���Y��<.<k��h��G�G���N���Z��#��a�
�;���ޱ;oṪN���fސc2�͠�D&��l9���I��n��V�[��8E1?\�fO�����t���q��<(�"h�e���͈��)�� <4�S�:=�?���i൓ X��sQ=K�5�
���z*�mʍ`�\���|�<]}���\��o��UX!{�(��}���<�e���ᾡ���v9�^�#�u���Àc�k�D�ڍH���1*�s�^B�Y�d>����Ŧ������ `NF@�.d�M�)_y����b����S`�A������j��<�|���;��{|�!b�4�k?�6t)s"���ӈ��a2�m��J�%���n�d�q�q�������ZV'�Fm �jW\�(.Q�7u�mi!&b�q�����^ڡ��􂭽%4��A�"ך�>� "�t|vg�Z�f���L.��Lbg�:Nj���{X��W�){e\`�!�����YZ��U��c�W!9l@�+Xt��na�;)�VgXA",5Ä�P�� �������P��Q�5v���r�t�ݙA�↥ Ġh�av�;��o���������Q��%�֣�=�S+���ej��+]�UYd[��Ui(�W��~|��]ꙘR�E�(f� �,H���ꯤ��R��M�%G�9_hY�V����i��"ų�ط�K#��k2��1Ë�c���-��}{�f�P!�C�_��+C��8��p�C�w �Q�������am��7a�q������l�����,����S�"���s�X�����$��:U��	�m����໲�ȶnw
��0�cW˸0B��AKUO�	���ӾW!ޗ�kf#`#u�/wK)$��mӑA��E��p{��� (�e}IW_�r�:����d�F�ՙLUm��E��TFn�W���z�{D�cYM���&^��Y�&I2�5�⨍ru�_�az&����y2�.��������0V���"H�dܓ6P��7�ұ�q<Lv�,�A8�o�Y>�jF�������"���(�12�:���I;��o��ˠ�(3eg:�\<р����%��[j�S�s��9�,��FPm�S�
�.�8�vY[�Yu+9�vK'!F%U�"���ibӷ]
@a�Gyӿ�f�u�i.�T�\��^~Q"B�}�-X>k�+�1 qЊ�ۥ�nݳc=tؿ9j�Q�F����+X����=� 9I�����(�X;e�(MPn�9�������2ݥ�h7�|�i�{>I�&�T?���z�(�~����Y���# �_]��:ʌ�f�[ϭu�S��ڻ�+�gJ/��ԅ휯%޸ ڮԆG�;M���DK#X�$�S��>�� Xg;��'"p��r�Z�j&>(��A�`f^`�^Id
�h���i�9��p�7���"�oe�����o�]�����"=Z2z&�����VJj�����)sK}��g���8�� d��1�b���\��?��R���8�!���m�Z6���2��BKՈ�қ�[Si�2�R�NO��j�`8�,�C9��`�l� �*Z�oi-=>�[k�W�l��hU�ܛ�?|%����vF�۫���t2`6)����k����M���Y]�w��I)�7ME�Q�,�z	�]�Y����ps��5}�W�k|��R�������{?��>i����`%z�N�)l0j,���g����K�&,x��z2����`b2[mj�ƪ�$����BJj�~T9I5z���M��{R4FEWs�	MM���Tk�m����KC�Oߙ���[$�cu� �79�!��������)�ܒ�����gF�հ^�-q[$�ڮ��a��k�B��#�w��[h�=�L�&�Hsi����rs���緾�m�������hӊZ�cf�|$� {����e<Q��_`H�2��Yd>�&����lɏjIr���(��� ��q�i9�$�<�:��j-���c�y���WڃTǇ㰕zc~wIlk0��cn��w��_Ć��|����R��]kT3@D��&Q�W̚�~�>�=�Eհ�_w��{����_H2�L�Y ��gR�D�4FL�W��0G��k�#2���Os�=�q[��	�Ji�;fܙ����V��\'�&3�n�N�@@�CJ s�~5��"l�d��<��v���\�n��5����{u[z��6iZ`?<�G)�Tou2")����<��)��C�J5W��BP��9hږέC�y���Ȱ�J_�{��3����D�!Þ	b,R���ܘ�x��4��n�٠�Z�2�r'\\z������k+(Ɛ��H�����|JZ�U�m�N�h�N�������cH���Sӄ��ig��Ż�g� ��*z6-��]+��V";�L���{�}�+o�[s�>��ջ��������..��2[�d%b��HK�#$*תX	��n�#@�[�>�o�%{����J���<q#��0Qԛ��k.�ddX����W��(ܘa�F\B®KV��K3w������9� �5�]>��9:��*�مñ��IAQ�4L6͉ܿ��$Ӗάq��/2jôX :�� �̖r����/��{��d$���6�>j�$0��ym�O|7��n����ʨ��Ën��{���G��P.Ư�{N�A�����*�{�[�qᷦ��_c�45P��X�HQ�u��nqh��U��~�8�\Ͱ��G��	{�q���g8P�>4��S���H���~c�� �	*���)D9��$�a'$Y�BD8#ǌ�2h���b��~��W��Ǎ{���0��.RT6a�����G0�[�!��k�>,R����H�Cu�X�����c�Լ�&w�F��gvх��cuz$x�59:���"��˒�\�"�<Ia�P�l��|~��2�����3�l��Gơ�ԷA�\W(OJ�p���5���C�TԳ� ÷p �֥W��s�,1�o��w�1L:�I
#j�=��7-U��RCaE��͛����+��Bov��}�&⚁�j��!�� �T,Lp!�~D�8�w��
���\<d����Q|%s?3�{��*�:���P��~$�_��ꕕ?��b����,�!������w9O�����&G�!Q�O4����n� ��ˣ��P�Pd�a�!Cg�й��~������h�6{�bN��iZ��ǎ���Ibm9GF�1�.U�B��*��e7 �_����n(h�`�,|���V6�JfjY�0�մ��r<\���Ali\t@�������r%b��yYQ�\��h �Y!�M|�6[��
����M�W���wI�e�x�=�g��^����I�	�?�����>���x_����<y:�7��uPܾ�	e���A��]^�[�󇁥��r��Z�"��y�����e݅XV ��q�X�_M>�4���@�q)M�YdcSDn&T'r����d�/�G��ȡ�hL���T1�(�rA!+�[�
&��OB1�$9���k����WjC�&��Tcx8���gk�Z���q쏝_���Ul(�	��nץ����ܐ?�X��#F�?���兿���Ig�4j2�ɫ��-u���_8���sQN|/��qs1B�a��x��������wN�;1���P4- 9�Lv�����E���q�5�m��j�<�k`B|J�`��m�L�1d�ٹ���^�O�����4``xN�(�|[hUĠ��Ir9�'�]�b 5@{�1��L*rÏ:E��̚H��<���=���Kmg{�)����dl�PP.��9�Y\ ��ҥw�)��bN�q�$@]u���a5��aOP�*�������&��7����B��-�V�\Q�7��s�G��W����⪪:�Wk%&�|Tޏ����L��E�9���}3�N)�"ǝ�qÛZL�(s\d���b�c�&���>J��	��ś��\����y�5S���7��5��o)��Z7�g���oq�a��C�)��|t�*���\&�qZ�W/T��UV�u�ĉ�_V�	�f�?X�ܠC�n�'���o��L ��ވ�9��s�������5E��r΋�\��c�o�FB��FT*g{?�{ʏ����Km�Vz���7]��1&mrSK�,�j�IV��t>�2l�� 1�
xʚ)�i��+�ʇ�6��;	NG.�t�qrC���0��?�~| 	B^*:	�6�.�5R��-��]���<���w4�y��fe~/ܙ��rltɭIЫ>>"gN/{ܱ'�ӯ��
[�Ca^�fR�y���b�%�o�Aw���=�:�Dն�n���j�M���{����1�:�3(/�J�F^�(� hskGs���h�Ib�4�lHz2�h2K���vd,�p�k