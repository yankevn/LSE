��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]呙���疄k��Y����Y�bp\����A!T�3v��Y!�#m굯�H��Ij�	�R��nT�p��z�A��E~�X�P�)�n0�Ӭ���ON�a�: A�,��$9��&>�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�V'w?b�G�F��`�~8Q��	�jv�A��v�q6~���%%���ї�j�t'������E�����eZ���I���Om��W�����mt�auE(+T���c �k
D��.����q5�b�tM7�=	6,6INR}�[��>u�O�G'�mLa��,ǅ���?j�* �?�J�f���l؀����e�_����������<�D���.�!���wf�A��]��~��?p��bBo�>)��4DiEq����Qwj2���Iwƈ�]}`�͝�O�T�t���<��B;�sn�9�ڶ<�k����3ZƦx��&A>��07|�$�%+��`γ`����NG*��*&!W��a��Q�n޼o�3�5L��I���NX#��dǌC��2')�Oc��޷[���gꦧ�p"QE&a:W�L0��g�&����a�n����0�S���tJ�, x���N����%QM�Q�=LRgĞ;$�~u�Y�S��pv%۠@�W���b-�f�W�%3��W�%+����8=��|D(���d�[ 49(�Ei�H��~�� #��in�V�6{y������Ź�P��O�����-TM��3�� b��R�X�H��үPLX�3�l&F�щ(�ź�	ng�"G�tcA�z���0pc�
7K���H_���仰�{�FƮ'�|��"�����(�]��|w6�"��^��	�2�aѵ�D�_���c�,?+��O�).F(������B���p�Hr�ӻ^,�'x/��	�O�j�e&���ݓ����,�󣚪�Q\?��P�$0M�&��[T�.���t��4#�0���{V�LwB�v@���/>��b���w{s)!4��`��p��Y@�.�F�+5��[�n:|*�
��!�'A�jKbyFx�~B�T�a2�"T?�`�K(f��'��HIS�t�}It*/���k�Q#e������\�N�#�3�J1e����i\���O�(�/�F�%t5u�*V��/���j7u��6W�&�0L<�}��<����?᳁S��pȰ�������a�WE�T%�r�1`?�Hd0�c@o�Hh�q�»��+q/Ih��d�����0���*M���Iw��A�⚙\R���=�"�䯁%7��ߞ�E�S�~4Sl4��(�1D�j?�܉��T�X��~��*��J�м�j����v9!���G����FԇQ5J�7���
XB`��[�6%�3Y�!ٴT|��@�7#��_�$sjF��ާ*�;��	����R4ʻ*�H����1e�:.'x*��<�^���Ҋ�s*%:$�^�q�]��;�G�7�������WCYs�j��t�#k\檴'9���pC��K ή���q�e�:=&�T�c%	$�#?46Z��a�ޓ&���z1�nN����q)�2!q�u5VƢ�l�\uFGQ����Q��_+ɮi�w�LQ5���s_�f��`N�y.R��xq��g��}����-�v�d摴�I�^b[��g�e���O�P`�'�����R���0�j��o����OK������r�fնZx�c`)�U��?�f�F�{�4�7$�\�%�p2Q�7��P�G Ns���
�Q�~]a�^����gw�9®�c�}l5�x�V���IË�T�f)�k�o���e���^׾"�{ןf|�k��)����Uw��_q�� K�j����	�A��#�H<����L��
�6�-t��؃������`cƭ!O�r��f�����$x�k��[��[#�_�����,074�<פ���&�sIǴ(K�[rK4Ѥf�e�4D�3���>��|��ߥV���6�M����>���D�O�(���2���ڦQW��LovV���'��j'�>��2��|����Ql�64�f�x�1��z^(o��/���.���V��t�<#s��Kk�&oX%����LқXE�[y�/1#�*���--��%'_E*�j�u�]F�������p�!tI?�G_<���1g7�F���:�n���7���b�ʓcCbѿ�r,i蕜]*T�lK�lp���'.h0�;٤)��g˛��"}:�V���e2�2(-@5�ŒH��G?����/5�D�zF�#a%�r������#�n�6̅oof�L�"� (��},�ۯ�4�:biAD��'�q.f���b��u��&��)������=��XS�4vx�s=;)a��'8_&O���|$H�5���S������x��;��9�C�c�i���u�l�:LŇ�{�&e2�ݼ�#��ʚ#���RX���@�p��̔���9Lќ�e�FG>�v�5�B�OW3>�</3��i���H���	�<����T��<Hv�N�Qy� He���uX�C������Ka˝�l���Yu���N���ea� $�.�:!��*�Ȼ]�EZR*k�e|��M����K��%�֌�^��q��ɳ����h������]�W��V���J_�t�H1	e��y,n��5�|je?��9D�JП�d�ŕ1�}嘾�͑�Pڍ�ǯ���R�H��D��������(�[4\��L�?np4���ej�ژ	�ҷ�﫤��S����QuI{vc>2����\=F��p0 �սJo1��S����"��˱OT@8��-����7Q5���5�?�|���]?ぶ��R:	u�Ǎ��s<n�Fg�Q���x�4�W�����c/��
�G���'�_Q����y�u�>]�w�U��C�y'����S�M�f<���(�l���Q!���J����ጀf�5N�+=4q\,�Sr�s�Y�?�%����Z�P����ڼ텛5�</�S'���~��>#<�.��� �	��"�&��v����xxu6C�D�Yxgo�	��Z��(�11���=�Κ�c-Q�n5>�BDLK��v|Q���<�}R��:Z�DV��c�$u���� �׀|����-��"݀��'���.��̨�����E��SMUw�2C�|Г���X�Y� ܎lq�����